module real_aes_16618_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_1740;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_1767;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_733;
wire n_402;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1691;
wire n_640;
wire n_1721;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_1192;
wire n_518;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI221xp5_ASAP7_75t_L g1272 ( .A1(n_0), .A2(n_89), .B1(n_1000), .B2(n_1253), .C(n_1273), .Y(n_1272) );
AOI22xp33_ASAP7_75t_SL g1292 ( .A1(n_0), .A2(n_200), .B1(n_1293), .B2(n_1295), .Y(n_1292) );
INVx1_ASAP7_75t_L g883 ( .A(n_1), .Y(n_883) );
INVx1_ASAP7_75t_L g326 ( .A(n_2), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_2), .B(n_336), .Y(n_411) );
AND2x2_ASAP7_75t_L g597 ( .A(n_2), .B(n_217), .Y(n_597) );
AND2x2_ASAP7_75t_L g615 ( .A(n_2), .B(n_515), .Y(n_615) );
INVx1_ASAP7_75t_L g1221 ( .A(n_3), .Y(n_1221) );
AOI22xp5_ASAP7_75t_L g1241 ( .A1(n_3), .A2(n_8), .B1(n_626), .B2(n_988), .Y(n_1241) );
AOI22xp5_ASAP7_75t_L g1484 ( .A1(n_4), .A2(n_45), .B1(n_1459), .B2(n_1465), .Y(n_1484) );
INVx1_ASAP7_75t_L g1177 ( .A(n_5), .Y(n_1177) );
INVx1_ASAP7_75t_L g1262 ( .A(n_6), .Y(n_1262) );
OAI22xp33_ASAP7_75t_L g1299 ( .A1(n_6), .A2(n_79), .B1(n_908), .B2(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g692 ( .A(n_7), .Y(n_692) );
OA222x2_ASAP7_75t_L g716 ( .A1(n_7), .A2(n_121), .B1(n_150), .B2(n_717), .C1(n_719), .C2(n_725), .Y(n_716) );
INVx1_ASAP7_75t_L g1231 ( .A(n_8), .Y(n_1231) );
AOI221xp5_ASAP7_75t_L g1252 ( .A1(n_9), .A2(n_78), .B1(n_877), .B2(n_1122), .C(n_1253), .Y(n_1252) );
AOI22xp33_ASAP7_75t_SL g1298 ( .A1(n_9), .A2(n_172), .B1(n_777), .B2(n_1291), .Y(n_1298) );
INVx2_ASAP7_75t_L g365 ( .A(n_10), .Y(n_365) );
INVx1_ASAP7_75t_L g882 ( .A(n_11), .Y(n_882) );
OAI322xp33_ASAP7_75t_L g886 ( .A1(n_11), .A2(n_537), .A3(n_887), .B1(n_892), .B2(n_893), .C1(n_896), .C2(n_902), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g1328 ( .A(n_12), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_13), .A2(n_152), .B1(n_672), .B2(n_679), .Y(n_678) );
INVxp67_ASAP7_75t_SL g749 ( .A(n_13), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_14), .A2(n_198), .B1(n_735), .B2(n_874), .C(n_877), .Y(n_873) );
INVx1_ASAP7_75t_L g895 ( .A(n_14), .Y(n_895) );
INVx1_ASAP7_75t_L g984 ( .A(n_15), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_16), .A2(n_278), .B1(n_919), .B2(n_922), .Y(n_1178) );
INVxp67_ASAP7_75t_SL g1180 ( .A(n_16), .Y(n_1180) );
AOI22xp5_ASAP7_75t_L g1498 ( .A1(n_17), .A2(n_185), .B1(n_1455), .B2(n_1462), .Y(n_1498) );
INVx1_ASAP7_75t_L g1662 ( .A(n_17), .Y(n_1662) );
AOI22xp33_ASAP7_75t_L g1716 ( .A1(n_17), .A2(n_1717), .B1(n_1721), .B2(n_1768), .Y(n_1716) );
INVx1_ASAP7_75t_L g1744 ( .A(n_18), .Y(n_1744) );
AOI221xp5_ASAP7_75t_L g1758 ( .A1(n_18), .A2(n_119), .B1(n_925), .B2(n_1759), .C(n_1761), .Y(n_1758) );
INVx1_ASAP7_75t_L g1430 ( .A(n_19), .Y(n_1430) );
AOI221x1_ASAP7_75t_SL g1435 ( .A1(n_19), .A2(n_169), .B1(n_723), .B2(n_1367), .C(n_1436), .Y(n_1435) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_20), .Y(n_321) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_20), .B(n_319), .Y(n_1456) );
OA22x2_ASAP7_75t_L g343 ( .A1(n_21), .A2(n_344), .B1(n_528), .B2(n_529), .Y(n_343) );
INVxp67_ASAP7_75t_L g529 ( .A(n_21), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g1483 ( .A1(n_21), .A2(n_160), .B1(n_1455), .B2(n_1462), .Y(n_1483) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_22), .A2(n_194), .B1(n_683), .B2(n_790), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_22), .A2(n_262), .B1(n_752), .B2(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_23), .A2(n_261), .B1(n_861), .B2(n_879), .Y(n_878) );
INVxp67_ASAP7_75t_L g890 ( .A(n_23), .Y(n_890) );
INVx1_ASAP7_75t_L g1427 ( .A(n_24), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1440 ( .A1(n_24), .A2(n_153), .B1(n_497), .B2(n_861), .Y(n_1440) );
INVx1_ASAP7_75t_L g413 ( .A(n_25), .Y(n_413) );
INVx1_ASAP7_75t_L g1098 ( .A(n_26), .Y(n_1098) );
OAI22xp5_ASAP7_75t_L g1145 ( .A1(n_26), .A2(n_52), .B1(n_1146), .B2(n_1147), .Y(n_1145) );
INVx1_ASAP7_75t_L g847 ( .A(n_27), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g1489 ( .A1(n_27), .A2(n_242), .B1(n_1455), .B2(n_1462), .Y(n_1489) );
OAI211xp5_ASAP7_75t_SL g980 ( .A1(n_28), .A2(n_981), .B(n_983), .C(n_986), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_28), .A2(n_237), .B1(n_606), .B2(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1170 ( .A(n_29), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_30), .A2(n_259), .B1(n_861), .B2(n_862), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_30), .A2(n_198), .B1(n_675), .B2(n_777), .Y(n_901) );
INVx1_ASAP7_75t_L g1750 ( .A(n_31), .Y(n_1750) );
OAI22xp33_ASAP7_75t_L g1756 ( .A1(n_31), .A2(n_41), .B1(n_941), .B2(n_942), .Y(n_1756) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_32), .A2(n_1347), .B1(n_1348), .B2(n_1349), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_32), .Y(n_1347) );
AOI22xp5_ASAP7_75t_L g1478 ( .A1(n_32), .A2(n_98), .B1(n_1455), .B2(n_1462), .Y(n_1478) );
CKINVDCx5p33_ASAP7_75t_R g1425 ( .A(n_33), .Y(n_1425) );
AOI22xp33_ASAP7_75t_SL g668 ( .A1(n_34), .A2(n_234), .B1(n_669), .B2(n_672), .Y(n_668) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_34), .Y(n_737) );
INVx1_ASAP7_75t_L g937 ( .A(n_35), .Y(n_937) );
AOI22xp5_ASAP7_75t_L g1476 ( .A1(n_36), .A2(n_144), .B1(n_1465), .B2(n_1477), .Y(n_1476) );
OAI22xp5_ASAP7_75t_L g1315 ( .A1(n_37), .A2(n_939), .B1(n_1316), .B2(n_1319), .Y(n_1315) );
INVx1_ASAP7_75t_L g1334 ( .A(n_37), .Y(n_1334) );
INVx1_ASAP7_75t_L g934 ( .A(n_38), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_38), .A2(n_229), .B1(n_645), .B2(n_965), .C(n_966), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g993 ( .A1(n_39), .A2(n_100), .B1(n_994), .B2(n_995), .C(n_996), .Y(n_993) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_39), .A2(n_100), .B1(n_1023), .B2(n_1025), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_40), .A2(n_161), .B1(n_723), .B2(n_751), .Y(n_1368) );
INVx1_ASAP7_75t_L g1396 ( .A(n_40), .Y(n_1396) );
OAI221xp5_ASAP7_75t_L g1746 ( .A1(n_41), .A2(n_270), .B1(n_753), .B2(n_1147), .C(n_1201), .Y(n_1746) );
INVx1_ASAP7_75t_L g1156 ( .A(n_42), .Y(n_1156) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_43), .A2(n_220), .B1(n_1002), .B2(n_1003), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_43), .A2(n_302), .B1(n_560), .B2(n_777), .Y(n_1013) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_44), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g1112 ( .A1(n_46), .A2(n_291), .B1(n_682), .B2(n_685), .C(n_1113), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_46), .A2(n_149), .B1(n_1120), .B2(n_1122), .Y(n_1119) );
AOI21xp5_ASAP7_75t_L g1163 ( .A1(n_47), .A2(n_685), .B(n_777), .Y(n_1163) );
INVxp67_ASAP7_75t_SL g1189 ( .A(n_47), .Y(n_1189) );
INVx1_ASAP7_75t_L g1220 ( .A(n_48), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_48), .A2(n_156), .B1(n_626), .B2(n_965), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_49), .A2(n_170), .B1(n_793), .B2(n_939), .Y(n_1094) );
CKINVDCx5p33_ASAP7_75t_R g1129 ( .A(n_49), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g1739 ( .A(n_50), .Y(n_1739) );
INVx1_ASAP7_75t_L g1322 ( .A(n_51), .Y(n_1322) );
AOI22xp33_ASAP7_75t_L g1342 ( .A1(n_51), .A2(n_55), .B1(n_654), .B2(n_751), .Y(n_1342) );
INVx1_ASAP7_75t_L g1116 ( .A(n_52), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_53), .A2(n_189), .B1(n_826), .B2(n_1256), .Y(n_1370) );
INVx1_ASAP7_75t_L g1391 ( .A(n_53), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g1556 ( .A1(n_54), .A2(n_205), .B1(n_1459), .B2(n_1465), .Y(n_1556) );
AOI221xp5_ASAP7_75t_L g1310 ( .A1(n_55), .A2(n_295), .B1(n_684), .B2(n_1296), .C(n_1311), .Y(n_1310) );
INVxp67_ASAP7_75t_SL g1748 ( .A(n_56), .Y(n_1748) );
OAI22xp5_ASAP7_75t_L g1762 ( .A1(n_56), .A2(n_939), .B1(n_1763), .B2(n_1764), .Y(n_1762) );
OAI221xp5_ASAP7_75t_L g1157 ( .A1(n_57), .A2(n_218), .B1(n_694), .B2(n_941), .C(n_942), .Y(n_1157) );
OAI221xp5_ASAP7_75t_L g1200 ( .A1(n_57), .A2(n_278), .B1(n_753), .B2(n_1147), .C(n_1201), .Y(n_1200) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_58), .A2(n_248), .B1(n_793), .B2(n_939), .Y(n_938) );
INVxp67_ASAP7_75t_SL g945 ( .A(n_58), .Y(n_945) );
INVx1_ASAP7_75t_L g767 ( .A(n_59), .Y(n_767) );
INVx1_ASAP7_75t_L g1099 ( .A(n_60), .Y(n_1099) );
OAI21xp33_ASAP7_75t_L g1144 ( .A1(n_60), .A2(n_725), .B(n_753), .Y(n_1144) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_61), .Y(n_906) );
INVx1_ASAP7_75t_L g869 ( .A(n_62), .Y(n_869) );
OAI211xp5_ASAP7_75t_L g907 ( .A1(n_62), .A2(n_908), .B(n_909), .C(n_912), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g778 ( .A(n_63), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g1674 ( .A(n_64), .Y(n_1674) );
INVx1_ASAP7_75t_L g1752 ( .A(n_65), .Y(n_1752) );
OAI222xp33_ASAP7_75t_L g1755 ( .A1(n_65), .A2(n_255), .B1(n_270), .B2(n_477), .C1(n_488), .C2(n_1047), .Y(n_1755) );
AOI21xp33_ASAP7_75t_L g999 ( .A1(n_66), .A2(n_626), .B(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1009 ( .A(n_66), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_67), .A2(n_276), .B1(n_579), .B2(n_583), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_67), .A2(n_292), .B1(n_624), .B2(n_626), .C(n_628), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_68), .A2(n_147), .B1(n_1462), .B2(n_1465), .Y(n_1461) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_69), .A2(n_157), .B1(n_397), .B2(n_399), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_69), .A2(n_157), .B1(n_511), .B2(n_516), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g1454 ( .A1(n_70), .A2(n_265), .B1(n_1455), .B2(n_1459), .Y(n_1454) );
OAI221xp5_ASAP7_75t_L g1352 ( .A1(n_71), .A2(n_106), .B1(n_642), .B2(n_1070), .C(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1376 ( .A(n_71), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1104 ( .A(n_72), .Y(n_1104) );
AOI22xp5_ASAP7_75t_L g1501 ( .A1(n_73), .A2(n_127), .B1(n_1465), .B2(n_1474), .Y(n_1501) );
INVx1_ASAP7_75t_L g1694 ( .A(n_74), .Y(n_1694) );
OAI211xp5_ASAP7_75t_L g1703 ( .A1(n_74), .A2(n_1704), .B(n_1706), .C(n_1707), .Y(n_1703) );
INVx1_ASAP7_75t_L g452 ( .A(n_75), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g1279 ( .A1(n_76), .A2(n_175), .B1(n_602), .B2(n_606), .Y(n_1279) );
INVx1_ASAP7_75t_L g1355 ( .A(n_77), .Y(n_1355) );
OAI221xp5_ASAP7_75t_SL g1382 ( .A1(n_77), .A2(n_103), .B1(n_547), .B2(n_555), .C(n_570), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_78), .A2(n_236), .B1(n_1290), .B2(n_1291), .Y(n_1289) );
INVx1_ASAP7_75t_L g1260 ( .A(n_79), .Y(n_1260) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_80), .A2(n_283), .B1(n_925), .B2(n_1053), .C(n_1055), .Y(n_1052) );
INVx1_ASAP7_75t_L g1085 ( .A(n_80), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_81), .A2(n_97), .B1(n_682), .B2(n_683), .C(n_685), .Y(n_681) );
AOI22xp33_ASAP7_75t_SL g750 ( .A1(n_81), .A2(n_234), .B1(n_751), .B2(n_752), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g1557 ( .A1(n_82), .A2(n_288), .B1(n_1455), .B2(n_1462), .Y(n_1557) );
CKINVDCx5p33_ASAP7_75t_R g1740 ( .A(n_83), .Y(n_1740) );
INVx1_ASAP7_75t_L g928 ( .A(n_84), .Y(n_928) );
AOI221xp5_ASAP7_75t_L g957 ( .A1(n_84), .A2(n_166), .B1(n_958), .B2(n_959), .C(n_961), .Y(n_957) );
OAI22xp33_ASAP7_75t_L g1330 ( .A1(n_85), .A2(n_122), .B1(n_941), .B2(n_942), .Y(n_1330) );
OAI22xp5_ASAP7_75t_L g1343 ( .A1(n_85), .A2(n_253), .B1(n_1147), .B2(n_1201), .Y(n_1343) );
INVx1_ASAP7_75t_L g455 ( .A(n_86), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g1745 ( .A(n_87), .Y(n_1745) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_88), .A2(n_197), .B1(n_544), .B2(n_552), .C(n_558), .Y(n_543) );
OAI211xp5_ASAP7_75t_L g610 ( .A1(n_88), .A2(n_611), .B(n_616), .C(n_629), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g1297 ( .A1(n_89), .A2(n_240), .B1(n_787), .B2(n_790), .Y(n_1297) );
OAI211xp5_ASAP7_75t_L g1686 ( .A1(n_90), .A2(n_1687), .B(n_1688), .C(n_1691), .Y(n_1686) );
INVx1_ASAP7_75t_L g1710 ( .A(n_90), .Y(n_1710) );
INVx1_ASAP7_75t_L g319 ( .A(n_91), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g1722 ( .A1(n_92), .A2(n_1723), .B1(n_1724), .B2(n_1767), .Y(n_1722) );
CKINVDCx5p33_ASAP7_75t_R g1723 ( .A(n_92), .Y(n_1723) );
INVx1_ASAP7_75t_L g1318 ( .A(n_93), .Y(n_1318) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_93), .A2(n_295), .B1(n_723), .B2(n_751), .Y(n_1339) );
INVx1_ASAP7_75t_L g1749 ( .A(n_94), .Y(n_1749) );
OAI22xp33_ASAP7_75t_L g1697 ( .A1(n_95), .A2(n_258), .B1(n_513), .B2(n_520), .Y(n_1697) );
OAI22xp33_ASAP7_75t_L g1711 ( .A1(n_95), .A2(n_133), .B1(n_398), .B2(n_401), .Y(n_1711) );
AOI221xp5_ASAP7_75t_L g1369 ( .A1(n_96), .A2(n_126), .B1(n_735), .B2(n_990), .C(n_1367), .Y(n_1369) );
INVx1_ASAP7_75t_L g1386 ( .A(n_96), .Y(n_1386) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_97), .A2(n_135), .B1(n_733), .B2(n_735), .C(n_736), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_99), .A2(n_226), .B1(n_602), .B2(n_606), .Y(n_601) );
INVx1_ASAP7_75t_L g1229 ( .A(n_101), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_101), .A2(n_138), .B1(n_723), .B2(n_751), .Y(n_1242) );
XOR2x2_ASAP7_75t_L g1035 ( .A(n_102), .B(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1362 ( .A(n_103), .Y(n_1362) );
CKINVDCx5p33_ASAP7_75t_R g1217 ( .A(n_104), .Y(n_1217) );
INVx1_ASAP7_75t_L g1407 ( .A(n_105), .Y(n_1407) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_105), .A2(n_215), .B1(n_1147), .B2(n_1201), .Y(n_1441) );
INVx1_ASAP7_75t_L g1373 ( .A(n_106), .Y(n_1373) );
INVx1_ASAP7_75t_L g1050 ( .A(n_107), .Y(n_1050) );
INVx1_ASAP7_75t_L g1057 ( .A(n_108), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_109), .A2(n_203), .B1(n_752), .B2(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g1012 ( .A(n_109), .Y(n_1012) );
OAI221xp5_ASAP7_75t_L g1210 ( .A1(n_110), .A2(n_247), .B1(n_793), .B2(n_939), .C(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1245 ( .A(n_110), .Y(n_1245) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_111), .A2(n_764), .B1(n_765), .B2(n_842), .Y(n_763) );
INVx1_ASAP7_75t_L g842 ( .A(n_111), .Y(n_842) );
INVx1_ASAP7_75t_L g1056 ( .A(n_112), .Y(n_1056) );
INVx1_ASAP7_75t_L g1359 ( .A(n_113), .Y(n_1359) );
OAI21xp33_ASAP7_75t_L g1380 ( .A1(n_113), .A2(n_593), .B(n_1381), .Y(n_1380) );
AOI22xp33_ASAP7_75t_SL g1488 ( .A1(n_114), .A2(n_177), .B1(n_1459), .B2(n_1465), .Y(n_1488) );
CKINVDCx5p33_ASAP7_75t_R g1313 ( .A(n_115), .Y(n_1313) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_116), .A2(n_173), .B1(n_919), .B2(n_922), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_116), .A2(n_245), .B1(n_603), .B2(n_758), .Y(n_1066) );
INVx1_ASAP7_75t_L g866 ( .A(n_117), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_118), .A2(n_191), .B1(n_793), .B2(n_939), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g1064 ( .A(n_118), .Y(n_1064) );
INVx1_ASAP7_75t_L g1730 ( .A(n_119), .Y(n_1730) );
INVx1_ASAP7_75t_L g568 ( .A(n_120), .Y(n_568) );
INVx1_ASAP7_75t_L g709 ( .A(n_121), .Y(n_709) );
INVx1_ASAP7_75t_L g1335 ( .A(n_122), .Y(n_1335) );
AOI221xp5_ASAP7_75t_SL g1366 ( .A1(n_123), .A2(n_274), .B1(n_646), .B2(n_735), .C(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1393 ( .A(n_123), .Y(n_1393) );
CKINVDCx5p33_ASAP7_75t_R g1364 ( .A(n_124), .Y(n_1364) );
AOI221xp5_ASAP7_75t_L g854 ( .A1(n_125), .A2(n_180), .B1(n_855), .B2(n_856), .C(n_859), .Y(n_854) );
INVxp67_ASAP7_75t_L g888 ( .A(n_125), .Y(n_888) );
INVx1_ASAP7_75t_L g1397 ( .A(n_126), .Y(n_1397) );
AOI221xp5_ASAP7_75t_L g987 ( .A1(n_128), .A2(n_302), .B1(n_988), .B2(n_989), .C(n_990), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_128), .A2(n_220), .B1(n_777), .B2(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1105 ( .A(n_129), .Y(n_1105) );
AOI22xp33_ASAP7_75t_SL g1125 ( .A1(n_129), .A2(n_141), .B1(n_1126), .B2(n_1127), .Y(n_1125) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_130), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_130), .A2(n_219), .B1(n_624), .B2(n_645), .C(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g1213 ( .A(n_131), .Y(n_1213) );
OAI22xp5_ASAP7_75t_L g1239 ( .A1(n_131), .A2(n_287), .B1(n_603), .B2(n_758), .Y(n_1239) );
CKINVDCx5p33_ASAP7_75t_R g1419 ( .A(n_132), .Y(n_1419) );
OAI22xp33_ASAP7_75t_L g1695 ( .A1(n_133), .A2(n_235), .B1(n_517), .B2(n_1696), .Y(n_1695) );
CKINVDCx5p33_ASAP7_75t_R g1667 ( .A(n_134), .Y(n_1667) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_135), .A2(n_158), .B1(n_675), .B2(n_676), .C(n_677), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g930 ( .A1(n_136), .A2(n_166), .B1(n_925), .B2(n_931), .C(n_933), .Y(n_930) );
INVx1_ASAP7_75t_L g968 ( .A(n_136), .Y(n_968) );
INVxp67_ASAP7_75t_SL g772 ( .A(n_137), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g792 ( .A1(n_137), .A2(n_694), .B1(n_793), .B2(n_795), .C(n_803), .Y(n_792) );
INVx1_ASAP7_75t_L g1223 ( .A(n_138), .Y(n_1223) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_139), .A2(n_677), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g821 ( .A(n_139), .Y(n_821) );
INVx1_ASAP7_75t_L g802 ( .A(n_140), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_140), .A2(n_194), .B1(n_824), .B2(n_826), .Y(n_823) );
INVx1_ASAP7_75t_L g1111 ( .A(n_141), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_142), .A2(n_304), .B1(n_673), .B2(n_684), .Y(n_1173) );
INVxp67_ASAP7_75t_SL g1198 ( .A(n_142), .Y(n_1198) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_143), .A2(n_245), .B1(n_694), .B2(n_941), .C(n_942), .Y(n_1040) );
INVxp67_ASAP7_75t_SL g1062 ( .A(n_143), .Y(n_1062) );
INVx1_ASAP7_75t_L g600 ( .A(n_145), .Y(n_600) );
INVx1_ASAP7_75t_L g1324 ( .A(n_146), .Y(n_1324) );
INVx1_ASAP7_75t_L g1160 ( .A(n_148), .Y(n_1160) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_149), .A2(n_267), .B1(n_677), .B2(n_1053), .C(n_1107), .Y(n_1106) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_150), .A2(n_151), .B1(n_576), .B2(n_702), .C(n_705), .Y(n_701) );
INVxp67_ASAP7_75t_SL g727 ( .A(n_151), .Y(n_727) );
INVxp33_ASAP7_75t_SL g738 ( .A(n_152), .Y(n_738) );
INVx1_ASAP7_75t_L g1421 ( .A(n_153), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_154), .B(n_1458), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_154), .B(n_263), .Y(n_1460) );
INVx2_ASAP7_75t_L g1464 ( .A(n_154), .Y(n_1464) );
XNOR2xp5_ASAP7_75t_L g977 ( .A(n_155), .B(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g1228 ( .A(n_156), .Y(n_1228) );
INVx1_ASAP7_75t_L g746 ( .A(n_158), .Y(n_746) );
INVx1_ASAP7_75t_L g1246 ( .A(n_159), .Y(n_1246) );
AOI22xp5_ASAP7_75t_L g1472 ( .A1(n_159), .A2(n_212), .B1(n_1455), .B2(n_1465), .Y(n_1472) );
INVx1_ASAP7_75t_L g1385 ( .A(n_161), .Y(n_1385) );
INVx1_ASAP7_75t_L g1168 ( .A(n_162), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_163), .A2(n_171), .B1(n_1462), .B2(n_1474), .Y(n_1473) );
OAI221xp5_ASAP7_75t_L g940 ( .A1(n_164), .A2(n_241), .B1(n_694), .B2(n_941), .C(n_942), .Y(n_940) );
INVx1_ASAP7_75t_L g975 ( .A(n_164), .Y(n_975) );
OAI21xp5_ASAP7_75t_SL g1092 ( .A1(n_165), .A2(n_712), .B(n_1093), .Y(n_1092) );
INVx1_ASAP7_75t_L g1115 ( .A(n_165), .Y(n_1115) );
CKINVDCx5p33_ASAP7_75t_R g1673 ( .A(n_167), .Y(n_1673) );
CKINVDCx5p33_ASAP7_75t_R g1416 ( .A(n_168), .Y(n_1416) );
INVx1_ASAP7_75t_L g1423 ( .A(n_169), .Y(n_1423) );
INVx1_ASAP7_75t_L g1138 ( .A(n_170), .Y(n_1138) );
INVxp67_ASAP7_75t_SL g1271 ( .A(n_172), .Y(n_1271) );
OAI211xp5_ASAP7_75t_L g1059 ( .A1(n_173), .A2(n_712), .B(n_1060), .C(n_1063), .Y(n_1059) );
INVx1_ASAP7_75t_L g707 ( .A(n_174), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_174), .A2(n_201), .B1(n_603), .B2(n_758), .Y(n_757) );
OAI211xp5_ASAP7_75t_L g1250 ( .A1(n_175), .A2(n_652), .B(n_1251), .C(n_1259), .Y(n_1250) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_176), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g1668 ( .A(n_178), .Y(n_1668) );
INVx2_ASAP7_75t_L g349 ( .A(n_179), .Y(n_349) );
INVx1_ASAP7_75t_L g484 ( .A(n_179), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_179), .B(n_365), .Y(n_541) );
INVxp67_ASAP7_75t_L g899 ( .A(n_180), .Y(n_899) );
INVx1_ASAP7_75t_L g1028 ( .A(n_181), .Y(n_1028) );
OAI211xp5_ASAP7_75t_L g1095 ( .A1(n_182), .A2(n_694), .B(n_1096), .C(n_1097), .Y(n_1095) );
CKINVDCx5p33_ASAP7_75t_R g1143 ( .A(n_182), .Y(n_1143) );
AOI22xp5_ASAP7_75t_L g1502 ( .A1(n_183), .A2(n_298), .B1(n_1455), .B2(n_1462), .Y(n_1502) );
XOR2xp5_ASAP7_75t_L g1399 ( .A(n_184), .B(n_1400), .Y(n_1399) );
OAI221xp5_ASAP7_75t_SL g1265 ( .A1(n_186), .A2(n_264), .B1(n_1266), .B2(n_1267), .C(n_1268), .Y(n_1265) );
INVx1_ASAP7_75t_L g1283 ( .A(n_186), .Y(n_1283) );
INVx1_ASAP7_75t_L g1232 ( .A(n_187), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_187), .A2(n_281), .B1(n_863), .B2(n_992), .Y(n_1244) );
OAI22xp33_ASAP7_75t_L g1408 ( .A1(n_188), .A2(n_273), .B1(n_464), .B2(n_469), .Y(n_1408) );
INVx1_ASAP7_75t_L g1446 ( .A(n_188), .Y(n_1446) );
INVx1_ASAP7_75t_L g1394 ( .A(n_189), .Y(n_1394) );
INVx1_ASAP7_75t_L g432 ( .A(n_190), .Y(n_432) );
INVxp67_ASAP7_75t_SL g1061 ( .A(n_191), .Y(n_1061) );
BUFx3_ASAP7_75t_L g361 ( .A(n_192), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g1676 ( .A(n_193), .Y(n_1676) );
OAI221xp5_ASAP7_75t_L g1325 ( .A1(n_195), .A2(n_253), .B1(n_785), .B2(n_1326), .C(n_1327), .Y(n_1325) );
OAI211xp5_ASAP7_75t_L g1332 ( .A1(n_195), .A2(n_947), .B(n_1333), .C(n_1336), .Y(n_1332) );
CKINVDCx5p33_ASAP7_75t_R g1312 ( .A(n_196), .Y(n_1312) );
OAI221xp5_ASAP7_75t_SL g631 ( .A1(n_197), .A2(n_286), .B1(n_632), .B2(n_635), .C(n_639), .Y(n_631) );
XOR2xp5_ASAP7_75t_L g1247 ( .A(n_199), .B(n_1248), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_200), .A2(n_240), .B1(n_1255), .B2(n_1257), .Y(n_1254) );
INVx1_ASAP7_75t_L g690 ( .A(n_201), .Y(n_690) );
OAI211xp5_ASAP7_75t_SL g373 ( .A1(n_202), .A2(n_374), .B(n_381), .C(n_385), .Y(n_373) );
INVx1_ASAP7_75t_L g504 ( .A(n_202), .Y(n_504) );
INVx1_ASAP7_75t_L g1017 ( .A(n_203), .Y(n_1017) );
CKINVDCx5p33_ASAP7_75t_R g1278 ( .A(n_204), .Y(n_1278) );
INVx1_ASAP7_75t_L g1176 ( .A(n_206), .Y(n_1176) );
CKINVDCx5p33_ASAP7_75t_R g1670 ( .A(n_207), .Y(n_1670) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_208), .Y(n_771) );
INVx1_ASAP7_75t_L g1048 ( .A(n_209), .Y(n_1048) );
INVx1_ASAP7_75t_L g395 ( .A(n_210), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g491 ( .A1(n_210), .A2(n_492), .B(n_494), .C(n_499), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g1737 ( .A(n_211), .Y(n_1737) );
OAI211xp5_ASAP7_75t_L g1214 ( .A1(n_213), .A2(n_607), .B(n_694), .C(n_1215), .Y(n_1214) );
INVxp33_ASAP7_75t_SL g1238 ( .A(n_213), .Y(n_1238) );
INVx1_ASAP7_75t_L g1039 ( .A(n_214), .Y(n_1039) );
OAI221xp5_ASAP7_75t_L g1412 ( .A1(n_215), .A2(n_231), .B1(n_466), .B2(n_547), .C(n_555), .Y(n_1412) );
INVx1_ASAP7_75t_L g985 ( .A(n_216), .Y(n_985) );
BUFx3_ASAP7_75t_L g336 ( .A(n_217), .Y(n_336) );
INVx1_ASAP7_75t_L g515 ( .A(n_217), .Y(n_515) );
INVxp67_ASAP7_75t_SL g1204 ( .A(n_218), .Y(n_1204) );
INVx1_ASAP7_75t_L g573 ( .A(n_219), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_221), .B(n_838), .Y(n_837) );
CKINVDCx5p33_ASAP7_75t_R g1429 ( .A(n_222), .Y(n_1429) );
OAI322xp33_ASAP7_75t_SL g561 ( .A1(n_223), .A2(n_457), .A3(n_562), .B1(n_567), .B2(n_572), .C1(n_584), .C2(n_587), .Y(n_561) );
OAI22xp33_ASAP7_75t_SL g648 ( .A1(n_223), .A2(n_226), .B1(n_649), .B2(n_652), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g1354 ( .A(n_224), .Y(n_1354) );
INVx1_ASAP7_75t_L g780 ( .A(n_225), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g1320 ( .A(n_227), .Y(n_1320) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_228), .A2(n_290), .B1(n_579), .B2(n_925), .C(n_926), .Y(n_924) );
INVx1_ASAP7_75t_L g962 ( .A(n_228), .Y(n_962) );
INVx1_ASAP7_75t_L g927 ( .A(n_229), .Y(n_927) );
INVx1_ASAP7_75t_L g577 ( .A(n_230), .Y(n_577) );
OA222x2_ASAP7_75t_L g1442 ( .A1(n_231), .A2(n_244), .B1(n_293), .B2(n_717), .C1(n_725), .C2(n_1443), .Y(n_1442) );
XOR2xp5_ASAP7_75t_L g914 ( .A(n_232), .B(n_915), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_233), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g1700 ( .A1(n_235), .A2(n_258), .B1(n_359), .B2(n_1701), .Y(n_1700) );
INVxp67_ASAP7_75t_SL g1269 ( .A(n_236), .Y(n_1269) );
OAI22xp5_ASAP7_75t_SL g531 ( .A1(n_238), .A2(n_532), .B1(n_533), .B2(n_659), .Y(n_531) );
INVx1_ASAP7_75t_L g659 ( .A(n_238), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_238), .A2(n_532), .B1(n_533), .B2(n_659), .Y(n_661) );
AOI211xp5_ASAP7_75t_L g1043 ( .A1(n_239), .A2(n_682), .B(n_1044), .C(n_1046), .Y(n_1043) );
INVx1_ASAP7_75t_L g1079 ( .A(n_239), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g950 ( .A(n_241), .Y(n_950) );
INVx1_ASAP7_75t_L g363 ( .A(n_243), .Y(n_363) );
INVx1_ASAP7_75t_L g379 ( .A(n_243), .Y(n_379) );
INVx1_ASAP7_75t_L g1410 ( .A(n_244), .Y(n_1410) );
CKINVDCx5p33_ASAP7_75t_R g1734 ( .A(n_246), .Y(n_1734) );
INVxp67_ASAP7_75t_SL g1236 ( .A(n_247), .Y(n_1236) );
INVx1_ASAP7_75t_L g956 ( .A(n_248), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_249), .A2(n_280), .B1(n_919), .B2(n_922), .Y(n_918) );
INVx1_ASAP7_75t_L g951 ( .A(n_249), .Y(n_951) );
INVx1_ASAP7_75t_L g437 ( .A(n_250), .Y(n_437) );
AOI21xp33_ASAP7_75t_L g1172 ( .A1(n_251), .A2(n_470), .B(n_677), .Y(n_1172) );
INVxp67_ASAP7_75t_L g1192 ( .A(n_251), .Y(n_1192) );
INVx1_ASAP7_75t_L g441 ( .A(n_252), .Y(n_441) );
INVx1_ASAP7_75t_L g706 ( .A(n_254), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_254), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g1766 ( .A(n_255), .Y(n_1766) );
INVx1_ASAP7_75t_L g418 ( .A(n_256), .Y(n_418) );
AOI22xp5_ASAP7_75t_SL g1497 ( .A1(n_257), .A2(n_307), .B1(n_1465), .B2(n_1474), .Y(n_1497) );
INVxp33_ASAP7_75t_L g894 ( .A(n_259), .Y(n_894) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_260), .Y(n_997) );
INVx1_ASAP7_75t_L g900 ( .A(n_261), .Y(n_900) );
INVx1_ASAP7_75t_L g807 ( .A(n_262), .Y(n_807) );
INVx1_ASAP7_75t_L g1458 ( .A(n_263), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_263), .B(n_1464), .Y(n_1466) );
INVx1_ASAP7_75t_L g1285 ( .A(n_264), .Y(n_1285) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_266), .A2(n_311), .B1(n_357), .B2(n_366), .Y(n_356) );
OAI22xp33_ASAP7_75t_L g519 ( .A1(n_266), .A2(n_311), .B1(n_328), .B2(n_520), .Y(n_519) );
AOI221xp5_ASAP7_75t_SL g1130 ( .A1(n_267), .A2(n_269), .B1(n_1122), .B2(n_1131), .C(n_1132), .Y(n_1130) );
CKINVDCx5p33_ASAP7_75t_R g1671 ( .A(n_268), .Y(n_1671) );
INVx1_ASAP7_75t_L g1110 ( .A(n_269), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_271), .A2(n_1090), .B1(n_1091), .B2(n_1148), .Y(n_1089) );
INVx1_ASAP7_75t_L g1148 ( .A(n_271), .Y(n_1148) );
XOR2x2_ASAP7_75t_L g1152 ( .A(n_272), .B(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1445 ( .A(n_273), .Y(n_1445) );
INVx1_ASAP7_75t_L g1388 ( .A(n_274), .Y(n_1388) );
INVx1_ASAP7_75t_L g1045 ( .A(n_275), .Y(n_1045) );
INVxp67_ASAP7_75t_SL g643 ( .A(n_276), .Y(n_643) );
INVx1_ASAP7_75t_L g781 ( .A(n_277), .Y(n_781) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_277), .A2(n_725), .B1(n_828), .B2(n_833), .C(n_834), .Y(n_827) );
INVx1_ASAP7_75t_L g872 ( .A(n_279), .Y(n_872) );
INVxp67_ASAP7_75t_SL g971 ( .A(n_280), .Y(n_971) );
INVx1_ASAP7_75t_L g1225 ( .A(n_281), .Y(n_1225) );
INVx1_ASAP7_75t_L g391 ( .A(n_282), .Y(n_391) );
INVx1_ASAP7_75t_L g1072 ( .A(n_283), .Y(n_1072) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_284), .Y(n_332) );
INVx1_ASAP7_75t_L g1165 ( .A(n_285), .Y(n_1165) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_286), .Y(n_535) );
INVx1_ASAP7_75t_L g1216 ( .A(n_287), .Y(n_1216) );
CKINVDCx5p33_ASAP7_75t_R g1317 ( .A(n_289), .Y(n_1317) );
INVx1_ASAP7_75t_L g967 ( .A(n_290), .Y(n_967) );
INVx1_ASAP7_75t_L g1134 ( .A(n_291), .Y(n_1134) );
INVx1_ASAP7_75t_L g571 ( .A(n_292), .Y(n_571) );
INVx1_ASAP7_75t_L g1405 ( .A(n_293), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g1732 ( .A(n_294), .Y(n_1732) );
CKINVDCx5p33_ASAP7_75t_R g1693 ( .A(n_296), .Y(n_1693) );
INVx1_ASAP7_75t_L g761 ( .A(n_297), .Y(n_761) );
INVx1_ASAP7_75t_L g354 ( .A(n_299), .Y(n_354) );
INVx2_ASAP7_75t_L g410 ( .A(n_299), .Y(n_410) );
INVx1_ASAP7_75t_L g483 ( .A(n_299), .Y(n_483) );
INVx1_ASAP7_75t_L g935 ( .A(n_300), .Y(n_935) );
INVx1_ASAP7_75t_L g1306 ( .A(n_301), .Y(n_1306) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_303), .Y(n_783) );
INVxp67_ASAP7_75t_SL g1187 ( .A(n_304), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_305), .Y(n_851) );
OAI21xp33_ASAP7_75t_SL g1208 ( .A1(n_306), .A2(n_712), .B(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1212 ( .A(n_306), .Y(n_1212) );
INVx1_ASAP7_75t_L g566 ( .A(n_308), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g1677 ( .A(n_309), .Y(n_1677) );
INVx1_ASAP7_75t_L g426 ( .A(n_310), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_337), .B(n_1448), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_322), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g1715 ( .A(n_316), .B(n_325), .Y(n_1715) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g1720 ( .A(n_318), .B(n_321), .Y(n_1720) );
INVx1_ASAP7_75t_L g1771 ( .A(n_318), .Y(n_1771) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g1774 ( .A(n_321), .B(n_1771), .Y(n_1774) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g525 ( .A(n_325), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g447 ( .A(n_326), .B(n_336), .Y(n_447) );
AND2x4_ASAP7_75t_L g647 ( .A(n_326), .B(n_335), .Y(n_647) );
AND2x4_ASAP7_75t_SL g1714 ( .A(n_327), .B(n_1715), .Y(n_1714) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x6_ASAP7_75t_L g328 ( .A(n_329), .B(n_334), .Y(n_328) );
INVx1_ASAP7_75t_L g417 ( .A(n_329), .Y(n_417) );
OR2x6_ASAP7_75t_L g513 ( .A(n_329), .B(n_514), .Y(n_513) );
BUFx4f_ASAP7_75t_L g1731 ( .A(n_329), .Y(n_1731) );
INVxp67_ASAP7_75t_L g1743 ( .A(n_329), .Y(n_1743) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx4f_ASAP7_75t_L g451 ( .A(n_330), .Y(n_451) );
INVx3_ASAP7_75t_L g619 ( .A(n_330), .Y(n_619) );
INVx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx2_ASAP7_75t_L g424 ( .A(n_332), .Y(n_424) );
INVx2_ASAP7_75t_L g431 ( .A(n_332), .Y(n_431) );
NAND2x1_ASAP7_75t_L g435 ( .A(n_332), .B(n_333), .Y(n_435) );
AND2x2_ASAP7_75t_L g498 ( .A(n_332), .B(n_333), .Y(n_498) );
INVx1_ASAP7_75t_L g509 ( .A(n_332), .Y(n_509) );
AND2x2_ASAP7_75t_L g522 ( .A(n_332), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_333), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g430 ( .A(n_333), .B(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g503 ( .A(n_333), .Y(n_503) );
INVx2_ASAP7_75t_L g523 ( .A(n_333), .Y(n_523) );
INVx1_ASAP7_75t_L g599 ( .A(n_333), .Y(n_599) );
AND2x2_ASAP7_75t_L g655 ( .A(n_333), .B(n_424), .Y(n_655) );
OR2x6_ASAP7_75t_L g1696 ( .A(n_334), .B(n_619), .Y(n_1696) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g496 ( .A(n_335), .Y(n_496) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g502 ( .A(n_336), .Y(n_502) );
AND2x4_ASAP7_75t_L g507 ( .A(n_336), .B(n_508), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_339), .B1(n_1303), .B2(n_1447), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
XNOR2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_843), .Y(n_339) );
XNOR2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_662), .Y(n_340) );
AOI22x1_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_530), .B2(n_660), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g528 ( .A(n_344), .Y(n_528) );
OAI211xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_355), .B(n_404), .C(n_490), .Y(n_344) );
CKINVDCx14_ASAP7_75t_R g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_350), .Y(n_346) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_347), .B(n_350), .Y(n_1712) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp33_ASAP7_75t_SL g460 ( .A(n_349), .B(n_365), .Y(n_460) );
INVx1_ASAP7_75t_L g551 ( .A(n_349), .Y(n_551) );
AND2x2_ASAP7_75t_L g929 ( .A(n_349), .B(n_389), .Y(n_929) );
AND3x4_ASAP7_75t_L g1288 ( .A(n_349), .B(n_389), .C(n_811), .Y(n_1288) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g446 ( .A(n_352), .Y(n_446) );
OR2x2_ASAP7_75t_L g459 ( .A(n_352), .B(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g540 ( .A(n_352), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_SL g1082 ( .A(n_352), .B(n_447), .Y(n_1082) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g527 ( .A(n_353), .Y(n_527) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR3xp33_ASAP7_75t_SL g355 ( .A(n_356), .B(n_373), .C(n_396), .Y(n_355) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
OR2x4_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
OR2x4_ASAP7_75t_L g398 ( .A(n_360), .B(n_368), .Y(n_398) );
BUFx3_ASAP7_75t_L g464 ( .A(n_360), .Y(n_464) );
INVx2_ASAP7_75t_L g487 ( .A(n_360), .Y(n_487) );
BUFx4f_ASAP7_75t_L g801 ( .A(n_360), .Y(n_801) );
BUFx3_ASAP7_75t_L g1047 ( .A(n_360), .Y(n_1047) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx2_ASAP7_75t_L g372 ( .A(n_361), .Y(n_372) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_361), .Y(n_380) );
AND2x4_ASAP7_75t_L g383 ( .A(n_361), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_361), .B(n_379), .Y(n_403) );
INVx1_ASAP7_75t_L g582 ( .A(n_362), .Y(n_582) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g371 ( .A(n_363), .Y(n_371) );
INVx1_ASAP7_75t_L g368 ( .A(n_364), .Y(n_368) );
AND2x4_ASAP7_75t_L g382 ( .A(n_364), .B(n_383), .Y(n_382) );
OR2x6_ASAP7_75t_L g401 ( .A(n_364), .B(n_402), .Y(n_401) );
NAND3x1_ASAP7_75t_L g481 ( .A(n_364), .B(n_482), .C(n_484), .Y(n_481) );
AND2x4_ASAP7_75t_L g550 ( .A(n_364), .B(n_551), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g687 ( .A(n_364), .B(n_484), .Y(n_687) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx3_ASAP7_75t_L g389 ( .A(n_365), .Y(n_389) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_368), .B(n_369), .Y(n_1702) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_369), .Y(n_898) );
BUFx6f_ASAP7_75t_L g1016 ( .A(n_369), .Y(n_1016) );
INVx2_ASAP7_75t_L g1054 ( .A(n_369), .Y(n_1054) );
INVx2_ASAP7_75t_L g1314 ( .A(n_369), .Y(n_1314) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_370), .Y(n_470) );
INVx2_ASAP7_75t_L g477 ( .A(n_370), .Y(n_477) );
BUFx8_ASAP7_75t_L g542 ( .A(n_370), .Y(n_542) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AND2x4_ASAP7_75t_L g581 ( .A(n_372), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x6_ASAP7_75t_L g694 ( .A(n_376), .B(n_695), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g1316 ( .A1(n_376), .A2(n_686), .B1(n_801), .B2(n_1317), .C(n_1318), .Y(n_1316) );
INVx1_ASAP7_75t_L g1705 ( .A(n_376), .Y(n_1705) );
BUFx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_377), .Y(n_467) );
BUFx3_ASAP7_75t_L g570 ( .A(n_377), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
BUFx2_ASAP7_75t_L g394 ( .A(n_378), .Y(n_394) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g384 ( .A(n_379), .Y(n_384) );
BUFx2_ASAP7_75t_L g390 ( .A(n_380), .Y(n_390) );
INVx2_ASAP7_75t_L g547 ( .A(n_380), .Y(n_547) );
AND2x4_ASAP7_75t_L g673 ( .A(n_380), .B(n_557), .Y(n_673) );
CKINVDCx8_ASAP7_75t_R g381 ( .A(n_382), .Y(n_381) );
CKINVDCx8_ASAP7_75t_R g1706 ( .A(n_382), .Y(n_1706) );
BUFx2_ASAP7_75t_L g560 ( .A(n_383), .Y(n_560) );
BUFx2_ASAP7_75t_L g583 ( .A(n_383), .Y(n_583) );
BUFx2_ASAP7_75t_L g675 ( .A(n_383), .Y(n_675) );
BUFx3_ASAP7_75t_L g682 ( .A(n_383), .Y(n_682) );
BUFx2_ASAP7_75t_L g708 ( .A(n_383), .Y(n_708) );
AND2x2_ASAP7_75t_L g923 ( .A(n_383), .B(n_921), .Y(n_923) );
INVx2_ASAP7_75t_L g1020 ( .A(n_383), .Y(n_1020) );
INVx1_ASAP7_75t_L g557 ( .A(n_384), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_391), .B1(n_392), .B2(n_395), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
AND2x4_ASAP7_75t_L g393 ( .A(n_388), .B(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g1708 ( .A(n_388), .B(n_390), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_388), .B(n_394), .Y(n_1709) );
INVx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_391), .A2(n_500), .B1(n_504), .B2(n_505), .Y(n_499) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx3_ASAP7_75t_L g478 ( .A(n_402), .Y(n_478) );
INVx1_ASAP7_75t_L g704 ( .A(n_402), .Y(n_704) );
BUFx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g473 ( .A(n_403), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_456), .Y(n_404) );
OAI33xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_412), .A3(n_425), .B1(n_436), .B2(n_442), .B3(n_448), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_406), .A2(n_742), .B(n_753), .Y(n_741) );
INVx1_ASAP7_75t_L g1136 ( .A(n_406), .Y(n_1136) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx4_ASAP7_75t_L g817 ( .A(n_408), .Y(n_817) );
AOI222xp33_ASAP7_75t_L g952 ( .A1(n_408), .A2(n_740), .B1(n_953), .B2(n_956), .C1(n_957), .C2(n_964), .Y(n_952) );
INVx2_ASAP7_75t_L g1068 ( .A(n_408), .Y(n_1068) );
INVx2_ASAP7_75t_L g1185 ( .A(n_408), .Y(n_1185) );
HB1xp67_ASAP7_75t_L g1434 ( .A(n_408), .Y(n_1434) );
AND2x4_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g658 ( .A(n_409), .Y(n_658) );
OR2x2_ASAP7_75t_L g1398 ( .A(n_409), .B(n_687), .Y(n_1398) );
BUFx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_410), .B(n_597), .Y(n_756) );
INVx2_ASAP7_75t_L g811 ( .A(n_410), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_418), .B2(n_419), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g461 ( .A1(n_413), .A2(n_437), .B1(n_462), .B2(n_465), .Y(n_461) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_416), .A2(n_967), .B1(n_968), .B2(n_969), .Y(n_966) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_418), .A2(n_441), .B1(n_486), .B2(n_488), .Y(n_485) );
INVx5_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx6_ASAP7_75t_L g739 ( .A(n_420), .Y(n_739) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g454 ( .A(n_421), .Y(n_454) );
INVx4_ASAP7_75t_L g622 ( .A(n_421), .Y(n_622) );
INVx2_ASAP7_75t_SL g969 ( .A(n_421), .Y(n_969) );
INVx2_ASAP7_75t_L g1075 ( .A(n_421), .Y(n_1075) );
INVx1_ASAP7_75t_L g1270 ( .A(n_421), .Y(n_1270) );
INVx2_ASAP7_75t_L g1681 ( .A(n_421), .Y(n_1681) );
INVx8_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g518 ( .A(n_422), .B(n_502), .Y(n_518) );
BUFx2_ASAP7_75t_L g1190 ( .A(n_422), .Y(n_1190) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_432), .B2(n_433), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_426), .A2(n_452), .B1(n_469), .B2(n_471), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_427), .A2(n_437), .B1(n_438), .B2(n_441), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g828 ( .A1(n_427), .A2(n_783), .B1(n_798), .B2(n_829), .C(n_830), .Y(n_828) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g1070 ( .A(n_428), .Y(n_1070) );
INVx4_ASAP7_75t_L g1736 ( .A(n_428), .Y(n_1736) );
INVx4_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g745 ( .A(n_430), .Y(n_745) );
INVx2_ASAP7_75t_L g820 ( .A(n_430), .Y(n_820) );
INVx1_ASAP7_75t_L g1194 ( .A(n_430), .Y(n_1194) );
BUFx2_ASAP7_75t_L g1196 ( .A(n_430), .Y(n_1196) );
AND2x2_ASAP7_75t_L g598 ( .A(n_431), .B(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_432), .A2(n_455), .B1(n_475), .B2(n_478), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g1195 ( .A1(n_433), .A2(n_1160), .B1(n_1170), .B2(n_1196), .Y(n_1195) );
OAI221xp5_ASAP7_75t_L g1340 ( .A1(n_433), .A2(n_1312), .B1(n_1317), .B2(n_1341), .C(n_1342), .Y(n_1340) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx4_ASAP7_75t_L g748 ( .A(n_434), .Y(n_748) );
OR2x6_ASAP7_75t_L g753 ( .A(n_434), .B(n_754), .Y(n_753) );
BUFx4f_ASAP7_75t_L g822 ( .A(n_434), .Y(n_822) );
BUFx4f_ASAP7_75t_L g829 ( .A(n_434), .Y(n_829) );
BUFx4f_ASAP7_75t_L g998 ( .A(n_434), .Y(n_998) );
BUFx4f_ASAP7_75t_L g1071 ( .A(n_434), .Y(n_1071) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g440 ( .A(n_435), .Y(n_440) );
INVx5_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g493 ( .A(n_440), .Y(n_493) );
OR2x2_ASAP7_75t_L g725 ( .A(n_440), .B(n_722), .Y(n_725) );
OR2x2_ASAP7_75t_L g974 ( .A(n_440), .B(n_722), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g1683 ( .A1(n_440), .A2(n_1196), .B1(n_1668), .B2(n_1677), .Y(n_1683) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g1337 ( .A1(n_444), .A2(n_1185), .B1(n_1338), .B2(n_1340), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
AND2x4_ASAP7_75t_L g740 ( .A(n_445), .B(n_447), .Y(n_740) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx4_ASAP7_75t_L g628 ( .A(n_447), .Y(n_628) );
INVx4_ASAP7_75t_L g990 ( .A(n_447), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_452), .B1(n_453), .B2(n_455), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g1074 ( .A(n_450), .Y(n_1074) );
INVx2_ASAP7_75t_L g1133 ( .A(n_450), .Y(n_1133) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g642 ( .A(n_451), .Y(n_642) );
INVx4_ASAP7_75t_L g963 ( .A(n_451), .Y(n_963) );
BUFx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI33xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_461), .A3(n_468), .B1(n_474), .B2(n_479), .B3(n_485), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI33xp33_ASAP7_75t_L g1383 ( .A1(n_458), .A2(n_1384), .A3(n_1387), .B1(n_1392), .B2(n_1395), .B3(n_1398), .Y(n_1383) );
OAI33xp33_ASAP7_75t_L g1665 ( .A1(n_458), .A2(n_1398), .A3(n_1666), .B1(n_1669), .B2(n_1672), .B3(n_1675), .Y(n_1665) );
BUFx4f_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx8_ASAP7_75t_L g892 ( .A(n_459), .Y(n_892) );
BUFx2_ASAP7_75t_L g677 ( .A(n_460), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_462), .A2(n_568), .B1(n_569), .B2(n_571), .Y(n_567) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g1055 ( .A1(n_464), .A2(n_570), .B1(n_686), .B2(n_1056), .C(n_1057), .Y(n_1055) );
OAI221xp5_ASAP7_75t_L g1227 ( .A1(n_464), .A2(n_686), .B1(n_1161), .B2(n_1228), .C(n_1229), .Y(n_1227) );
OAI221xp5_ASAP7_75t_L g1763 ( .A1(n_464), .A2(n_570), .B1(n_686), .B2(n_1732), .C(n_1740), .Y(n_1763) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g1219 ( .A1(n_466), .A2(n_929), .B1(n_1008), .B2(n_1220), .C(n_1221), .Y(n_1219) );
OAI22xp33_ASAP7_75t_L g1384 ( .A1(n_466), .A2(n_801), .B1(n_1385), .B2(n_1386), .Y(n_1384) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g489 ( .A(n_467), .Y(n_489) );
OR2x2_ASAP7_75t_L g605 ( .A(n_467), .B(n_540), .Y(n_605) );
INVx4_ASAP7_75t_L g1162 ( .A(n_467), .Y(n_1162) );
OAI221xp5_ASAP7_75t_L g1311 ( .A1(n_467), .A2(n_929), .B1(n_1312), .B2(n_1313), .C(n_1314), .Y(n_1311) );
INVx2_ASAP7_75t_L g676 ( .A(n_469), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g926 ( .A1(n_469), .A2(n_570), .B1(n_927), .B2(n_928), .C(n_929), .Y(n_926) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g576 ( .A(n_470), .Y(n_576) );
INVx2_ASAP7_75t_SL g680 ( .A(n_470), .Y(n_680) );
INVx5_ASAP7_75t_L g1389 ( .A(n_470), .Y(n_1389) );
HB1xp67_ASAP7_75t_L g1418 ( .A(n_470), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1669 ( .A1(n_471), .A2(n_1054), .B1(n_1670), .B2(n_1671), .Y(n_1669) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
CKINVDCx8_ASAP7_75t_R g806 ( .A(n_472), .Y(n_806) );
INVx1_ASAP7_75t_L g1049 ( .A(n_472), .Y(n_1049) );
INVx3_ASAP7_75t_L g1226 ( .A(n_472), .Y(n_1226) );
INVx3_ASAP7_75t_L g1321 ( .A(n_472), .Y(n_1321) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g594 ( .A(n_473), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_475), .A2(n_1390), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g1672 ( .A1(n_475), .A2(n_1390), .B1(n_1673), .B2(n_1674), .Y(n_1672) );
OAI221xp5_ASAP7_75t_L g1761 ( .A1(n_475), .A2(n_570), .B1(n_929), .B2(n_1737), .C(n_1739), .Y(n_1761) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g1326 ( .A(n_476), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_476), .B(n_589), .Y(n_1377) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g565 ( .A(n_477), .Y(n_565) );
OR2x6_ASAP7_75t_SL g793 ( .A(n_477), .B(n_794), .Y(n_793) );
BUFx2_ASAP7_75t_L g1294 ( .A(n_477), .Y(n_1294) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_478), .A2(n_563), .B1(n_564), .B2(n_566), .Y(n_562) );
OAI221xp5_ASAP7_75t_L g572 ( .A1(n_478), .A2(n_573), .B1(n_574), .B2(n_577), .C(n_578), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g896 ( .A1(n_478), .A2(n_897), .B1(n_899), .B2(n_900), .C(n_901), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g1415 ( .A1(n_478), .A2(n_1416), .B1(n_1417), .B2(n_1419), .Y(n_1415) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g1021 ( .A(n_480), .Y(n_1021) );
AOI33xp33_ASAP7_75t_L g1286 ( .A1(n_480), .A2(n_1287), .A3(n_1289), .B1(n_1292), .B2(n_1297), .B3(n_1298), .Y(n_1286) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g586 ( .A(n_481), .Y(n_586) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g549 ( .A(n_483), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_483), .B(n_615), .Y(n_722) );
OR2x2_ASAP7_75t_L g587 ( .A(n_486), .B(n_588), .Y(n_587) );
OR2x6_ASAP7_75t_L g908 ( .A(n_486), .B(n_588), .Y(n_908) );
INVx2_ASAP7_75t_SL g1103 ( .A(n_486), .Y(n_1103) );
OAI22xp33_ASAP7_75t_L g1675 ( .A1(n_486), .A2(n_570), .B1(n_1676), .B2(n_1677), .Y(n_1675) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g1224 ( .A(n_487), .Y(n_1224) );
OAI22xp33_ASAP7_75t_L g893 ( .A1(n_488), .A2(n_799), .B1(n_894), .B2(n_895), .Y(n_893) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g785 ( .A(n_489), .Y(n_785) );
INVx3_ASAP7_75t_L g1171 ( .A(n_489), .Y(n_1171) );
OAI31xp33_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_510), .A3(n_519), .B(n_524), .Y(n_490) );
BUFx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g1191 ( .A1(n_493), .A2(n_1165), .B1(n_1192), .B2(n_1193), .Y(n_1191) );
OAI22xp5_ASAP7_75t_L g1436 ( .A1(n_493), .A2(n_1416), .B1(n_1425), .B2(n_1437), .Y(n_1436) );
OAI22xp5_ASAP7_75t_L g1738 ( .A1(n_493), .A2(n_1077), .B1(n_1739), .B2(n_1740), .Y(n_1738) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_496), .B(n_1690), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_496), .B(n_503), .Y(n_1692) );
AND2x4_ASAP7_75t_SL g614 ( .A(n_497), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g625 ( .A(n_497), .Y(n_625) );
AND2x6_ASAP7_75t_L g630 ( .A(n_497), .B(n_597), .Y(n_630) );
BUFx3_ASAP7_75t_L g735 ( .A(n_497), .Y(n_735) );
BUFx3_ASAP7_75t_L g855 ( .A(n_497), .Y(n_855) );
BUFx3_ASAP7_75t_L g965 ( .A(n_497), .Y(n_965) );
BUFx3_ASAP7_75t_L g988 ( .A(n_497), .Y(n_988) );
BUFx6f_ASAP7_75t_L g1124 ( .A(n_497), .Y(n_1124) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g1275 ( .A(n_498), .Y(n_1275) );
BUFx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g637 ( .A(n_503), .Y(n_637) );
INVx1_ASAP7_75t_L g760 ( .A(n_503), .Y(n_760) );
BUFx2_ASAP7_75t_L g865 ( .A(n_503), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g1691 ( .A1(n_505), .A2(n_1692), .B1(n_1693), .B2(n_1694), .Y(n_1691) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_508), .B(n_597), .Y(n_604) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g521 ( .A(n_514), .B(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_522), .Y(n_627) );
BUFx3_ASAP7_75t_L g645 ( .A(n_522), .Y(n_645) );
INVx2_ASAP7_75t_L g734 ( .A(n_522), .Y(n_734) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx2_ASAP7_75t_L g1698 ( .A(n_525), .Y(n_1698) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g603 ( .A(n_527), .B(n_604), .Y(n_603) );
INVxp67_ASAP7_75t_L g608 ( .A(n_527), .Y(n_608) );
INVx1_ASAP7_75t_L g714 ( .A(n_527), .Y(n_714) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_527), .B(n_604), .Y(n_1147) );
INVxp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND3x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_590), .C(n_609), .Y(n_533) );
AOI211xp5_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_536), .B(n_543), .C(n_561), .Y(n_534) );
INVxp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_538), .A2(n_984), .B1(n_985), .B2(n_1032), .Y(n_1031) );
INVx2_ASAP7_75t_L g1300 ( .A(n_538), .Y(n_1300) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .Y(n_538) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_539), .B(n_1033), .Y(n_1032) );
AND2x4_ASAP7_75t_L g1374 ( .A(n_539), .B(n_1033), .Y(n_1374) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g589 ( .A(n_540), .Y(n_589) );
OR2x2_ASAP7_75t_L g593 ( .A(n_540), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g700 ( .A(n_541), .Y(n_700) );
INVx1_ASAP7_75t_L g921 ( .A(n_541), .Y(n_921) );
INVx3_ASAP7_75t_L g788 ( .A(n_542), .Y(n_788) );
INVx2_ASAP7_75t_SL g804 ( .A(n_542), .Y(n_804) );
INVx2_ASAP7_75t_SL g932 ( .A(n_542), .Y(n_932) );
INVx3_ASAP7_75t_L g1008 ( .A(n_542), .Y(n_1008) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
AND2x6_ASAP7_75t_L g689 ( .A(n_546), .B(n_550), .Y(n_689) );
NAND2x1_ASAP7_75t_L g911 ( .A(n_546), .B(n_548), .Y(n_911) );
AND2x4_ASAP7_75t_SL g1024 ( .A(n_546), .B(n_548), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_546), .B(n_548), .Y(n_1284) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x4_ASAP7_75t_L g553 ( .A(n_548), .B(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g559 ( .A(n_548), .B(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_SL g1026 ( .A(n_548), .B(n_554), .Y(n_1026) );
A2O1A1Ixp33_ASAP7_75t_L g1381 ( .A1(n_548), .A2(n_777), .B(n_1354), .C(n_1382), .Y(n_1381) );
AND2x4_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
OR2x2_ASAP7_75t_L g595 ( .A(n_549), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g954 ( .A(n_549), .Y(n_954) );
NAND2x1p5_ASAP7_75t_L g607 ( .A(n_550), .B(n_581), .Y(n_607) );
AND2x2_ASAP7_75t_L g691 ( .A(n_550), .B(n_556), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_550), .Y(n_695) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_553), .A2(n_866), .B1(n_872), .B2(n_910), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_553), .A2(n_1283), .B1(n_1284), .B2(n_1285), .Y(n_1282) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx3_ASAP7_75t_L g912 ( .A(n_559), .Y(n_912) );
NOR3xp33_ASAP7_75t_L g1005 ( .A(n_559), .B(n_1006), .C(n_1022), .Y(n_1005) );
BUFx2_ASAP7_75t_L g1291 ( .A(n_560), .Y(n_1291) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g889 ( .A(n_565), .Y(n_889) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_566), .A2(n_577), .B1(n_617), .B2(n_620), .C(n_623), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g639 ( .A1(n_568), .A2(n_620), .B1(n_640), .B2(n_643), .C(n_644), .Y(n_639) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g797 ( .A(n_570), .Y(n_797) );
OAI221xp5_ASAP7_75t_L g933 ( .A1(n_570), .A2(n_686), .B1(n_801), .B2(n_934), .C(n_935), .Y(n_933) );
OAI22xp33_ASAP7_75t_L g1395 ( .A1(n_570), .A2(n_801), .B1(n_1396), .B2(n_1397), .Y(n_1395) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_576), .A2(n_1320), .B1(n_1321), .B2(n_1322), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_579), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_705) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx8_ASAP7_75t_L g777 ( .A(n_580), .Y(n_777) );
INVx2_ASAP7_75t_L g1033 ( .A(n_580), .Y(n_1033) );
INVx3_ASAP7_75t_L g1411 ( .A(n_580), .Y(n_1411) );
INVx8_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx3_ASAP7_75t_L g671 ( .A(n_581), .Y(n_671) );
BUFx3_ASAP7_75t_L g684 ( .A(n_581), .Y(n_684) );
AND2x2_ASAP7_75t_L g920 ( .A(n_581), .B(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx2_ASAP7_75t_L g903 ( .A(n_586), .Y(n_903) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_600), .B(n_601), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g904 ( .A1(n_591), .A2(n_883), .B1(n_905), .B2(n_906), .C(n_907), .Y(n_904) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_591), .A2(n_1028), .B(n_1029), .Y(n_1027) );
AOI21xp5_ASAP7_75t_L g1277 ( .A1(n_591), .A2(n_1278), .B(n_1279), .Y(n_1277) );
INVx8_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
BUFx3_ASAP7_75t_L g891 ( .A(n_594), .Y(n_891) );
INVx1_ASAP7_75t_L g1167 ( .A(n_594), .Y(n_1167) );
INVx1_ASAP7_75t_L g718 ( .A(n_595), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_595), .B(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g955 ( .A(n_596), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g638 ( .A(n_597), .Y(n_638) );
AND2x2_ASAP7_75t_L g864 ( .A(n_597), .B(n_865), .Y(n_864) );
AND2x2_ASAP7_75t_L g651 ( .A(n_598), .B(n_615), .Y(n_651) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_598), .Y(n_751) );
INVx3_ASAP7_75t_L g825 ( .A(n_598), .Y(n_825) );
INVx2_ASAP7_75t_L g850 ( .A(n_602), .Y(n_850) );
AND2x4_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx2_ASAP7_75t_SL g836 ( .A(n_603), .Y(n_836) );
AND2x4_ASAP7_75t_L g1030 ( .A(n_603), .B(n_605), .Y(n_1030) );
INVx1_ASAP7_75t_L g1363 ( .A(n_604), .Y(n_1363) );
INVx2_ASAP7_75t_L g1378 ( .A(n_605), .Y(n_1378) );
INVx3_ASAP7_75t_L g905 ( .A(n_606), .Y(n_905) );
OR2x6_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx2_ASAP7_75t_L g710 ( .A(n_607), .Y(n_710) );
OR2x2_ASAP7_75t_L g769 ( .A(n_607), .B(n_608), .Y(n_769) );
OAI31xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_631), .A3(n_648), .B(n_656), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g994 ( .A(n_612), .Y(n_994) );
INVx2_ASAP7_75t_L g1266 ( .A(n_612), .Y(n_1266) );
INVx4_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx3_ASAP7_75t_L g871 ( .A(n_614), .Y(n_871) );
AND2x4_ASAP7_75t_L g634 ( .A(n_615), .B(n_627), .Y(n_634) );
AND2x4_ASAP7_75t_L g653 ( .A(n_615), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g730 ( .A(n_615), .B(n_627), .Y(n_730) );
AND2x2_ASAP7_75t_L g982 ( .A(n_615), .B(n_723), .Y(n_982) );
BUFx2_ASAP7_75t_L g1356 ( .A(n_615), .Y(n_1356) );
OAI22xp5_ASAP7_75t_L g1197 ( .A1(n_617), .A2(n_1168), .B1(n_1190), .B2(n_1198), .Y(n_1197) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
BUFx3_ASAP7_75t_L g1084 ( .A(n_619), .Y(n_1084) );
BUFx6f_ASAP7_75t_L g1188 ( .A(n_619), .Y(n_1188) );
BUFx3_ASAP7_75t_L g1437 ( .A(n_619), .Y(n_1437) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_622), .A2(n_935), .B1(n_962), .B2(n_963), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g1684 ( .A1(n_622), .A2(n_963), .B1(n_1671), .B2(n_1674), .Y(n_1684) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g958 ( .A(n_625), .Y(n_958) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g858 ( .A(n_627), .Y(n_858) );
HB1xp67_ASAP7_75t_SL g877 ( .A(n_628), .Y(n_877) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_630), .A2(n_871), .B1(n_872), .B2(n_873), .C(n_878), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g986 ( .A1(n_630), .A2(n_987), .B(n_991), .Y(n_986) );
AOI21xp5_ASAP7_75t_L g1251 ( .A1(n_630), .A2(n_1252), .B(n_1254), .Y(n_1251) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx6f_ASAP7_75t_L g881 ( .A(n_634), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_634), .A2(n_650), .B1(n_984), .B2(n_985), .Y(n_983) );
INVx1_ASAP7_75t_L g1264 ( .A(n_634), .Y(n_1264) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g995 ( .A(n_636), .Y(n_995) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g1360 ( .A(n_638), .Y(n_1360) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_642), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g960 ( .A(n_645), .Y(n_960) );
BUFx2_ASAP7_75t_L g1253 ( .A(n_645), .Y(n_1253) );
INVx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g859 ( .A(n_647), .Y(n_859) );
INVx2_ASAP7_75t_L g1000 ( .A(n_647), .Y(n_1000) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
HB1xp67_ASAP7_75t_L g1261 ( .A(n_650), .Y(n_1261) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_L g713 ( .A(n_651), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g868 ( .A(n_651), .Y(n_868) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g880 ( .A1(n_653), .A2(n_881), .B1(n_882), .B2(n_883), .Y(n_880) );
BUFx2_ASAP7_75t_L g826 ( .A(n_654), .Y(n_826) );
INVx1_ASAP7_75t_L g1258 ( .A(n_654), .Y(n_1258) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g724 ( .A(n_655), .Y(n_724) );
BUFx3_ASAP7_75t_L g752 ( .A(n_655), .Y(n_752) );
BUFx3_ASAP7_75t_L g863 ( .A(n_655), .Y(n_863) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_657), .A2(n_666), .B(n_711), .Y(n_665) );
INVx2_ASAP7_75t_L g943 ( .A(n_657), .Y(n_943) );
OAI31xp33_ASAP7_75t_SL g1093 ( .A1(n_657), .A2(n_1094), .A3(n_1095), .B(n_1100), .Y(n_1093) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_658), .B(n_841), .Y(n_840) );
AOI21xp5_ASAP7_75t_SL g1350 ( .A1(n_658), .A2(n_1351), .B(n_1365), .Y(n_1350) );
INVx1_ASAP7_75t_L g1432 ( .A(n_658), .Y(n_1432) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
XNOR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_763), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_761), .B(n_762), .Y(n_663) );
AND3x1_ASAP7_75t_L g664 ( .A(n_665), .B(n_715), .C(n_731), .Y(n_664) );
AOI31xp33_ASAP7_75t_L g762 ( .A1(n_665), .A2(n_715), .A3(n_731), .B(n_761), .Y(n_762) );
NAND3xp33_ASAP7_75t_SL g666 ( .A(n_667), .B(n_688), .C(n_696), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_674), .B1(n_678), .B2(n_681), .Y(n_667) );
BUFx2_ASAP7_75t_SL g1290 ( .A(n_669), .Y(n_1290) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
BUFx3_ASAP7_75t_L g1113 ( .A(n_671), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_671), .B(n_1328), .Y(n_1327) );
BUFx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx5_ASAP7_75t_L g791 ( .A(n_673), .Y(n_791) );
AND2x4_ASAP7_75t_L g841 ( .A(n_673), .B(n_700), .Y(n_841) );
BUFx3_ASAP7_75t_L g925 ( .A(n_673), .Y(n_925) );
BUFx12f_ASAP7_75t_L g1296 ( .A(n_673), .Y(n_1296) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_675), .A2(n_771), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g1760 ( .A(n_684), .Y(n_1760) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g795 ( .A1(n_686), .A2(n_796), .B1(n_798), .B2(n_799), .C(n_802), .Y(n_795) );
OAI221xp5_ASAP7_75t_L g1420 ( .A1(n_686), .A2(n_1047), .B1(n_1421), .B2(n_1422), .C(n_1423), .Y(n_1420) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_691), .B2(n_692), .C(n_693), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_689), .A2(n_691), .B1(n_780), .B2(n_781), .Y(n_779) );
INVx4_ASAP7_75t_L g941 ( .A(n_689), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_689), .A2(n_691), .B1(n_1098), .B2(n_1099), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_689), .A2(n_691), .B1(n_1216), .B2(n_1217), .Y(n_1215) );
INVx2_ASAP7_75t_L g942 ( .A(n_691), .Y(n_942) );
NOR3xp33_ASAP7_75t_L g1309 ( .A(n_693), .B(n_1310), .C(n_1315), .Y(n_1309) );
NOR3xp33_ASAP7_75t_L g1757 ( .A(n_693), .B(n_1758), .C(n_1762), .Y(n_1757) );
CKINVDCx5p33_ASAP7_75t_R g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g1413 ( .A(n_695), .Y(n_1413) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_701), .B1(n_709), .B2(n_710), .Y(n_696) );
INVxp67_ASAP7_75t_L g775 ( .A(n_697), .Y(n_775) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
BUFx2_ASAP7_75t_L g1329 ( .A(n_699), .Y(n_1329) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g794 ( .A(n_700), .Y(n_794) );
OAI21xp33_ASAP7_75t_L g1011 ( .A1(n_702), .A2(n_1012), .B(n_1013), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1424 ( .A1(n_702), .A2(n_1425), .B1(n_1426), .B2(n_1427), .Y(n_1424) );
INVx3_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g1390 ( .A(n_704), .Y(n_1390) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_708), .Y(n_1107) );
AOI211xp5_ASAP7_75t_SL g936 ( .A1(n_710), .A2(n_937), .B(n_938), .C(n_940), .Y(n_936) );
AOI211xp5_ASAP7_75t_L g1038 ( .A1(n_710), .A2(n_1039), .B(n_1040), .C(n_1041), .Y(n_1038) );
INVx2_ASAP7_75t_L g1096 ( .A(n_710), .Y(n_1096) );
AOI211xp5_ASAP7_75t_L g1155 ( .A1(n_710), .A2(n_1156), .B(n_1157), .C(n_1158), .Y(n_1155) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_710), .A2(n_1324), .B1(n_1325), .B2(n_1329), .C(n_1330), .Y(n_1323) );
AOI221xp5_ASAP7_75t_L g1754 ( .A1(n_710), .A2(n_1329), .B1(n_1749), .B2(n_1755), .C(n_1756), .Y(n_1754) );
INVx1_ASAP7_75t_L g1181 ( .A(n_712), .Y(n_1181) );
INVx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI222xp33_ASAP7_75t_L g766 ( .A1(n_713), .A2(n_729), .B1(n_767), .B2(n_768), .C1(n_771), .C2(n_772), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_713), .B(n_971), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_713), .B(n_1328), .Y(n_1331) );
AOI22xp33_ASAP7_75t_SL g1444 ( .A1(n_713), .A2(n_729), .B1(n_1445), .B2(n_1446), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1751 ( .A(n_713), .B(n_1752), .Y(n_1751) );
AND2x4_ASAP7_75t_L g729 ( .A(n_714), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_726), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g770 ( .A(n_720), .Y(n_770) );
AOI222xp33_ASAP7_75t_L g949 ( .A1(n_720), .A2(n_835), .B1(n_836), .B2(n_937), .C1(n_950), .C2(n_951), .Y(n_949) );
AOI222xp33_ASAP7_75t_L g1060 ( .A1(n_720), .A2(n_953), .B1(n_973), .B2(n_1039), .C1(n_1061), .C2(n_1062), .Y(n_1060) );
AOI211xp5_ASAP7_75t_L g1142 ( .A1(n_720), .A2(n_1143), .B(n_1144), .C(n_1145), .Y(n_1142) );
AOI222xp33_ASAP7_75t_L g1203 ( .A1(n_720), .A2(n_953), .B1(n_973), .B2(n_1156), .C1(n_1177), .C2(n_1204), .Y(n_1203) );
AOI21xp33_ASAP7_75t_L g1237 ( .A1(n_720), .A2(n_1238), .B(n_1239), .Y(n_1237) );
INVx1_ASAP7_75t_L g1443 ( .A(n_720), .Y(n_1443) );
AOI222xp33_ASAP7_75t_L g1747 ( .A1(n_720), .A2(n_953), .B1(n_973), .B2(n_1748), .C1(n_1749), .C2(n_1750), .Y(n_1747) );
AND2x4_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
AOI332xp33_ASAP7_75t_L g1333 ( .A1(n_721), .A2(n_723), .A3(n_954), .B1(n_955), .B2(n_973), .B3(n_1324), .C1(n_1334), .C2(n_1335), .Y(n_1333) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx3_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g1003 ( .A(n_724), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g947 ( .A(n_729), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_729), .B(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1140 ( .A(n_729), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_729), .B(n_1176), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_729), .B(n_1236), .Y(n_1235) );
NAND2xp33_ASAP7_75t_SL g1765 ( .A(n_729), .B(n_1766), .Y(n_1765) );
AOI211xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_740), .B(n_741), .C(n_757), .Y(n_731) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g876 ( .A(n_734), .Y(n_876) );
OAI221xp5_ASAP7_75t_L g1439 ( .A1(n_739), .A2(n_1193), .B1(n_1419), .B2(n_1429), .C(n_1440), .Y(n_1439) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_740), .Y(n_833) );
AOI322xp5_ASAP7_75t_L g1118 ( .A1(n_740), .A2(n_953), .A3(n_1119), .B1(n_1125), .B2(n_1129), .C1(n_1130), .C2(n_1136), .Y(n_1118) );
AOI332xp33_ASAP7_75t_L g1240 ( .A1(n_740), .A2(n_816), .A3(n_953), .B1(n_1241), .B2(n_1242), .B3(n_1243), .C1(n_1244), .C2(n_1245), .Y(n_1240) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_746), .B1(n_747), .B2(n_749), .C(n_750), .Y(n_742) );
INVx3_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_745), .A2(n_822), .B1(n_1313), .B2(n_1320), .C(n_1339), .Y(n_1338) );
OAI22xp5_ASAP7_75t_L g1682 ( .A1(n_747), .A2(n_1341), .B1(n_1670), .B2(n_1673), .Y(n_1682) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g1080 ( .A(n_748), .Y(n_1080) );
INVx1_ASAP7_75t_L g1687 ( .A(n_748), .Y(n_1687) );
INVx2_ASAP7_75t_L g1735 ( .A(n_748), .Y(n_1735) );
INVx3_ASAP7_75t_L g832 ( .A(n_751), .Y(n_832) );
BUFx6f_ASAP7_75t_L g1256 ( .A(n_751), .Y(n_1256) );
OAI21xp5_ASAP7_75t_SL g813 ( .A1(n_753), .A2(n_814), .B(n_818), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g976 ( .A(n_753), .Y(n_976) );
OAI21xp5_ASAP7_75t_L g1438 ( .A1(n_753), .A2(n_833), .B(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NAND2x2_ASAP7_75t_L g758 ( .A(n_755), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g835 ( .A(n_758), .Y(n_835) );
HB1xp67_ASAP7_75t_L g1146 ( .A(n_758), .Y(n_1146) );
INVx2_ASAP7_75t_SL g1202 ( .A(n_758), .Y(n_1202) );
INVx2_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_773), .C(n_812), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
OAI21xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_792), .B(n_808), .Y(n_773) );
OAI211xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_776), .B(n_779), .C(n_782), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_778), .A2(n_780), .B1(n_835), .B2(n_836), .Y(n_834) );
OAI211xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B(n_786), .C(n_789), .Y(n_782) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g1764 ( .A1(n_788), .A2(n_1226), .B1(n_1734), .B2(n_1745), .Y(n_1764) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g1175 ( .A(n_793), .Y(n_1175) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g1666 ( .A1(n_801), .A2(n_1171), .B1(n_1667), .B2(n_1668), .Y(n_1666) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_805), .B1(n_806), .B2(n_807), .Y(n_803) );
OAI221xp5_ASAP7_75t_L g818 ( .A1(n_805), .A2(n_819), .B1(n_821), .B2(n_822), .C(n_823), .Y(n_818) );
OAI221xp5_ASAP7_75t_L g1014 ( .A1(n_806), .A2(n_997), .B1(n_1015), .B2(n_1017), .C(n_1018), .Y(n_1014) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g885 ( .A(n_809), .Y(n_885) );
A2O1A1Ixp33_ASAP7_75t_SL g1154 ( .A1(n_809), .A2(n_1155), .B(n_1174), .C(n_1179), .Y(n_1154) );
BUFx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_810), .Y(n_1004) );
BUFx2_ASAP7_75t_L g1276 ( .A(n_810), .Y(n_1276) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI31xp33_ASAP7_75t_SL g1209 ( .A1(n_811), .A2(n_1210), .A3(n_1214), .B(n_1218), .Y(n_1209) );
NOR3xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_827), .C(n_837), .Y(n_812) );
INVxp67_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
BUFx2_ASAP7_75t_L g1078 ( .A(n_820), .Y(n_1078) );
INVx2_ASAP7_75t_L g1341 ( .A(n_820), .Y(n_1341) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g861 ( .A(n_825), .Y(n_861) );
INVx2_ASAP7_75t_SL g992 ( .A(n_825), .Y(n_992) );
INVx1_ASAP7_75t_L g1002 ( .A(n_825), .Y(n_1002) );
INVx1_ASAP7_75t_L g1126 ( .A(n_825), .Y(n_1126) );
A2O1A1Ixp33_ASAP7_75t_L g1358 ( .A1(n_831), .A2(n_855), .B(n_1359), .C(n_1360), .Y(n_1358) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx3_ASAP7_75t_L g939 ( .A(n_841), .Y(n_939) );
AOI221xp5_ASAP7_75t_L g1174 ( .A1(n_841), .A2(n_1175), .B1(n_1176), .B2(n_1177), .C(n_1178), .Y(n_1174) );
XNOR2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_1087), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_1034), .B1(n_1035), .B2(n_1086), .Y(n_844) );
INVx1_ASAP7_75t_L g1086 ( .A(n_845), .Y(n_1086) );
XOR2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_913), .Y(n_845) );
XNOR2x1_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
AND2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_904), .Y(n_848) );
AOI221xp5_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_851), .B1(n_852), .B2(n_884), .C(n_886), .Y(n_849) );
NAND3xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_870), .C(n_880), .Y(n_852) );
AOI222xp33_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_860), .B1(n_864), .B2(n_866), .C1(n_867), .C2(n_869), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_855), .A2(n_863), .B1(n_1354), .B2(n_1355), .Y(n_1353) );
BUFx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g989 ( .A(n_858), .Y(n_989) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_863), .Y(n_879) );
INVx1_ASAP7_75t_SL g1128 ( .A(n_863), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g1361 ( .A1(n_864), .A2(n_1362), .B1(n_1363), .B2(n_1364), .Y(n_1361) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g1121 ( .A(n_876), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1131 ( .A(n_876), .Y(n_1131) );
INVx2_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_890), .B2(n_891), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g1101 ( .A1(n_891), .A2(n_1102), .B1(n_1104), .B2(n_1105), .C(n_1106), .Y(n_1101) );
OAI221xp5_ASAP7_75t_L g1108 ( .A1(n_891), .A2(n_1109), .B1(n_1110), .B2(n_1111), .C(n_1112), .Y(n_1108) );
CKINVDCx20_ASAP7_75t_R g1010 ( .A(n_892), .Y(n_1010) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g1109 ( .A(n_898), .Y(n_1109) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_SL g1301 ( .A(n_912), .Y(n_1301) );
XNOR2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_977), .Y(n_913) );
OR2x2_ASAP7_75t_L g915 ( .A(n_916), .B(n_948), .Y(n_915) );
A2O1A1Ixp33_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_936), .B(n_943), .C(n_944), .Y(n_916) );
NOR3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_924), .C(n_930), .Y(n_917) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_920), .A2(n_923), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
AOI22xp5_ASAP7_75t_L g1211 ( .A1(n_920), .A2(n_923), .B1(n_1212), .B2(n_1213), .Y(n_1211) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
AOI221xp5_ASAP7_75t_SL g1404 ( .A1(n_925), .A2(n_1405), .B1(n_1406), .B2(n_1407), .C(n_1408), .Y(n_1404) );
OAI21xp33_ASAP7_75t_L g1044 ( .A1(n_929), .A2(n_1008), .B(n_1045), .Y(n_1044) );
OAI221xp5_ASAP7_75t_L g1428 ( .A1(n_929), .A2(n_1015), .B1(n_1161), .B2(n_1429), .C(n_1430), .Y(n_1428) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_932), .A2(n_1165), .B1(n_1166), .B2(n_1168), .Y(n_1164) );
INVx1_ASAP7_75t_L g1058 ( .A(n_943), .Y(n_1058) );
A2O1A1Ixp33_ASAP7_75t_L g1753 ( .A1(n_943), .A2(n_1754), .B(n_1757), .C(n_1765), .Y(n_1753) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
NAND4xp25_ASAP7_75t_L g948 ( .A(n_949), .B(n_952), .C(n_970), .D(n_972), .Y(n_948) );
AND2x4_ASAP7_75t_L g953 ( .A(n_954), .B(n_955), .Y(n_953) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g1679 ( .A1(n_963), .A2(n_1667), .B1(n_1676), .B2(n_1680), .Y(n_1679) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_969), .A2(n_1050), .B1(n_1084), .B2(n_1085), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g1135 ( .A(n_969), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g1729 ( .A1(n_969), .A2(n_1730), .B1(n_1731), .B2(n_1732), .Y(n_1729) );
OAI22xp5_ASAP7_75t_L g1741 ( .A1(n_969), .A2(n_1742), .B1(n_1744), .B2(n_1745), .Y(n_1741) );
AOI21xp5_ASAP7_75t_L g972 ( .A1(n_973), .A2(n_975), .B(n_976), .Y(n_972) );
AOI21xp5_ASAP7_75t_L g1234 ( .A1(n_973), .A2(n_976), .B(n_1217), .Y(n_1234) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
OR3x1_ASAP7_75t_L g1065 ( .A(n_976), .B(n_1066), .C(n_1067), .Y(n_1065) );
NOR3xp33_ASAP7_75t_L g1336 ( .A(n_976), .B(n_1337), .C(n_1343), .Y(n_1336) );
AND4x1_ASAP7_75t_L g978 ( .A(n_979), .B(n_1005), .C(n_1027), .D(n_1031), .Y(n_978) );
OAI21xp33_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_993), .B(n_1004), .Y(n_979) );
INVx2_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
BUFx2_ASAP7_75t_L g1267 ( .A(n_995), .Y(n_1267) );
OAI211xp5_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_998), .B(n_999), .C(n_1001), .Y(n_996) );
A2O1A1Ixp33_ASAP7_75t_L g1308 ( .A1(n_1004), .A2(n_1309), .B(n_1323), .C(n_1331), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1011), .B1(n_1014), .B2(n_1021), .Y(n_1006) );
OAI21xp5_ASAP7_75t_L g1007 ( .A1(n_1008), .A2(n_1009), .B(n_1010), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_1008), .A2(n_1166), .B1(n_1231), .B2(n_1232), .Y(n_1230) );
INVx2_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1020), .Y(n_1406) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
AOI211x1_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1058), .B(n_1059), .C(n_1065), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1042), .Y(n_1037) );
NOR3xp33_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1051), .C(n_1052), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_1045), .A2(n_1070), .B1(n_1071), .B2(n_1072), .Y(n_1069) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1048), .B1(n_1049), .B2(n_1050), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_1048), .A2(n_1057), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_1056), .A2(n_1077), .B1(n_1079), .B2(n_1080), .Y(n_1076) );
OAI33xp33_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1069), .A3(n_1073), .B1(n_1076), .B2(n_1081), .B3(n_1083), .Y(n_1067) );
INVx4_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
OAI33xp33_ASAP7_75t_L g1678 ( .A1(n_1081), .A2(n_1185), .A3(n_1679), .B1(n_1682), .B2(n_1683), .B3(n_1684), .Y(n_1678) );
OAI33xp33_ASAP7_75t_L g1728 ( .A1(n_1081), .A2(n_1185), .A3(n_1729), .B1(n_1733), .B2(n_1738), .B3(n_1741), .Y(n_1728) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1082), .Y(n_1199) );
OA22x2_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1149), .B1(n_1150), .B2(n_1302), .Y(n_1087) );
HB1xp67_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1089), .Y(n_1302) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
NOR2x1_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1117), .Y(n_1091) );
NAND3xp33_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1108), .C(n_1114), .Y(n_1100) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
OAI22xp5_ASAP7_75t_SL g1132 ( .A1(n_1104), .A2(n_1133), .B1(n_1134), .B2(n_1135), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1137), .Y(n_1117) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1121), .Y(n_1367) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_SL g1127 ( .A(n_1128), .Y(n_1127) );
OAI221xp5_ASAP7_75t_L g1268 ( .A1(n_1133), .A2(n_1269), .B1(n_1270), .B2(n_1271), .C(n_1272), .Y(n_1268) );
AOI21xp5_ASAP7_75t_L g1137 ( .A1(n_1138), .A2(n_1139), .B(n_1141), .Y(n_1137) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
XNOR2xp5_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1247), .Y(n_1150) );
XNOR2xp5_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1206), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1182), .Y(n_1153) );
OAI21xp33_ASAP7_75t_L g1158 ( .A1(n_1159), .A2(n_1164), .B(n_1169), .Y(n_1158) );
OAI21xp33_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1161), .B(n_1163), .Y(n_1159) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1162), .Y(n_1422) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
OAI211xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1171), .B(n_1172), .C(n_1173), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1181), .Y(n_1179) );
NAND3xp33_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1203), .C(n_1205), .Y(n_1182) );
NOR2xp33_ASAP7_75t_SL g1183 ( .A(n_1184), .B(n_1200), .Y(n_1183) );
OAI33xp33_ASAP7_75t_L g1184 ( .A1(n_1185), .A2(n_1186), .A3(n_1191), .B1(n_1195), .B2(n_1197), .B3(n_1199), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g1186 ( .A1(n_1187), .A2(n_1188), .B1(n_1189), .B2(n_1190), .Y(n_1186) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
XOR2x2_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1246), .Y(n_1206) );
NOR2xp33_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1233), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1222), .B1(n_1227), .B2(n_1230), .Y(n_1218) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1224), .B1(n_1225), .B2(n_1226), .Y(n_1222) );
BUFx4f_ASAP7_75t_SL g1426 ( .A(n_1224), .Y(n_1426) );
NAND4xp25_ASAP7_75t_SL g1233 ( .A(n_1234), .B(n_1235), .C(n_1237), .D(n_1240), .Y(n_1233) );
NAND3xp33_ASAP7_75t_SL g1248 ( .A(n_1249), .B(n_1277), .C(n_1280), .Y(n_1248) );
OAI21xp33_ASAP7_75t_L g1249 ( .A1(n_1250), .A2(n_1265), .B(n_1276), .Y(n_1249) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_1260), .A2(n_1261), .B1(n_1262), .B2(n_1263), .Y(n_1259) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
BUFx2_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1275), .Y(n_1690) );
NOR3xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1299), .C(n_1301), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1286), .Y(n_1281) );
BUFx3_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
BUFx2_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVxp67_ASAP7_75t_SL g1447 ( .A(n_1303), .Y(n_1447) );
XOR2xp5_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1344), .Y(n_1303) );
HB1xp67_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
XNOR2x1_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1307), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1332), .Y(n_1307) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1329), .Y(n_1403) );
HB1xp67_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
XNOR2xp5_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1399), .Y(n_1345) );
INVx2_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1371), .Y(n_1349) );
AOI21xp5_ASAP7_75t_L g1351 ( .A1(n_1352), .A2(n_1356), .B(n_1357), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1361), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1375 ( .A1(n_1364), .A2(n_1376), .B1(n_1377), .B2(n_1378), .Y(n_1375) );
AOI22xp5_ASAP7_75t_L g1365 ( .A1(n_1366), .A2(n_1368), .B1(n_1369), .B2(n_1370), .Y(n_1365) );
NAND3xp33_ASAP7_75t_SL g1371 ( .A(n_1372), .B(n_1375), .C(n_1379), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1373), .B(n_1374), .Y(n_1372) );
NOR2xp33_ASAP7_75t_SL g1379 ( .A(n_1380), .B(n_1383), .Y(n_1379) );
OAI22xp5_ASAP7_75t_L g1387 ( .A1(n_1388), .A2(n_1389), .B1(n_1390), .B2(n_1391), .Y(n_1387) );
NAND4xp75_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1433), .C(n_1442), .D(n_1444), .Y(n_1400) );
OAI21x1_ASAP7_75t_L g1401 ( .A1(n_1402), .A2(n_1414), .B(n_1431), .Y(n_1401) );
OAI21xp5_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1404), .B(n_1409), .Y(n_1402) );
A2O1A1Ixp33_ASAP7_75t_L g1409 ( .A1(n_1410), .A2(n_1411), .B(n_1412), .C(n_1413), .Y(n_1409) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_1415), .A2(n_1420), .B1(n_1424), .B2(n_1428), .Y(n_1414) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
AOI211x1_ASAP7_75t_L g1433 ( .A1(n_1434), .A2(n_1435), .B(n_1438), .C(n_1441), .Y(n_1433) );
OAI221xp5_ASAP7_75t_L g1448 ( .A1(n_1449), .A2(n_1656), .B1(n_1659), .B2(n_1713), .C(n_1716), .Y(n_1448) );
AOI211xp5_ASAP7_75t_L g1449 ( .A1(n_1450), .A2(n_1570), .B(n_1616), .C(n_1640), .Y(n_1449) );
OAI211xp5_ASAP7_75t_L g1450 ( .A1(n_1451), .A2(n_1467), .B(n_1512), .C(n_1558), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1451), .B(n_1591), .Y(n_1590) );
OAI211xp5_ASAP7_75t_L g1640 ( .A1(n_1451), .A2(n_1641), .B(n_1643), .C(n_1649), .Y(n_1640) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
OAI221xp5_ASAP7_75t_L g1542 ( .A1(n_1452), .A2(n_1543), .B1(n_1549), .B2(n_1552), .C(n_1554), .Y(n_1542) );
OAI32xp33_ASAP7_75t_L g1608 ( .A1(n_1452), .A2(n_1513), .A3(n_1530), .B1(n_1565), .B2(n_1609), .Y(n_1608) );
OAI221xp5_ASAP7_75t_L g1616 ( .A1(n_1452), .A2(n_1541), .B1(n_1617), .B2(n_1624), .C(n_1626), .Y(n_1616) );
INVx3_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
INVx3_ASAP7_75t_L g1536 ( .A(n_1453), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1453), .B(n_1540), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1453), .B(n_1486), .Y(n_1553) );
OR2x2_ASAP7_75t_L g1575 ( .A(n_1453), .B(n_1508), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1453), .B(n_1499), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1453), .B(n_1524), .Y(n_1632) );
NAND2xp5_ASAP7_75t_L g1639 ( .A(n_1453), .B(n_1508), .Y(n_1639) );
NOR2xp33_ASAP7_75t_L g1644 ( .A(n_1453), .B(n_1645), .Y(n_1644) );
AND2x4_ASAP7_75t_SL g1453 ( .A(n_1454), .B(n_1461), .Y(n_1453) );
AND2x6_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1457), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1456), .B(n_1460), .Y(n_1459) );
AND2x4_ASAP7_75t_L g1462 ( .A(n_1456), .B(n_1463), .Y(n_1462) );
AND2x6_ASAP7_75t_L g1465 ( .A(n_1456), .B(n_1466), .Y(n_1465) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1456), .B(n_1460), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1456), .B(n_1460), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1456), .B(n_1463), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1458), .B(n_1464), .Y(n_1463) );
HB1xp67_ASAP7_75t_L g1772 ( .A(n_1463), .Y(n_1772) );
AOI221xp5_ASAP7_75t_L g1467 ( .A1(n_1468), .A2(n_1479), .B1(n_1490), .B2(n_1507), .C(n_1509), .Y(n_1467) );
A2O1A1Ixp33_ASAP7_75t_SL g1537 ( .A1(n_1468), .A2(n_1518), .B(n_1538), .C(n_1539), .Y(n_1537) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1468), .Y(n_1568) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1469), .B(n_1475), .Y(n_1468) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
OR2x2_ASAP7_75t_L g1530 ( .A(n_1470), .B(n_1475), .Y(n_1530) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
OR2x2_ASAP7_75t_L g1494 ( .A(n_1471), .B(n_1495), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1471), .B(n_1495), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1521 ( .A(n_1471), .B(n_1496), .Y(n_1521) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1471), .Y(n_1533) );
NOR2xp33_ASAP7_75t_L g1545 ( .A(n_1471), .B(n_1475), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1473), .Y(n_1471) );
NOR2xp33_ASAP7_75t_L g1492 ( .A(n_1475), .B(n_1482), .Y(n_1492) );
CKINVDCx5p33_ASAP7_75t_R g1506 ( .A(n_1475), .Y(n_1506) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1475), .B(n_1482), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1548 ( .A(n_1475), .B(n_1505), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1475), .B(n_1521), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1475), .B(n_1533), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1622 ( .A(n_1475), .B(n_1623), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1478), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1476), .B(n_1478), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1485), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1480), .B(n_1532), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1544 ( .A(n_1480), .B(n_1545), .Y(n_1544) );
OR2x2_ASAP7_75t_L g1585 ( .A(n_1480), .B(n_1548), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1480), .B(n_1524), .Y(n_1615) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1480), .B(n_1513), .Y(n_1650) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1503 ( .A(n_1481), .B(n_1504), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1481), .B(n_1510), .Y(n_1559) );
NOR2xp33_ASAP7_75t_L g1563 ( .A(n_1481), .B(n_1530), .Y(n_1563) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1481), .B(n_1513), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1481), .B(n_1577), .Y(n_1576) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1481), .B(n_1520), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1588 ( .A(n_1481), .B(n_1515), .Y(n_1588) );
INVx3_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx2_ASAP7_75t_L g1518 ( .A(n_1482), .Y(n_1518) );
NAND2xp5_ASAP7_75t_L g1603 ( .A(n_1482), .B(n_1486), .Y(n_1603) );
OR2x2_ASAP7_75t_L g1645 ( .A(n_1482), .B(n_1515), .Y(n_1645) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1484), .Y(n_1482) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1486), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1624 ( .A(n_1486), .B(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1487), .B(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1487), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1487), .B(n_1508), .Y(n_1524) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1487), .Y(n_1541) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1489), .Y(n_1487) );
OAI32xp33_ASAP7_75t_L g1490 ( .A1(n_1491), .A2(n_1493), .A3(n_1499), .B1(n_1500), .B2(n_1503), .Y(n_1490) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1492), .B(n_1510), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1493), .B(n_1551), .Y(n_1550) );
NAND2xp5_ASAP7_75t_SL g1565 ( .A(n_1493), .B(n_1518), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1493), .B(n_1506), .Y(n_1607) );
OAI21xp5_ASAP7_75t_L g1612 ( .A1(n_1493), .A2(n_1613), .B(n_1615), .Y(n_1612) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1493), .B(n_1511), .Y(n_1619) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1495), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1495), .B(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1496), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1497), .B(n_1498), .Y(n_1496) );
OAI21xp33_ASAP7_75t_L g1561 ( .A1(n_1499), .A2(n_1562), .B(n_1564), .Y(n_1561) );
AOI221xp5_ASAP7_75t_L g1649 ( .A1(n_1499), .A2(n_1531), .B1(n_1650), .B2(n_1651), .C(n_1652), .Y(n_1649) );
INVx2_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
AOI22xp33_ASAP7_75t_L g1543 ( .A1(n_1500), .A2(n_1544), .B1(n_1546), .B2(n_1547), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1500), .B(n_1515), .Y(n_1546) );
CKINVDCx6p67_ASAP7_75t_R g1594 ( .A(n_1500), .Y(n_1594) );
AND2x4_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1502), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1501), .B(n_1502), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1505), .B(n_1506), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1506), .B(n_1521), .Y(n_1520) );
OR2x2_ASAP7_75t_L g1525 ( .A(n_1506), .B(n_1526), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1506), .B(n_1532), .Y(n_1531) );
OR2x2_ASAP7_75t_L g1564 ( .A(n_1506), .B(n_1565), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1506), .B(n_1629), .Y(n_1628) );
OR2x2_ASAP7_75t_L g1535 ( .A(n_1507), .B(n_1536), .Y(n_1535) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1507), .Y(n_1610) );
OR2x2_ASAP7_75t_L g1514 ( .A(n_1508), .B(n_1515), .Y(n_1514) );
AOI21xp33_ASAP7_75t_L g1583 ( .A1(n_1508), .A2(n_1554), .B(n_1584), .Y(n_1583) );
NAND2xp5_ASAP7_75t_SL g1599 ( .A(n_1508), .B(n_1600), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1508), .B(n_1536), .Y(n_1655) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1509), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1642 ( .A(n_1509), .B(n_1540), .Y(n_1642) );
AND2x2_ASAP7_75t_L g1651 ( .A(n_1509), .B(n_1541), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1511), .Y(n_1509) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1510), .Y(n_1526) );
AOI211xp5_ASAP7_75t_L g1512 ( .A1(n_1513), .A2(n_1516), .B(n_1522), .C(n_1542), .Y(n_1512) );
INVx2_ASAP7_75t_SL g1513 ( .A(n_1514), .Y(n_1513) );
NOR2xp33_ASAP7_75t_L g1597 ( .A(n_1514), .B(n_1598), .Y(n_1597) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
OR2x2_ASAP7_75t_L g1517 ( .A(n_1518), .B(n_1519), .Y(n_1517) );
INVx2_ASAP7_75t_L g1529 ( .A(n_1518), .Y(n_1529) );
NAND2xp5_ASAP7_75t_SL g1582 ( .A(n_1518), .B(n_1546), .Y(n_1582) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1518), .B(n_1602), .Y(n_1636) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1521), .Y(n_1631) );
OAI211xp5_ASAP7_75t_L g1522 ( .A1(n_1523), .A2(n_1525), .B(n_1527), .C(n_1537), .Y(n_1522) );
CKINVDCx14_ASAP7_75t_R g1523 ( .A(n_1524), .Y(n_1523) );
NOR2xp33_ASAP7_75t_L g1572 ( .A(n_1525), .B(n_1535), .Y(n_1572) );
OR2x2_ASAP7_75t_L g1614 ( .A(n_1526), .B(n_1551), .Y(n_1614) );
OAI21xp5_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1531), .B(n_1534), .Y(n_1527) );
NOR2xp33_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1530), .Y(n_1528) );
AOI311xp33_ASAP7_75t_L g1604 ( .A1(n_1529), .A2(n_1574), .A3(n_1605), .B(n_1608), .C(n_1611), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1529), .B(n_1531), .Y(n_1638) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1531), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1532), .B(n_1551), .Y(n_1577) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1532), .Y(n_1630) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
NAND2xp5_ASAP7_75t_L g1609 ( .A(n_1536), .B(n_1610), .Y(n_1609) );
AOI221xp5_ASAP7_75t_L g1578 ( .A1(n_1539), .A2(n_1579), .B1(n_1581), .B2(n_1590), .C(n_1592), .Y(n_1578) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1540), .Y(n_1566) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
AOI21xp5_ASAP7_75t_L g1652 ( .A1(n_1549), .A2(n_1653), .B(n_1654), .Y(n_1652) );
CKINVDCx5p33_ASAP7_75t_R g1549 ( .A(n_1550), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1551), .B(n_1559), .Y(n_1627) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1554), .Y(n_1591) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1556), .B(n_1557), .Y(n_1555) );
AOI221xp5_ASAP7_75t_L g1558 ( .A1(n_1559), .A2(n_1560), .B1(n_1561), .B2(n_1566), .C(n_1567), .Y(n_1558) );
INVxp33_ASAP7_75t_SL g1562 ( .A(n_1563), .Y(n_1562) );
OAI31xp33_ASAP7_75t_L g1634 ( .A1(n_1566), .A2(n_1584), .A3(n_1613), .B(n_1635), .Y(n_1634) );
NOR2xp33_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1569), .Y(n_1567) );
OAI211xp5_ASAP7_75t_L g1581 ( .A1(n_1568), .A2(n_1582), .B(n_1583), .C(n_1586), .Y(n_1581) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_1568), .B(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1569), .Y(n_1646) );
NAND3xp33_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1578), .C(n_1604), .Y(n_1570) );
NOR2xp33_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1573), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1574), .B(n_1576), .Y(n_1573) );
AOI22xp33_ASAP7_75t_SL g1617 ( .A1(n_1574), .A2(n_1618), .B1(n_1620), .B2(n_1621), .Y(n_1617) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1577), .Y(n_1648) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1589), .Y(n_1586) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
OAI211xp5_ASAP7_75t_L g1592 ( .A1(n_1593), .A2(n_1595), .B(n_1596), .C(n_1599), .Y(n_1592) );
CKINVDCx6p67_ASAP7_75t_R g1593 ( .A(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
INVxp33_ASAP7_75t_SL g1653 ( .A(n_1600), .Y(n_1653) );
NOR2xp33_ASAP7_75t_L g1600 ( .A(n_1601), .B(n_1603), .Y(n_1600) );
CKINVDCx14_ASAP7_75t_R g1601 ( .A(n_1602), .Y(n_1601) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
INVxp67_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1614), .B(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
O2A1O1Ixp33_ASAP7_75t_L g1626 ( .A1(n_1627), .A2(n_1628), .B(n_1632), .C(n_1633), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1631), .Y(n_1629) );
AOI21xp5_ASAP7_75t_L g1633 ( .A1(n_1634), .A2(n_1637), .B(n_1639), .Y(n_1633) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
OAI21xp33_ASAP7_75t_L g1643 ( .A1(n_1644), .A2(n_1646), .B(n_1647), .Y(n_1643) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
CKINVDCx20_ASAP7_75t_R g1656 ( .A(n_1657), .Y(n_1656) );
CKINVDCx5p33_ASAP7_75t_R g1657 ( .A(n_1658), .Y(n_1657) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
HB1xp67_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
XNOR2xp5_ASAP7_75t_L g1661 ( .A(n_1662), .B(n_1663), .Y(n_1661) );
AND3x1_ASAP7_75t_L g1663 ( .A(n_1664), .B(n_1685), .C(n_1699), .Y(n_1663) );
NOR2xp33_ASAP7_75t_SL g1664 ( .A(n_1665), .B(n_1678), .Y(n_1664) );
BUFx6f_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
OAI31xp33_ASAP7_75t_L g1685 ( .A1(n_1686), .A2(n_1695), .A3(n_1697), .B(n_1698), .Y(n_1685) );
INVx2_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
AOI22xp33_ASAP7_75t_SL g1707 ( .A1(n_1693), .A2(n_1708), .B1(n_1709), .B2(n_1710), .Y(n_1707) );
OAI31xp33_ASAP7_75t_SL g1699 ( .A1(n_1700), .A2(n_1703), .A3(n_1711), .B(n_1712), .Y(n_1699) );
INVx2_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
INVx3_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
HB1xp67_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
BUFx3_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
BUFx3_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
INVxp33_ASAP7_75t_SL g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1724), .Y(n_1767) );
INVxp67_ASAP7_75t_SL g1724 ( .A(n_1725), .Y(n_1724) );
NOR2x1_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1753), .Y(n_1725) );
NAND3xp33_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1747), .C(n_1751), .Y(n_1726) );
NOR2xp33_ASAP7_75t_L g1727 ( .A(n_1728), .B(n_1746), .Y(n_1727) );
OAI22xp5_ASAP7_75t_L g1733 ( .A1(n_1734), .A2(n_1735), .B1(n_1736), .B2(n_1737), .Y(n_1733) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
HB1xp67_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
HB1xp67_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
OAI21xp5_ASAP7_75t_L g1770 ( .A1(n_1771), .A2(n_1772), .B(n_1773), .Y(n_1770) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
endmodule