module fake_jpeg_19256_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_21),
.B1(n_32),
.B2(n_22),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_53),
.B1(n_54),
.B2(n_62),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_32),
.B1(n_21),
.B2(n_16),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_21),
.B1(n_32),
.B2(n_18),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_26),
.B1(n_18),
.B2(n_25),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_20),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_26),
.B1(n_25),
.B2(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_28),
.B1(n_20),
.B2(n_33),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_16),
.B1(n_41),
.B2(n_28),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_82),
.Y(n_108)
);

NAND2xp67_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_38),
.Y(n_66)
);

XNOR2x1_ASAP7_75t_SL g109 ( 
.A(n_66),
.B(n_49),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_15),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_28),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_50),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_45),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_80),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_15),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_28),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_45),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_59),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_33),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_48),
.C(n_59),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_109),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_70),
.B1(n_65),
.B2(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_112),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_47),
.B(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_107),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_86),
.B1(n_74),
.B2(n_84),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_104),
.B1(n_110),
.B2(n_89),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g103 ( 
.A(n_66),
.B(n_55),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_55),
.B1(n_63),
.B2(n_49),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_52),
.C(n_48),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_65),
.C(n_27),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_48),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_49),
.B1(n_31),
.B2(n_27),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_31),
.Y(n_112)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_27),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_24),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_72),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_123),
.B1(n_134),
.B2(n_90),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_87),
.B1(n_65),
.B2(n_82),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_76),
.B1(n_88),
.B2(n_78),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_135),
.Y(n_152)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_70),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_110),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_88),
.B1(n_71),
.B2(n_3),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_69),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_92),
.B(n_108),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_99),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_161),
.B1(n_1),
.B2(n_2),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_148),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_163),
.B1(n_133),
.B2(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_98),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_113),
.B(n_91),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_160),
.B(n_24),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_154),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_91),
.C(n_108),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_131),
.C(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_162),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_108),
.B(n_105),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_95),
.B1(n_93),
.B2(n_111),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_93),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_97),
.B(n_114),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_164),
.A2(n_121),
.B(n_118),
.C(n_114),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_159),
.B(n_116),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_117),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_174),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

AO21x1_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_125),
.B(n_128),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_175),
.B1(n_183),
.B2(n_185),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_126),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_181),
.Y(n_187)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_114),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_149),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_1),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_184),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_5),
.B(n_6),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_151),
.C(n_156),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_193),
.C(n_147),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_154),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_204),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_156),
.C(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_150),
.B1(n_158),
.B2(n_155),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_171),
.B1(n_175),
.B2(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_162),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_160),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_158),
.B1(n_164),
.B2(n_149),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_207),
.A2(n_218),
.B1(n_219),
.B2(n_188),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_172),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_212),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_180),
.B(n_183),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_213),
.B(n_187),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_198),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_175),
.B(n_185),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_175),
.C(n_165),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_190),
.C(n_200),
.Y(n_224)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_215),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_14),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_208),
.B(n_198),
.CI(n_192),
.CON(n_220),
.SN(n_220)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_221),
.B(n_222),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_196),
.CI(n_205),
.CON(n_222),
.SN(n_222)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_227),
.C(n_229),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_201),
.B1(n_188),
.B2(n_202),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_228),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_199),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_238),
.Y(n_240)
);

OA21x2_ASAP7_75t_SL g237 ( 
.A1(n_229),
.A2(n_209),
.B(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_225),
.A2(n_213),
.B(n_219),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_226),
.Y(n_239)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_243),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_224),
.B(n_238),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_221),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_242),
.B(n_231),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_249),
.A3(n_240),
.B1(n_222),
.B2(n_220),
.C1(n_227),
.C2(n_10),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_5),
.B(n_7),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_232),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_250),
.A2(n_252),
.A3(n_248),
.B1(n_247),
.B2(n_10),
.C1(n_11),
.C2(n_8),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_253),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_254),
.B1(n_9),
.B2(n_12),
.Y(n_256)
);

XNOR2x2_ASAP7_75t_SL g257 ( 
.A(n_256),
.B(n_9),
.Y(n_257)
);


endmodule