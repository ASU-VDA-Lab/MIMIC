module fake_jpeg_7449_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_26),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_31),
.B1(n_29),
.B2(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_46),
.A2(n_17),
.B1(n_33),
.B2(n_22),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_29),
.B1(n_31),
.B2(n_16),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_21),
.B1(n_42),
.B2(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_60),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_22),
.B(n_33),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_32),
.B1(n_26),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_43),
.B1(n_18),
.B2(n_22),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_23),
.B1(n_28),
.B2(n_42),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_67),
.B1(n_50),
.B2(n_42),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_68),
.A2(n_57),
.B1(n_64),
.B2(n_59),
.Y(n_113)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_77),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_36),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_82),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_87),
.B1(n_33),
.B2(n_16),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_17),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_36),
.Y(n_91)
);

NOR2x1_ASAP7_75t_R g92 ( 
.A(n_81),
.B(n_78),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_93),
.B(n_37),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_40),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_94),
.A2(n_88),
.B1(n_89),
.B2(n_30),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_40),
.C(n_41),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_116),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_23),
.B1(n_28),
.B2(n_42),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_102),
.B1(n_74),
.B2(n_77),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_98),
.A2(n_30),
.B1(n_19),
.B2(n_15),
.Y(n_147)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_109),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_108),
.B(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_36),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_87),
.B1(n_83),
.B2(n_74),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_118),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_82),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_71),
.B1(n_72),
.B2(n_68),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_125),
.B1(n_130),
.B2(n_138),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_128),
.B1(n_133),
.B2(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_123),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_126),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_67),
.B1(n_38),
.B2(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_127),
.B(n_135),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_38),
.B1(n_69),
.B2(n_77),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_75),
.A3(n_90),
.B1(n_85),
.B2(n_74),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_132),
.B(n_118),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_77),
.B1(n_69),
.B2(n_59),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_76),
.A3(n_19),
.B1(n_37),
.B2(n_41),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_141),
.B1(n_146),
.B2(n_117),
.Y(n_158)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_114),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_38),
.B1(n_69),
.B2(n_53),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_99),
.B1(n_105),
.B2(n_113),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_108),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_69),
.B1(n_45),
.B2(n_41),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_93),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_110),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_37),
.B1(n_36),
.B2(n_21),
.Y(n_143)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_155),
.B(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_159),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_166),
.B1(n_178),
.B2(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_161),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_93),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_175),
.C(n_177),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_20),
.B1(n_84),
.B2(n_24),
.Y(n_195)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_167),
.Y(n_200)
);

AO21x2_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_95),
.B(n_100),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_112),
.B1(n_37),
.B2(n_100),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_124),
.B(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_136),
.B(n_12),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_131),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_107),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_107),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_20),
.B(n_37),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_0),
.B(n_1),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_49),
.C(n_37),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_141),
.C(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_20),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_177),
.C(n_174),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_192),
.C(n_203),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_190),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_187),
.A2(n_191),
.B1(n_197),
.B2(n_171),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

XOR2x2_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_147),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_13),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_164),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_127),
.B1(n_128),
.B2(n_135),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_146),
.C(n_84),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_165),
.B1(n_178),
.B2(n_148),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_84),
.B1(n_27),
.B2(n_24),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_202),
.B(n_169),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_R g202 ( 
.A(n_166),
.B(n_14),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_15),
.Y(n_203)
);

XOR2x2_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_14),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_204),
.A2(n_157),
.B(n_172),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_14),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_163),
.C(n_155),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_0),
.Y(n_226)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_207),
.B(n_162),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_205),
.C(n_186),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_218),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_193),
.C(n_183),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_214),
.C(n_217),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_160),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_225),
.B1(n_233),
.B2(n_199),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_160),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_219),
.A2(n_220),
.B(n_224),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_150),
.C(n_179),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_223),
.C(n_196),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_156),
.C(n_167),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_167),
.B1(n_153),
.B2(n_161),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_182),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_232),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_230),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_13),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_189),
.A2(n_13),
.B(n_12),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_194),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_184),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_203),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_238),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_184),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_204),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_220),
.B1(n_230),
.B2(n_228),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_191),
.B1(n_200),
.B2(n_187),
.Y(n_242)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_250),
.C(n_251),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_197),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_221),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_252),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_201),
.C(n_196),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_12),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_234),
.C(n_237),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_262),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_222),
.B1(n_225),
.B2(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_211),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_265),
.Y(n_275)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_267),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_219),
.C(n_233),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_269),
.C(n_270),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_1),
.C(n_3),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_251),
.C(n_250),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_281),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_235),
.C(n_246),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_10),
.C(n_9),
.Y(n_289)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_257),
.B(n_253),
.CI(n_240),
.CON(n_279),
.SN(n_279)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_283),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_253),
.B(n_244),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_9),
.Y(n_290)
);

AO22x1_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_240),
.B1(n_234),
.B2(n_5),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_262),
.B1(n_267),
.B2(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_260),
.CI(n_11),
.CON(n_283),
.SN(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_260),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_287),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_10),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_294),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_278),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_6),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_1),
.C(n_3),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_296),
.B(n_284),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_9),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_279),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_3),
.C(n_5),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_302),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_305),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_277),
.Y(n_302)
);

NOR2x1_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_281),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_304),
.B1(n_295),
.B2(n_291),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_271),
.B1(n_279),
.B2(n_283),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_310),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_293),
.B(n_285),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_307),
.A2(n_308),
.B(n_298),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_296),
.B(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_298),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_314),
.B(n_308),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_313),
.B(n_309),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_277),
.C(n_7),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_7),
.C(n_8),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_7),
.Y(n_320)
);


endmodule