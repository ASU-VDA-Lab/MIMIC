module real_jpeg_2045_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_285, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_285;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_1),
.A2(n_74),
.B1(n_75),
.B2(n_81),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_1),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_81),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_81),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_81),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_3),
.A2(n_36),
.B1(n_74),
.B2(n_75),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_3),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_3),
.A2(n_36),
.B1(n_64),
.B2(n_65),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_74),
.B1(n_75),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_4),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_135),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_135),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_135),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_5),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_127)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_40),
.B1(n_64),
.B2(n_65),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_10),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_40),
.B1(n_74),
.B2(n_75),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_12),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_13),
.A2(n_74),
.B1(n_75),
.B2(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_13),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_164),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_164),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_164),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_14),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_14),
.B(n_83),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_14),
.B(n_64),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_14),
.A2(n_74),
.B(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_14),
.B(n_33),
.C(n_49),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_155),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_14),
.B(n_111),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_14),
.B(n_29),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_14),
.B(n_57),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g254 ( 
.A1(n_14),
.A2(n_64),
.B(n_188),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_20),
.B(n_114),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_86),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.C(n_71),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_24),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_25),
.A2(n_26),
.B1(n_42),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_27),
.A2(n_41),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_33),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_28),
.A2(n_31),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_28),
.A2(n_38),
.B(n_152),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_28),
.A2(n_91),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_29),
.B(n_39),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_29),
.A2(n_41),
.B1(n_127),
.B2(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_29),
.A2(n_41),
.B1(n_155),
.B2(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_29),
.A2(n_41),
.B1(n_235),
.B2(n_238),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_31),
.A2(n_91),
.B(n_128),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_33),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_33),
.B(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_42),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_43),
.A2(n_54),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_43),
.A2(n_93),
.B(n_106),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_43),
.A2(n_56),
.B1(n_184),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_44),
.B(n_94),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_44),
.A2(n_105),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_44),
.A2(n_57),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_44),
.A2(n_57),
.B1(n_221),
.B2(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_46),
.B(n_60),
.C(n_65),
.Y(n_189)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_47),
.A2(n_61),
.B(n_187),
.C(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_47),
.B(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_52),
.A2(n_56),
.B(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_57),
.B(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_58),
.B(n_71),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B(n_66),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_59),
.A2(n_69),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_59),
.A2(n_69),
.B1(n_175),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_70)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_63),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_65),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_64),
.B(n_75),
.C(n_78),
.Y(n_156)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_65),
.A2(n_77),
.B(n_154),
.C(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_67),
.B(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_68),
.A2(n_111),
.B1(n_159),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_69),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_69),
.A2(n_158),
.B(n_160),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_80),
.B(n_82),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_79),
.B1(n_80),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_72),
.A2(n_79),
.B1(n_134),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_72),
.A2(n_79),
.B1(n_163),
.B2(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_79),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_75),
.B(n_155),
.Y(n_154)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_101),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_102),
.B2(n_103),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_95),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_92),
.B1(n_96),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_126),
.B(n_128),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_109),
.B(n_113),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_111),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_121),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_122),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.C(n_133),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_124),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_125),
.B(n_129),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_133),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_169),
.B(n_283),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_165),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_140),
.B(n_165),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_146),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_141),
.B(n_144),
.Y(n_266)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_146),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_157),
.C(n_162),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_147),
.A2(n_148),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_157),
.B(n_162),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI321xp33_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_264),
.A3(n_275),
.B1(n_281),
.B2(n_282),
.C(n_285),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_210),
.B(n_263),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_191),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_172),
.B(n_191),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_182),
.C(n_185),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_173),
.B(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_178),
.C(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_182),
.B(n_185),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_190),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_203),
.B2(n_204),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_192),
.B(n_205),
.C(n_208),
.Y(n_276)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_194),
.B(n_198),
.C(n_202),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_258),
.B(n_262),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_248),
.B(n_257),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_229),
.B(n_247),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_226),
.C(n_228),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_241),
.B(n_246),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_236),
.B(n_240),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_239),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_245),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_250),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_253),
.C(n_255),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_267),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.C(n_274),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_269),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);


endmodule