module fake_ariane_840_n_1926 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1926);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1926;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_16),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_1),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_49),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_89),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_19),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_73),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_150),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_99),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_69),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_60),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_83),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_58),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_163),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_79),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_28),
.Y(n_204)
);

INVxp33_ASAP7_75t_R g205 ( 
.A(n_37),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_147),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_135),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_64),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_32),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_75),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_61),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_2),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_95),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_26),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_71),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_15),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_103),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_48),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_19),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_175),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_148),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_0),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_166),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_15),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_31),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_156),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_169),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_171),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_61),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_106),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_114),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_57),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_21),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_167),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_58),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_60),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_104),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_100),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_77),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_45),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_66),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_118),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_102),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_76),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_90),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_68),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_158),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_52),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_180),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_26),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_32),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_50),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_98),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_40),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_128),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_37),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_3),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_172),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_139),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_109),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_112),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_134),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_111),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_161),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_130),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_145),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_93),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_125),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_153),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_45),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_17),
.Y(n_279)
);

BUFx8_ASAP7_75t_SL g280 ( 
.A(n_23),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_140),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_85),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_17),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_84),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_162),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_40),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_30),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_124),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_108),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_21),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_74),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_157),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_55),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_91),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_119),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_54),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_126),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_80),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_30),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_160),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_8),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_170),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_53),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_55),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_35),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_136),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_51),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_0),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_52),
.Y(n_309)
);

BUFx10_ASAP7_75t_L g310 ( 
.A(n_38),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_1),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_87),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_48),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_129),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_94),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_137),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_27),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_24),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_63),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_168),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_115),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_144),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_101),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_78),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_152),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_63),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_36),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_178),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_25),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_113),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_96),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_3),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_110),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_23),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_92),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_121),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_47),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_7),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_29),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_81),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_105),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_49),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_29),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_82),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_116),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_44),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_44),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_176),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_6),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_11),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_138),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_22),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_173),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_131),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_164),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_9),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_88),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_43),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_59),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_39),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_127),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_177),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_308),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_234),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_234),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_230),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_280),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_215),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_226),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_234),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_235),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_286),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_308),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_243),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_254),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_276),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_206),
.B(n_231),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_234),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_234),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_246),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_240),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_246),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_335),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_278),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_344),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_361),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_278),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_356),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_223),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_273),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_273),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_190),
.B(n_181),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_224),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_287),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_182),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_293),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_305),
.B(n_4),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_227),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_311),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_229),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_295),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_237),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_241),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_240),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_295),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_189),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_302),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_186),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_182),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_302),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_242),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_240),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_257),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_251),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_183),
.B(n_4),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_354),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_310),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_198),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_194),
.B(n_5),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_258),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_251),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_259),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_251),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_252),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_261),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_219),
.B(n_5),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_252),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_209),
.B(n_6),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_218),
.B(n_8),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_186),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_263),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_183),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_238),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_264),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_310),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_255),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_268),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_303),
.Y(n_440)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_184),
.B(n_9),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_313),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_317),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_318),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_279),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_222),
.B(n_10),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_283),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_326),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_310),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_296),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_329),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_239),
.B(n_10),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_334),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_338),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_375),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_376),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_383),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_364),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_364),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_363),
.B(n_252),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_395),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_373),
.B(n_260),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_185),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_365),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_397),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_386),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_369),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_365),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_400),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_371),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_370),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_378),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_409),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_374),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_385),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_367),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_389),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_378),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_368),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_394),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_399),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_381),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_381),
.B(n_266),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_405),
.Y(n_487)
);

NAND2x1_ASAP7_75t_L g488 ( 
.A(n_391),
.B(n_185),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g490 ( 
.A(n_372),
.B(n_184),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_401),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_403),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_430),
.A2(n_282),
.B(n_267),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_409),
.B(n_285),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_404),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_412),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_413),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_408),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_407),
.B(n_438),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_408),
.B(n_193),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_434),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_411),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_377),
.B(n_294),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_414),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_453),
.B(n_266),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_417),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_415),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_L g516 ( 
.A(n_417),
.B(n_220),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_419),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_419),
.Y(n_518)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_380),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_380),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_382),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_382),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_384),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_384),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_387),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_423),
.B(n_266),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_387),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_420),
.B(n_275),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_434),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_388),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_388),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_390),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_474),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_459),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_459),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_478),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_482),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_507),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_529),
.B(n_422),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_529),
.B(n_435),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_458),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_458),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_474),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_507),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_459),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_472),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_459),
.Y(n_548)
);

BUFx4f_ASAP7_75t_L g549 ( 
.A(n_507),
.Y(n_549)
);

AND3x1_ASAP7_75t_L g550 ( 
.A(n_510),
.B(n_431),
.C(n_421),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g551 ( 
.A(n_460),
.B(n_193),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_507),
.A2(n_393),
.B1(n_446),
.B2(n_366),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_505),
.B(n_435),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_461),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_472),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_505),
.B(n_439),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_499),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_479),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_465),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_507),
.A2(n_452),
.B1(n_428),
.B2(n_410),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_455),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_479),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_460),
.B(n_424),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_474),
.B(n_418),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_520),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_483),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_499),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_473),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_512),
.B(n_508),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_508),
.B(n_427),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_469),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_473),
.Y(n_572)
);

AND3x2_ASAP7_75t_L g573 ( 
.A(n_486),
.B(n_449),
.C(n_437),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_483),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_481),
.B(n_396),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_SL g578 ( 
.A(n_484),
.B(n_491),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_506),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_507),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_468),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_468),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_507),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_SL g584 ( 
.A(n_494),
.B(n_433),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_506),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_L g586 ( 
.A1(n_527),
.A2(n_290),
.B1(n_221),
.B2(n_217),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_499),
.Y(n_587)
);

INVxp67_ASAP7_75t_SL g588 ( 
.A(n_506),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_499),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_519),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_470),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_498),
.B(n_436),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_499),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_500),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_512),
.B(n_439),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_508),
.B(n_530),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_519),
.A2(n_301),
.B1(n_416),
.B2(n_441),
.Y(n_597)
);

BUFx6f_ASAP7_75t_SL g598 ( 
.A(n_485),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_488),
.B(n_428),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_508),
.B(n_440),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_511),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_499),
.Y(n_602)
);

OR2x6_ASAP7_75t_L g603 ( 
.A(n_488),
.B(n_454),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_462),
.B(n_445),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_470),
.Y(n_606)
);

BUFx4f_ASAP7_75t_L g607 ( 
.A(n_520),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_530),
.B(n_447),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_519),
.Y(n_609)
);

INVx4_ASAP7_75t_SL g610 ( 
.A(n_519),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_464),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_530),
.B(n_440),
.Y(n_612)
);

INVx6_ASAP7_75t_L g613 ( 
.A(n_530),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_475),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_456),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_480),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_480),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_520),
.A2(n_343),
.B1(n_359),
.B2(n_426),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_457),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_502),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_464),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_497),
.B(n_450),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_464),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_490),
.B(n_187),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_502),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_516),
.B(n_442),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_516),
.B(n_442),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_502),
.B(n_443),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_509),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_509),
.Y(n_631)
);

AND2x6_ASAP7_75t_L g632 ( 
.A(n_509),
.B(n_197),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_489),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_464),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_464),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_464),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_520),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_463),
.B(n_443),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_521),
.B(n_522),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_520),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_489),
.B(n_425),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_466),
.B(n_187),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_492),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_463),
.B(n_444),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_467),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_520),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_492),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_526),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_L g649 ( 
.A(n_526),
.B(n_277),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_471),
.B(n_476),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_493),
.B(n_444),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_521),
.B(n_448),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_526),
.Y(n_653)
);

BUFx4f_ASAP7_75t_L g654 ( 
.A(n_526),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_493),
.B(n_429),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_526),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_496),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_496),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_503),
.B(n_448),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_L g660 ( 
.A(n_526),
.B(n_277),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_503),
.B(n_451),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_504),
.A2(n_349),
.B1(n_337),
.B2(n_339),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_504),
.B(n_451),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_495),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_531),
.B(n_188),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_531),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_513),
.B(n_454),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_513),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_514),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_487),
.Y(n_670)
);

INVx4_ASAP7_75t_SL g671 ( 
.A(n_531),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_514),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_531),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_522),
.B(n_390),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_531),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_523),
.B(n_398),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_517),
.B(n_518),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_531),
.A2(n_314),
.B1(n_275),
.B2(n_271),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_517),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_532),
.Y(n_680)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_518),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_551),
.A2(n_524),
.B1(n_525),
.B2(n_528),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_538),
.B(n_501),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_680),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_577),
.Y(n_685)
);

INVx8_ASAP7_75t_L g686 ( 
.A(n_639),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_680),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_664),
.A2(n_495),
.B(n_523),
.Y(n_688)
);

INVx8_ASAP7_75t_L g689 ( 
.A(n_639),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_538),
.B(n_515),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_680),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_542),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_581),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_623),
.B(n_528),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_563),
.B(n_205),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_664),
.B(n_277),
.Y(n_696)
);

INVxp67_ASAP7_75t_SL g697 ( 
.A(n_579),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_540),
.B(n_200),
.Y(n_698)
);

BUFx6f_ASAP7_75t_SL g699 ( 
.A(n_645),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_541),
.B(n_533),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_592),
.B(n_277),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_545),
.B(n_188),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_542),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_554),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_581),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_551),
.A2(n_525),
.B1(n_524),
.B2(n_533),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_582),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_582),
.Y(n_708)
);

AND2x6_ASAP7_75t_SL g709 ( 
.A(n_641),
.B(n_398),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_543),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_541),
.B(n_532),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_639),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_627),
.B(n_628),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_639),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_543),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_550),
.A2(n_216),
.B1(n_213),
.B2(n_357),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_545),
.B(n_191),
.Y(n_717)
);

BUFx12f_ASAP7_75t_L g718 ( 
.A(n_645),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_604),
.B(n_200),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_577),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_627),
.B(n_532),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_547),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_591),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_604),
.B(n_204),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_655),
.B(n_204),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_592),
.B(n_211),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_547),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_545),
.B(n_191),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_555),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_555),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_550),
.A2(n_360),
.B1(n_358),
.B2(n_211),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_L g732 ( 
.A(n_552),
.B(n_337),
.C(n_214),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_627),
.B(n_192),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_642),
.B(n_564),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_564),
.B(n_214),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_SL g736 ( 
.A(n_594),
.B(n_339),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_627),
.B(n_628),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_628),
.B(n_195),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_628),
.B(n_195),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_616),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_564),
.B(n_342),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_558),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_558),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_617),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_617),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_681),
.B(n_196),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_595),
.B(n_196),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_562),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_SL g749 ( 
.A(n_561),
.B(n_275),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_562),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_553),
.B(n_297),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_535),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_551),
.A2(n_357),
.B1(n_201),
.B2(n_353),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_595),
.B(n_199),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_566),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_583),
.B(n_199),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_633),
.A2(n_342),
.B1(n_360),
.B2(n_358),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_553),
.B(n_201),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_559),
.B(n_346),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_535),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_618),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_549),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_594),
.B(n_346),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_536),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_583),
.B(n_202),
.Y(n_765)
);

AND2x4_ASAP7_75t_SL g766 ( 
.A(n_605),
.B(n_314),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_551),
.A2(n_314),
.B1(n_347),
.B2(n_352),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_551),
.A2(n_556),
.B1(n_612),
.B2(n_600),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_605),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_566),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_537),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_633),
.A2(n_350),
.B1(n_347),
.B2(n_349),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_564),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_573),
.Y(n_774)
);

NOR2xp67_ASAP7_75t_L g775 ( 
.A(n_650),
.B(n_202),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_571),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_584),
.B(n_578),
.C(n_662),
.Y(n_777)
);

AND2x4_ASAP7_75t_SL g778 ( 
.A(n_605),
.B(n_537),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_583),
.B(n_203),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_679),
.A2(n_569),
.B1(n_621),
.B2(n_618),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_551),
.A2(n_350),
.B1(n_352),
.B2(n_316),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_556),
.A2(n_312),
.B(n_355),
.C(n_322),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_600),
.B(n_203),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_551),
.A2(n_353),
.B1(n_208),
.B2(n_348),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_679),
.A2(n_351),
.B1(n_324),
.B2(n_325),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_536),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_546),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_612),
.B(n_207),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_575),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_570),
.B(n_207),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_546),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_625),
.B(n_299),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_549),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_629),
.A2(n_340),
.B(n_330),
.C(n_309),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_548),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_548),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_618),
.B(n_210),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_568),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_621),
.B(n_210),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_621),
.B(n_212),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_575),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_631),
.B(n_212),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_631),
.B(n_213),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_601),
.B(n_327),
.C(n_304),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_586),
.B(n_307),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_615),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_643),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_650),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_590),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_603),
.B(n_11),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_643),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_601),
.B(n_319),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_568),
.Y(n_813)
);

AOI221xp5_ASAP7_75t_L g814 ( 
.A1(n_662),
.A2(n_332),
.B1(n_348),
.B2(n_345),
.C(n_341),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_677),
.B(n_272),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_SL g816 ( 
.A(n_615),
.B(n_272),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_659),
.B(n_336),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_590),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_626),
.A2(n_341),
.B(n_345),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_647),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_565),
.B(n_666),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_661),
.B(n_225),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_630),
.B(n_228),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_614),
.B(n_12),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_537),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_630),
.B(n_232),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_646),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_572),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_647),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_657),
.B(n_233),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_572),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_574),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_657),
.A2(n_362),
.B(n_333),
.C(n_331),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_620),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_658),
.B(n_236),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_658),
.A2(n_328),
.B(n_323),
.C(n_321),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_565),
.B(n_277),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_565),
.B(n_277),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_574),
.Y(n_839)
);

OAI22xp33_ASAP7_75t_L g840 ( 
.A1(n_597),
.A2(n_320),
.B1(n_315),
.B2(n_306),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_560),
.A2(n_300),
.B1(n_298),
.B2(n_292),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_565),
.B(n_277),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_670),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_676),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_626),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_668),
.B(n_291),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_694),
.B(n_652),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_692),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_714),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_725),
.B(n_608),
.C(n_667),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_703),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_710),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_810),
.A2(n_672),
.B1(n_668),
.B2(n_669),
.Y(n_853)
);

AO21x1_ASAP7_75t_L g854 ( 
.A1(n_696),
.A2(n_669),
.B(n_672),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_714),
.B(n_620),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_696),
.A2(n_576),
.B(n_654),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_688),
.A2(n_576),
.B(n_587),
.Y(n_857)
);

AOI21x1_ASAP7_75t_L g858 ( 
.A1(n_821),
.A2(n_587),
.B(n_593),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_685),
.B(n_720),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_780),
.A2(n_821),
.B(n_799),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_719),
.B(n_674),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_724),
.B(n_674),
.Y(n_862)
);

BUFx4f_ASAP7_75t_L g863 ( 
.A(n_718),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_715),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_806),
.B(n_620),
.Y(n_865)
);

AO32x1_ASAP7_75t_L g866 ( 
.A1(n_722),
.A2(n_606),
.A3(n_675),
.B1(n_673),
.B2(n_648),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_727),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_731),
.A2(n_663),
.B(n_651),
.C(n_665),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_698),
.B(n_619),
.Y(n_869)
);

BUFx12f_ASAP7_75t_L g870 ( 
.A(n_718),
.Y(n_870)
);

BUFx4f_ASAP7_75t_L g871 ( 
.A(n_778),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_799),
.A2(n_607),
.B(n_654),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_761),
.A2(n_607),
.B(n_654),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_776),
.Y(n_874)
);

OAI21xp33_ASAP7_75t_L g875 ( 
.A1(n_816),
.A2(n_597),
.B(n_678),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_761),
.A2(n_607),
.B(n_588),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_805),
.A2(n_676),
.B1(n_599),
.B2(n_606),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_700),
.B(n_603),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_726),
.B(n_603),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_729),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_702),
.A2(n_596),
.B(n_637),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_695),
.B(n_645),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_730),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_843),
.B(n_598),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_704),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_714),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_742),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_845),
.Y(n_888)
);

AO21x1_ASAP7_75t_L g889 ( 
.A1(n_701),
.A2(n_649),
.B(n_660),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_717),
.A2(n_567),
.B(n_640),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_734),
.B(n_598),
.Y(n_891)
);

NOR2x1_ASAP7_75t_L g892 ( 
.A(n_777),
.B(n_534),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_728),
.A2(n_602),
.B(n_637),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_815),
.A2(n_603),
.B(n_602),
.C(n_557),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_751),
.B(n_534),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_728),
.A2(n_602),
.B(n_557),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_751),
.B(n_544),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_686),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_756),
.A2(n_779),
.B(n_765),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_751),
.B(n_544),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_773),
.B(n_579),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_743),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_845),
.A2(n_593),
.B(n_673),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_758),
.A2(n_656),
.B(n_589),
.C(n_644),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_778),
.B(n_610),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_714),
.B(n_609),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_SL g907 ( 
.A(n_814),
.B(n_638),
.C(n_244),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_810),
.A2(n_599),
.B1(n_656),
.B2(n_609),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_747),
.A2(n_599),
.B(n_635),
.C(n_611),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_L g910 ( 
.A(n_749),
.B(n_609),
.C(n_646),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_810),
.A2(n_599),
.B1(n_646),
.B2(n_611),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_779),
.A2(n_611),
.B(n_635),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_797),
.A2(n_635),
.B(n_675),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_768),
.A2(n_648),
.B(n_653),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_800),
.A2(n_653),
.B(n_580),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_773),
.B(n_585),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_802),
.A2(n_539),
.B(n_580),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_808),
.B(n_598),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_686),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_686),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_776),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_803),
.A2(n_539),
.B(n_580),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_712),
.B(n_666),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_733),
.B(n_585),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_754),
.A2(n_649),
.B(n_660),
.C(n_634),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_844),
.B(n_666),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_771),
.B(n_834),
.Y(n_927)
);

AO21x1_ASAP7_75t_L g928 ( 
.A1(n_701),
.A2(n_622),
.B(n_624),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_817),
.B(n_711),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_752),
.A2(n_539),
.B(n_636),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_713),
.B(n_666),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_748),
.A2(n_634),
.B1(n_624),
.B2(n_613),
.Y(n_932)
);

AO32x1_ASAP7_75t_L g933 ( 
.A1(n_750),
.A2(n_632),
.A3(n_671),
.B1(n_14),
.B2(n_16),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_760),
.A2(n_269),
.B(n_245),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_760),
.A2(n_270),
.B(n_247),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_763),
.B(n_610),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_737),
.A2(n_613),
.B1(n_610),
.B2(n_671),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_764),
.A2(n_274),
.B(n_248),
.Y(n_938)
);

INVx4_ASAP7_75t_L g939 ( 
.A(n_686),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_683),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_771),
.B(n_613),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_764),
.A2(n_281),
.B(n_249),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_834),
.B(n_613),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_712),
.B(n_689),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_689),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_786),
.A2(n_632),
.B(n_284),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_689),
.A2(n_610),
.B1(n_671),
.B2(n_632),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_689),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_755),
.B(n_770),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_833),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_789),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_736),
.B(n_671),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_801),
.B(n_807),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_774),
.B(n_289),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_L g955 ( 
.A(n_736),
.B(n_690),
.C(n_804),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_812),
.B(n_288),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_786),
.A2(n_265),
.B(n_256),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_766),
.B(n_253),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_769),
.B(n_250),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_787),
.A2(n_262),
.B(n_197),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_769),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_811),
.B(n_632),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_787),
.A2(n_262),
.B(n_197),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_820),
.B(n_632),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_790),
.A2(n_632),
.B(n_18),
.C(n_20),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_791),
.A2(n_262),
.B(n_197),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_829),
.B(n_632),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_825),
.B(n_262),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_833),
.A2(n_836),
.B(n_782),
.C(n_746),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_836),
.A2(n_13),
.B(n_18),
.C(n_22),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_782),
.A2(n_735),
.B(n_741),
.C(n_772),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_766),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_732),
.A2(n_197),
.B1(n_27),
.B2(n_28),
.Y(n_973)
);

CKINVDCx10_ASAP7_75t_R g974 ( 
.A(n_699),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_759),
.B(n_24),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_809),
.B(n_818),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_716),
.B(n_31),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_822),
.B(n_33),
.Y(n_978)
);

AND2x2_ASAP7_75t_SL g979 ( 
.A(n_767),
.B(n_33),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_721),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_980)
);

AND2x2_ASAP7_75t_SL g981 ( 
.A(n_781),
.B(n_34),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_809),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_818),
.Y(n_983)
);

AND2x2_ASAP7_75t_SL g984 ( 
.A(n_753),
.B(n_784),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_697),
.B(n_38),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_824),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_762),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_738),
.B(n_739),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_795),
.A2(n_65),
.B(n_165),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_783),
.B(n_41),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_840),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_795),
.A2(n_42),
.B(n_46),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_792),
.A2(n_46),
.B(n_47),
.C(n_50),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_682),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_796),
.A2(n_86),
.B(n_146),
.Y(n_995)
);

BUFx4f_ASAP7_75t_L g996 ( 
.A(n_699),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_706),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_796),
.A2(n_97),
.B(n_141),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_788),
.B(n_56),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_798),
.A2(n_123),
.B(n_67),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_757),
.A2(n_62),
.B(n_70),
.C(n_72),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_813),
.A2(n_831),
.B(n_832),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_775),
.B(n_62),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_823),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_828),
.A2(n_832),
.B(n_831),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_L g1006 ( 
.A(n_826),
.B(n_846),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_839),
.A2(n_684),
.B(n_687),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_830),
.A2(n_835),
.B(n_839),
.C(n_794),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_684),
.A2(n_687),
.B(n_691),
.C(n_841),
.Y(n_1009)
);

NOR2xp67_ASAP7_75t_L g1010 ( 
.A(n_819),
.B(n_785),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_693),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_709),
.B(n_699),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_693),
.B(n_705),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_705),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_762),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_827),
.A2(n_707),
.B(n_708),
.C(n_723),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_708),
.B(n_723),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_837),
.A2(n_842),
.B(n_838),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_762),
.B(n_793),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_929),
.A2(n_838),
.B(n_793),
.Y(n_1020)
);

O2A1O1Ixp5_ASAP7_75t_L g1021 ( 
.A1(n_854),
.A2(n_740),
.B(n_744),
.C(n_745),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_857),
.A2(n_745),
.B(n_762),
.Y(n_1022)
);

AOI221x1_ASAP7_75t_L g1023 ( 
.A1(n_977),
.A2(n_793),
.B1(n_899),
.B2(n_992),
.C(n_853),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_847),
.B(n_861),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_956),
.A2(n_862),
.B(n_975),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_853),
.A2(n_856),
.B(n_879),
.Y(n_1026)
);

AO21x2_ASAP7_75t_L g1027 ( 
.A1(n_1016),
.A2(n_903),
.B(n_914),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_848),
.Y(n_1028)
);

NAND2x1p5_ASAP7_75t_L g1029 ( 
.A(n_898),
.B(n_920),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_948),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_898),
.B(n_920),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_984),
.B(n_911),
.Y(n_1032)
);

BUFx4_ASAP7_75t_SL g1033 ( 
.A(n_874),
.Y(n_1033)
);

AO31x2_ASAP7_75t_L g1034 ( 
.A1(n_889),
.A2(n_1018),
.A3(n_1002),
.B(n_1005),
.Y(n_1034)
);

NOR2x1_ASAP7_75t_SL g1035 ( 
.A(n_939),
.B(n_1015),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_988),
.A2(n_903),
.B(n_1008),
.Y(n_1036)
);

CKINVDCx11_ASAP7_75t_R g1037 ( 
.A(n_870),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_948),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_969),
.A2(n_878),
.B(n_1007),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_913),
.A2(n_1007),
.B(n_915),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_921),
.B(n_939),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_859),
.B(n_882),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_949),
.A2(n_953),
.B1(n_869),
.B2(n_971),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_948),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_926),
.B(n_877),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1006),
.A2(n_978),
.B(n_894),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_904),
.A2(n_909),
.B(n_872),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_851),
.B(n_852),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_932),
.A2(n_892),
.B(n_881),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_864),
.B(n_867),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_880),
.B(n_883),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_873),
.A2(n_876),
.B(n_896),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_885),
.B(n_940),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_890),
.A2(n_893),
.B(n_912),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_930),
.A2(n_917),
.B(n_922),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_887),
.B(n_902),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_911),
.B(n_908),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_951),
.B(n_865),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_875),
.B(n_891),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_SL g1060 ( 
.A(n_1015),
.B(n_908),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_990),
.A2(n_999),
.B(n_952),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_986),
.B(n_927),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_919),
.Y(n_1063)
);

AND2x6_ASAP7_75t_L g1064 ( 
.A(n_947),
.B(n_919),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_871),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_976),
.B(n_1004),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_1013),
.A2(n_960),
.B(n_966),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_868),
.A2(n_931),
.B(n_925),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_963),
.A2(n_1019),
.B(n_989),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_945),
.B(n_976),
.Y(n_1070)
);

AND2x6_ASAP7_75t_L g1071 ( 
.A(n_945),
.B(n_1015),
.Y(n_1071)
);

CKINVDCx6p67_ASAP7_75t_R g1072 ( 
.A(n_974),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_995),
.A2(n_1000),
.B(n_998),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_850),
.A2(n_866),
.B(n_964),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_941),
.B(n_943),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_992),
.A2(n_979),
.B(n_981),
.C(n_993),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_905),
.B(n_961),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_888),
.A2(n_967),
.B(n_962),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_987),
.B(n_1010),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_895),
.B(n_900),
.Y(n_1080)
);

AO21x1_ASAP7_75t_L g1081 ( 
.A1(n_1001),
.A2(n_950),
.B(n_970),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_972),
.B(n_918),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1014),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_897),
.B(n_958),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_946),
.A2(n_923),
.B(n_987),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_991),
.A2(n_980),
.B1(n_985),
.B2(n_994),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_849),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_866),
.A2(n_1003),
.B(n_924),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_866),
.A2(n_933),
.B(n_938),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1017),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_936),
.B(n_954),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_884),
.B(n_1012),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_849),
.B(n_886),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_955),
.B(n_961),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_907),
.A2(n_944),
.B1(n_997),
.B2(n_994),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_L g1096 ( 
.A1(n_968),
.A2(n_906),
.B(n_934),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_871),
.B(n_863),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_863),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_933),
.A2(n_942),
.B(n_935),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_855),
.A2(n_901),
.B(n_916),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_996),
.B(n_983),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_SL g1102 ( 
.A1(n_997),
.A2(n_973),
.B(n_957),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_910),
.A2(n_905),
.B1(n_983),
.B2(n_982),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_982),
.B(n_983),
.Y(n_1104)
);

AOI21xp33_ASAP7_75t_L g1105 ( 
.A1(n_959),
.A2(n_937),
.B(n_982),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_849),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_886),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_933),
.A2(n_965),
.B(n_886),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_996),
.A2(n_854),
.A3(n_928),
.B(n_1016),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_861),
.A2(n_862),
.B(n_977),
.C(n_725),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_854),
.A2(n_928),
.A3(n_1016),
.B(n_1009),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_859),
.B(n_685),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_977),
.A2(n_971),
.B(n_869),
.C(n_992),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_929),
.A2(n_847),
.B(n_696),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_929),
.A2(n_847),
.B(n_696),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_859),
.B(n_685),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_SL g1117 ( 
.A1(n_854),
.A2(n_992),
.B(n_853),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_847),
.B(n_861),
.Y(n_1118)
);

NAND2x1_ASAP7_75t_L g1119 ( 
.A(n_987),
.B(n_712),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_977),
.A2(n_971),
.B(n_869),
.C(n_992),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_847),
.B(n_861),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_847),
.B(n_861),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_848),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_929),
.A2(n_847),
.B(n_696),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_874),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_859),
.B(n_685),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_857),
.A2(n_688),
.B(n_858),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_848),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_859),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_847),
.A2(n_853),
.B1(n_862),
.B2(n_861),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_859),
.B(n_685),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_854),
.A2(n_928),
.A3(n_1016),
.B(n_1009),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_859),
.B(n_685),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_929),
.A2(n_1009),
.B(n_988),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_898),
.B(n_939),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_874),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_977),
.A2(n_971),
.B(n_869),
.C(n_992),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_848),
.Y(n_1138)
);

AOI221x1_ASAP7_75t_L g1139 ( 
.A1(n_977),
.A2(n_899),
.B1(n_860),
.B2(n_992),
.C(n_853),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_857),
.A2(n_688),
.B(n_858),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_929),
.A2(n_847),
.B(n_696),
.Y(n_1141)
);

NAND2x1p5_ASAP7_75t_L g1142 ( 
.A(n_898),
.B(n_939),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_859),
.B(n_685),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_848),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_848),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_929),
.A2(n_847),
.B(n_696),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_859),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1011),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_847),
.B(n_861),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_857),
.A2(n_688),
.B(n_858),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_847),
.B(n_861),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_929),
.A2(n_847),
.B(n_696),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_857),
.A2(n_688),
.B(n_858),
.Y(n_1153)
);

AOI21x1_ASAP7_75t_L g1154 ( 
.A1(n_860),
.A2(n_854),
.B(n_928),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_857),
.A2(n_688),
.B(n_858),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_847),
.B(n_844),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_879),
.B(n_714),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_848),
.Y(n_1158)
);

NAND2xp33_ASAP7_75t_SL g1159 ( 
.A(n_853),
.B(n_714),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_859),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_888),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_874),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_847),
.B(n_861),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_871),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1028),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1156),
.B(n_1112),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1025),
.A2(n_1110),
.B(n_1113),
.C(n_1137),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1077),
.Y(n_1168)
);

OAI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1042),
.A2(n_1095),
.B1(n_1163),
.B2(n_1118),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1114),
.A2(n_1124),
.B(n_1115),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1077),
.B(n_1097),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1156),
.B(n_1024),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1033),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1087),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1059),
.A2(n_1032),
.B1(n_1086),
.B2(n_1159),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1114),
.A2(n_1124),
.B(n_1115),
.Y(n_1176)
);

NAND2x1p5_ASAP7_75t_L g1177 ( 
.A(n_1101),
.B(n_1070),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1129),
.B(n_1147),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_1037),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1113),
.A2(n_1137),
.B(n_1120),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1116),
.B(n_1126),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1059),
.A2(n_1032),
.B1(n_1159),
.B2(n_1045),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1110),
.A2(n_1120),
.B(n_1130),
.C(n_1076),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1123),
.Y(n_1185)
);

BUFx4f_ASAP7_75t_SL g1186 ( 
.A(n_1072),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1143),
.B(n_1129),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1121),
.B(n_1122),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1029),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1033),
.Y(n_1190)
);

OAI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1149),
.A2(n_1151),
.B1(n_1058),
.B2(n_1084),
.Y(n_1191)
);

OR2x2_ASAP7_75t_SL g1192 ( 
.A(n_1082),
.B(n_1147),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1128),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_1071),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1160),
.B(n_1062),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1138),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1043),
.B(n_1090),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1076),
.A2(n_1146),
.B(n_1141),
.C(n_1152),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1075),
.A2(n_1026),
.B(n_1036),
.Y(n_1199)
);

OR2x6_ASAP7_75t_L g1200 ( 
.A(n_1065),
.B(n_1164),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1144),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1145),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1026),
.A2(n_1134),
.B(n_1068),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1139),
.A2(n_1052),
.B(n_1047),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1090),
.B(n_1057),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1160),
.B(n_1092),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1057),
.A2(n_1050),
.B1(n_1048),
.B2(n_1051),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1041),
.B(n_1030),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1053),
.B(n_1125),
.Y(n_1209)
);

AO21x1_ASAP7_75t_L g1210 ( 
.A1(n_1046),
.A2(n_1079),
.B(n_1157),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1029),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1039),
.A2(n_1023),
.B(n_1073),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1080),
.B(n_1056),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1158),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1060),
.A2(n_1102),
.B1(n_1091),
.B2(n_1117),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1099),
.A2(n_1088),
.B(n_1074),
.C(n_1108),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1064),
.B(n_1083),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1064),
.B(n_1157),
.Y(n_1218)
);

INVxp67_ASAP7_75t_SL g1219 ( 
.A(n_1066),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1064),
.B(n_1148),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1064),
.B(n_1071),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1055),
.A2(n_1074),
.B(n_1020),
.Y(n_1222)
);

INVx5_ASAP7_75t_L g1223 ( 
.A(n_1071),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1094),
.B(n_1105),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1136),
.A2(n_1162),
.B1(n_1081),
.B2(n_1098),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1136),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1041),
.A2(n_1063),
.B1(n_1108),
.B2(n_1103),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1020),
.A2(n_1040),
.B(n_1054),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1104),
.Y(n_1229)
);

NOR2x1_ASAP7_75t_L g1230 ( 
.A(n_1038),
.B(n_1044),
.Y(n_1230)
);

OR2x6_ASAP7_75t_L g1231 ( 
.A(n_1041),
.B(n_1142),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1106),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1093),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1037),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1093),
.Y(n_1235)
);

CKINVDCx11_ASAP7_75t_R g1236 ( 
.A(n_1087),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1087),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1038),
.B(n_1044),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1035),
.B(n_1063),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1087),
.Y(n_1240)
);

INVx5_ASAP7_75t_L g1241 ( 
.A(n_1071),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1064),
.B(n_1071),
.Y(n_1242)
);

NOR2xp67_ASAP7_75t_L g1243 ( 
.A(n_1107),
.B(n_1079),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1107),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1107),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1107),
.B(n_1031),
.Y(n_1246)
);

OAI33xp33_ASAP7_75t_L g1247 ( 
.A1(n_1021),
.A2(n_1061),
.A3(n_1109),
.B1(n_1154),
.B2(n_1132),
.B3(n_1111),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1031),
.B(n_1142),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1127),
.A2(n_1155),
.B(n_1153),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1119),
.B(n_1135),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1100),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1109),
.B(n_1085),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1027),
.B(n_1135),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1027),
.B(n_1078),
.Y(n_1254)
);

BUFx8_ASAP7_75t_L g1255 ( 
.A(n_1109),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1049),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1109),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1089),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1111),
.B(n_1132),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1021),
.B(n_1096),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1111),
.B(n_1132),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1140),
.A2(n_1150),
.B(n_1022),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1069),
.B(n_1067),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1132),
.A2(n_1120),
.B(n_1113),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1034),
.A2(n_1130),
.B1(n_1076),
.B2(n_1110),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1072),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1028),
.Y(n_1267)
);

BUFx8_ASAP7_75t_L g1268 ( 
.A(n_1097),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1028),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1156),
.B(n_1112),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1156),
.B(n_1024),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1028),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1156),
.B(n_1112),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1156),
.B(n_1112),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1028),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1129),
.B(n_1147),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1028),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1077),
.B(n_898),
.Y(n_1278)
);

BUFx4_ASAP7_75t_SL g1279 ( 
.A(n_1136),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1130),
.A2(n_1076),
.B1(n_1110),
.B2(n_1024),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1066),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1077),
.B(n_898),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1130),
.A2(n_1076),
.B1(n_1110),
.B2(n_1024),
.Y(n_1283)
);

NOR2x1_ASAP7_75t_SL g1284 ( 
.A(n_1057),
.B(n_853),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1072),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1024),
.B(n_1118),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1024),
.B(n_1118),
.Y(n_1287)
);

OR2x6_ASAP7_75t_SL g1288 ( 
.A(n_1042),
.B(n_467),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1025),
.A2(n_725),
.B1(n_977),
.B2(n_1156),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1029),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1028),
.Y(n_1291)
);

BUFx4f_ASAP7_75t_L g1292 ( 
.A(n_1072),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1077),
.B(n_898),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1114),
.A2(n_1124),
.B(n_1115),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1029),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1136),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1042),
.B(n_670),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1025),
.A2(n_725),
.B1(n_977),
.B2(n_1156),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1024),
.B(n_1118),
.Y(n_1299)
);

BUFx4_ASAP7_75t_SL g1300 ( 
.A(n_1136),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1025),
.A2(n_725),
.B1(n_981),
.B2(n_979),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1114),
.A2(n_1124),
.B(n_1115),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1033),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1130),
.A2(n_1076),
.B1(n_1110),
.B2(n_1024),
.Y(n_1304)
);

BUFx12f_ASAP7_75t_L g1305 ( 
.A(n_1037),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1077),
.B(n_898),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1028),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1161),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1114),
.A2(n_1124),
.B(n_1115),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1114),
.A2(n_1124),
.B(n_1115),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1028),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1301),
.A2(n_1289),
.B1(n_1298),
.B2(n_1175),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1194),
.B(n_1223),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1172),
.B(n_1271),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1188),
.B(n_1286),
.Y(n_1315)
);

BUFx2_ASAP7_75t_R g1316 ( 
.A(n_1266),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_1285),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1165),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1185),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1252),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1193),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1279),
.Y(n_1322)
);

AO21x1_ASAP7_75t_L g1323 ( 
.A1(n_1280),
.A2(n_1304),
.B(n_1283),
.Y(n_1323)
);

CKINVDCx11_ASAP7_75t_R g1324 ( 
.A(n_1179),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1180),
.B(n_1284),
.Y(n_1325)
);

NAND2x1p5_ASAP7_75t_L g1326 ( 
.A(n_1194),
.B(n_1223),
.Y(n_1326)
);

AOI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1228),
.A2(n_1176),
.B(n_1170),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1225),
.A2(n_1283),
.B1(n_1280),
.B2(n_1304),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1180),
.B(n_1182),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1196),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1260),
.A2(n_1212),
.B(n_1222),
.Y(n_1331)
);

AO21x1_ASAP7_75t_L g1332 ( 
.A1(n_1265),
.A2(n_1167),
.B(n_1183),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1178),
.Y(n_1333)
);

AO21x2_ASAP7_75t_L g1334 ( 
.A1(n_1216),
.A2(n_1262),
.B(n_1310),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1201),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1194),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1202),
.Y(n_1337)
);

AOI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1294),
.A2(n_1309),
.B(n_1302),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1220),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1214),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1300),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1267),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1265),
.A2(n_1169),
.B(n_1207),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1269),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1204),
.A2(n_1203),
.B(n_1199),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_SL g1346 ( 
.A1(n_1207),
.A2(n_1221),
.B(n_1242),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1251),
.A2(n_1224),
.B(n_1253),
.Y(n_1347)
);

BUFx2_ASAP7_75t_R g1348 ( 
.A(n_1288),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1297),
.A2(n_1255),
.B1(n_1191),
.B2(n_1166),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_1186),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1188),
.A2(n_1286),
.B1(n_1287),
.B2(n_1299),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1272),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1220),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1206),
.B(n_1205),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1194),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1234),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1259),
.B(n_1261),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1264),
.A2(n_1198),
.B(n_1197),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1223),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1275),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1276),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1277),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1263),
.A2(n_1254),
.B(n_1259),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1254),
.A2(n_1261),
.B(n_1210),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1255),
.A2(n_1273),
.B1(n_1270),
.B2(n_1274),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1287),
.A2(n_1299),
.B1(n_1215),
.B2(n_1258),
.Y(n_1366)
);

BUFx2_ASAP7_75t_R g1367 ( 
.A(n_1237),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1291),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1252),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1307),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1205),
.B(n_1187),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1268),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1311),
.Y(n_1373)
);

INVx6_ASAP7_75t_L g1374 ( 
.A(n_1268),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1305),
.Y(n_1375)
);

AO21x1_ASAP7_75t_L g1376 ( 
.A1(n_1197),
.A2(n_1227),
.B(n_1213),
.Y(n_1376)
);

AO21x1_ASAP7_75t_L g1377 ( 
.A1(n_1227),
.A2(n_1213),
.B(n_1217),
.Y(n_1377)
);

AO21x1_ASAP7_75t_L g1378 ( 
.A1(n_1217),
.A2(n_1218),
.B(n_1221),
.Y(n_1378)
);

INVx5_ASAP7_75t_L g1379 ( 
.A(n_1241),
.Y(n_1379)
);

NAND2x1p5_ASAP7_75t_L g1380 ( 
.A(n_1241),
.B(n_1242),
.Y(n_1380)
);

BUFx2_ASAP7_75t_SL g1381 ( 
.A(n_1173),
.Y(n_1381)
);

OR2x6_ASAP7_75t_L g1382 ( 
.A(n_1218),
.B(n_1257),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1249),
.A2(n_1243),
.B(n_1245),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1192),
.A2(n_1181),
.B1(n_1184),
.B2(n_1226),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1308),
.A2(n_1219),
.B1(n_1281),
.B2(n_1195),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1209),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1236),
.Y(n_1387)
);

AO21x1_ASAP7_75t_L g1388 ( 
.A1(n_1232),
.A2(n_1240),
.B(n_1235),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1200),
.A2(n_1296),
.B1(n_1231),
.B2(n_1303),
.Y(n_1389)
);

BUFx2_ASAP7_75t_SL g1390 ( 
.A(n_1190),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1281),
.A2(n_1229),
.B1(n_1171),
.B2(n_1168),
.Y(n_1391)
);

CKINVDCx16_ASAP7_75t_R g1392 ( 
.A(n_1171),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1278),
.A2(n_1293),
.B1(n_1282),
.B2(n_1200),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1177),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1292),
.Y(n_1395)
);

AO21x1_ASAP7_75t_SL g1396 ( 
.A1(n_1250),
.A2(n_1233),
.B(n_1247),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1177),
.Y(n_1397)
);

AOI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1231),
.A2(n_1244),
.B(n_1246),
.Y(n_1398)
);

AND2x4_ASAP7_75t_SL g1399 ( 
.A(n_1278),
.B(n_1282),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1174),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1231),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1168),
.A2(n_1208),
.B1(n_1293),
.B2(n_1256),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1256),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1174),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1168),
.A2(n_1200),
.B1(n_1208),
.B2(n_1239),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1174),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1238),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1292),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1189),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1306),
.A2(n_1211),
.B1(n_1290),
.B2(n_1295),
.Y(n_1410)
);

BUFx2_ASAP7_75t_SL g1411 ( 
.A(n_1248),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1211),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1230),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1289),
.A2(n_1298),
.B1(n_1301),
.B2(n_1025),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_SL g1415 ( 
.A1(n_1284),
.A2(n_1183),
.B(n_1180),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1252),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1172),
.B(n_1271),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1194),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1178),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1301),
.A2(n_1025),
.B1(n_981),
.B2(n_979),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1165),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1252),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1186),
.Y(n_1423)
);

BUFx4f_ASAP7_75t_SL g1424 ( 
.A(n_1179),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1289),
.A2(n_1298),
.B1(n_1301),
.B2(n_1025),
.Y(n_1425)
);

AO21x1_ASAP7_75t_L g1426 ( 
.A1(n_1280),
.A2(n_1304),
.B(n_1283),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1165),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1180),
.B(n_1284),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1179),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1194),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1165),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1180),
.B(n_1284),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1284),
.A2(n_527),
.B1(n_486),
.B2(n_369),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1165),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1165),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1289),
.A2(n_1298),
.B1(n_1301),
.B2(n_1025),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1252),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1357),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1320),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1320),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1339),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1354),
.B(n_1371),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1339),
.Y(n_1443)
);

BUFx3_ASAP7_75t_L g1444 ( 
.A(n_1369),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1354),
.B(n_1371),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1353),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1378),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1378),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1325),
.B(n_1428),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1336),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1333),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1437),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1437),
.B(n_1369),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1416),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1416),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1386),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1422),
.B(n_1325),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1422),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1388),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1327),
.A2(n_1338),
.B(n_1345),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1428),
.B(n_1432),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1388),
.Y(n_1462)
);

CKINVDCx11_ASAP7_75t_R g1463 ( 
.A(n_1350),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1411),
.B(n_1382),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1361),
.Y(n_1465)
);

INVx5_ASAP7_75t_L g1466 ( 
.A(n_1379),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1334),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1347),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1419),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1364),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1432),
.B(n_1382),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1364),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1324),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1364),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1336),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1346),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1382),
.B(n_1379),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1382),
.B(n_1379),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1384),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1412),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1329),
.B(n_1363),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1343),
.A2(n_1328),
.B(n_1358),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1363),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1346),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1329),
.B(n_1363),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1412),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1336),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_R g1488 ( 
.A(n_1324),
.B(n_1429),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1318),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1319),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1321),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1331),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1330),
.Y(n_1493)
);

AO21x2_ASAP7_75t_L g1494 ( 
.A1(n_1376),
.A2(n_1383),
.B(n_1377),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1314),
.B(n_1351),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1376),
.B(n_1315),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1322),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1335),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1337),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1334),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1340),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1429),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1342),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1433),
.A2(n_1420),
.B1(n_1366),
.B2(n_1436),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1338),
.A2(n_1377),
.B(n_1323),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1344),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1352),
.B(n_1360),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1362),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1331),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1368),
.B(n_1370),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1323),
.B(n_1426),
.Y(n_1511)
);

BUFx4f_ASAP7_75t_L g1512 ( 
.A(n_1326),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1426),
.B(n_1373),
.Y(n_1513)
);

AO21x2_ASAP7_75t_L g1514 ( 
.A1(n_1383),
.A2(n_1332),
.B(n_1331),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1435),
.Y(n_1515)
);

INVxp33_ASAP7_75t_SL g1516 ( 
.A(n_1341),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1421),
.B(n_1427),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1431),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1332),
.A2(n_1415),
.B(n_1403),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1434),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1414),
.A2(n_1425),
.B(n_1312),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1334),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1407),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1417),
.B(n_1385),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1404),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1415),
.A2(n_1398),
.B(n_1409),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1396),
.B(n_1406),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1372),
.Y(n_1528)
);

INVxp67_ASAP7_75t_SL g1529 ( 
.A(n_1470),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1471),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1481),
.B(n_1396),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1470),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1489),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1496),
.B(n_1349),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1489),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1482),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1481),
.B(n_1406),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1485),
.B(n_1400),
.Y(n_1538)
);

NOR2x1_ASAP7_75t_L g1539 ( 
.A(n_1482),
.B(n_1413),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1439),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1439),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1440),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1490),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1521),
.A2(n_1393),
.B1(n_1365),
.B2(n_1374),
.C(n_1372),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1485),
.B(n_1389),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1449),
.B(n_1404),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1451),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1444),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1465),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1440),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1471),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1461),
.B(n_1442),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1490),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1454),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1444),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1472),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1454),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1469),
.Y(n_1558)
);

NAND2x1_ASAP7_75t_L g1559 ( 
.A(n_1476),
.B(n_1313),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1496),
.B(n_1380),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1445),
.B(n_1505),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1513),
.B(n_1430),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1504),
.A2(n_1372),
.B1(n_1374),
.B2(n_1375),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1511),
.A2(n_1348),
.B1(n_1374),
.B2(n_1372),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1495),
.B(n_1374),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1455),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1505),
.B(n_1430),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1505),
.B(n_1492),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1505),
.B(n_1430),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1472),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1493),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1457),
.B(n_1514),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1455),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1482),
.A2(n_1375),
.B1(n_1387),
.B2(n_1397),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1474),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1493),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1444),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1513),
.B(n_1359),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1511),
.B(n_1359),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1498),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1491),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1498),
.Y(n_1582)
);

OAI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1447),
.A2(n_1448),
.B(n_1459),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1514),
.B(n_1418),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1514),
.B(n_1418),
.Y(n_1585)
);

BUFx12f_ASAP7_75t_L g1586 ( 
.A(n_1463),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1501),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1483),
.B(n_1359),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1525),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1501),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1483),
.B(n_1355),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1581),
.B(n_1547),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1438),
.Y(n_1593)
);

NAND3xp33_ASAP7_75t_L g1594 ( 
.A(n_1536),
.B(n_1448),
.C(n_1447),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1564),
.B(n_1528),
.Y(n_1595)
);

OA21x2_ASAP7_75t_L g1596 ( 
.A1(n_1583),
.A2(n_1460),
.B(n_1462),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1586),
.B(n_1516),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1564),
.B(n_1528),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1565),
.B(n_1512),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1574),
.A2(n_1479),
.B1(n_1456),
.B2(n_1497),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1581),
.B(n_1523),
.Y(n_1601)
);

OAI221xp5_ASAP7_75t_SL g1602 ( 
.A1(n_1574),
.A2(n_1462),
.B1(n_1524),
.B2(n_1453),
.C(n_1523),
.Y(n_1602)
);

OAI221xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1563),
.A2(n_1524),
.B1(n_1453),
.B2(n_1484),
.C(n_1476),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1547),
.B(n_1499),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1563),
.A2(n_1484),
.B1(n_1458),
.B2(n_1452),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1552),
.B(n_1458),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1552),
.B(n_1458),
.Y(n_1607)
);

OAI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1536),
.A2(n_1464),
.B1(n_1392),
.B2(n_1466),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1549),
.B(n_1558),
.Y(n_1609)
);

AND2x2_ASAP7_75t_SL g1610 ( 
.A(n_1536),
.B(n_1477),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1549),
.B(n_1507),
.Y(n_1611)
);

OAI21xp33_ASAP7_75t_SL g1612 ( 
.A1(n_1552),
.A2(n_1452),
.B(n_1486),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1558),
.B(n_1561),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1561),
.B(n_1531),
.Y(n_1614)
);

NOR3xp33_ASAP7_75t_L g1615 ( 
.A(n_1536),
.B(n_1467),
.C(n_1522),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1534),
.A2(n_1515),
.B1(n_1508),
.B2(n_1506),
.C(n_1503),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1534),
.A2(n_1526),
.B1(n_1527),
.B2(n_1391),
.Y(n_1617)
);

NOR3xp33_ASAP7_75t_L g1618 ( 
.A(n_1536),
.B(n_1522),
.C(n_1467),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_SL g1619 ( 
.A(n_1544),
.B(n_1488),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1545),
.A2(n_1526),
.B1(n_1527),
.B2(n_1397),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1545),
.A2(n_1526),
.B1(n_1394),
.B2(n_1401),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1545),
.A2(n_1394),
.B1(n_1401),
.B2(n_1443),
.Y(n_1622)
);

NOR3xp33_ASAP7_75t_L g1623 ( 
.A(n_1539),
.B(n_1467),
.C(n_1522),
.Y(n_1623)
);

AOI211xp5_ASAP7_75t_L g1624 ( 
.A1(n_1544),
.A2(n_1488),
.B(n_1502),
.C(n_1473),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1531),
.B(n_1480),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1531),
.B(n_1480),
.Y(n_1626)
);

OAI221xp5_ASAP7_75t_L g1627 ( 
.A1(n_1583),
.A2(n_1539),
.B1(n_1565),
.B2(n_1568),
.C(n_1560),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1538),
.B(n_1486),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1538),
.B(n_1541),
.Y(n_1629)
);

OAI21xp5_ASAP7_75t_SL g1630 ( 
.A1(n_1568),
.A2(n_1399),
.B(n_1387),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1538),
.B(n_1507),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1541),
.B(n_1510),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1560),
.B(n_1512),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1579),
.B(n_1512),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1568),
.A2(n_1494),
.B1(n_1477),
.B2(n_1478),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1579),
.B(n_1510),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1540),
.B(n_1517),
.Y(n_1637)
);

NAND3xp33_ASAP7_75t_L g1638 ( 
.A(n_1562),
.B(n_1519),
.C(n_1508),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1537),
.A2(n_1441),
.B1(n_1443),
.B2(n_1446),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1540),
.B(n_1517),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1540),
.B(n_1503),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1542),
.B(n_1506),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1542),
.B(n_1515),
.Y(n_1643)
);

OAI221xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1562),
.A2(n_1518),
.B1(n_1520),
.B2(n_1464),
.C(n_1405),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1542),
.B(n_1518),
.Y(n_1645)
);

OAI221xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1578),
.A2(n_1520),
.B1(n_1464),
.B2(n_1509),
.C(n_1468),
.Y(n_1646)
);

NAND3xp33_ASAP7_75t_L g1647 ( 
.A(n_1578),
.B(n_1519),
.C(n_1509),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1550),
.B(n_1519),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1550),
.B(n_1519),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1550),
.B(n_1525),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1554),
.B(n_1494),
.Y(n_1651)
);

NAND2xp33_ASAP7_75t_SL g1652 ( 
.A(n_1559),
.B(n_1350),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1638),
.B(n_1529),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1638),
.B(n_1593),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1614),
.B(n_1606),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1530),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1592),
.B(n_1554),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1593),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1613),
.B(n_1554),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1606),
.B(n_1557),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1611),
.B(n_1557),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1607),
.B(n_1557),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1641),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1607),
.B(n_1566),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1609),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1601),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1612),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1637),
.B(n_1566),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1648),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1640),
.B(n_1566),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1642),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1597),
.B(n_1586),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1612),
.Y(n_1673)
);

INVxp67_ASAP7_75t_SL g1674 ( 
.A(n_1649),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1651),
.B(n_1529),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1604),
.Y(n_1676)
);

INVx2_ASAP7_75t_SL g1677 ( 
.A(n_1650),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1625),
.B(n_1566),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1636),
.B(n_1573),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1643),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1596),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1625),
.B(n_1573),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1631),
.B(n_1573),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1626),
.B(n_1573),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1626),
.B(n_1572),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1645),
.B(n_1532),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1628),
.B(n_1572),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1596),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1628),
.B(n_1572),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1616),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1632),
.B(n_1537),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1629),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1619),
.B(n_1586),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1627),
.B(n_1537),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1596),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1619),
.A2(n_1494),
.B1(n_1551),
.B2(n_1530),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1647),
.Y(n_1697)
);

NAND3xp33_ASAP7_75t_L g1698 ( 
.A(n_1624),
.B(n_1587),
.C(n_1582),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1610),
.B(n_1530),
.Y(n_1699)
);

NOR2x1_ASAP7_75t_L g1700 ( 
.A(n_1630),
.B(n_1559),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1596),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1647),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1594),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1658),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1658),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1602),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1690),
.B(n_1582),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1667),
.B(n_1610),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1673),
.B(n_1655),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1686),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1686),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1690),
.B(n_1703),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1703),
.B(n_1582),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1663),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1663),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1693),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1681),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1697),
.B(n_1587),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1697),
.B(n_1587),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1702),
.B(n_1533),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1673),
.B(n_1610),
.Y(n_1721)
);

INVxp67_ASAP7_75t_SL g1722 ( 
.A(n_1653),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1665),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1681),
.Y(n_1724)
);

NAND4xp75_ASAP7_75t_L g1725 ( 
.A(n_1702),
.B(n_1598),
.C(n_1595),
.D(n_1624),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1655),
.B(n_1635),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1654),
.B(n_1589),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1656),
.B(n_1630),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1656),
.B(n_1546),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1702),
.B(n_1533),
.Y(n_1730)
);

NAND4xp25_ASAP7_75t_L g1731 ( 
.A(n_1698),
.B(n_1603),
.C(n_1594),
.D(n_1600),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1676),
.B(n_1535),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1671),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1654),
.B(n_1589),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1671),
.B(n_1535),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1666),
.B(n_1543),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1700),
.Y(n_1737)
);

NAND2x1p5_ASAP7_75t_L g1738 ( 
.A(n_1700),
.B(n_1466),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1680),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1681),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1680),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1672),
.B(n_1586),
.Y(n_1742)
);

NOR2x1p5_ASAP7_75t_L g1743 ( 
.A(n_1698),
.B(n_1559),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1708),
.B(n_1656),
.Y(n_1744)
);

NOR2x1_ASAP7_75t_L g1745 ( 
.A(n_1725),
.B(n_1423),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1724),
.Y(n_1746)
);

NAND2x1_ASAP7_75t_SL g1747 ( 
.A(n_1708),
.B(n_1721),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1725),
.A2(n_1653),
.B(n_1696),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1712),
.B(n_1661),
.Y(n_1749)
);

BUFx2_ASAP7_75t_SL g1750 ( 
.A(n_1737),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1732),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1723),
.B(n_1669),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1707),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1743),
.B(n_1699),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1736),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1737),
.A2(n_1706),
.B(n_1731),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1731),
.B(n_1661),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1706),
.B(n_1692),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1735),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1722),
.B(n_1710),
.Y(n_1760)
);

BUFx2_ASAP7_75t_SL g1761 ( 
.A(n_1743),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1710),
.B(n_1674),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1735),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1718),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1704),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1727),
.B(n_1692),
.Y(n_1766)
);

AOI22x1_ASAP7_75t_L g1767 ( 
.A1(n_1738),
.A2(n_1701),
.B1(n_1341),
.B2(n_1356),
.Y(n_1767)
);

NOR3x1_ASAP7_75t_L g1768 ( 
.A(n_1727),
.B(n_1694),
.C(n_1677),
.Y(n_1768)
);

NOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1742),
.B(n_1423),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1711),
.B(n_1694),
.Y(n_1770)
);

OAI32xp33_ASAP7_75t_L g1771 ( 
.A1(n_1721),
.A2(n_1695),
.A3(n_1688),
.B1(n_1675),
.B2(n_1659),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1738),
.A2(n_1699),
.B(n_1605),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1711),
.B(n_1677),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1734),
.B(n_1691),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1719),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1709),
.B(n_1687),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1734),
.B(n_1691),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1704),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1709),
.B(n_1656),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1716),
.B(n_1356),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1713),
.B(n_1657),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1728),
.B(n_1685),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1728),
.B(n_1424),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1724),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1705),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1705),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1738),
.A2(n_1683),
.B1(n_1679),
.B2(n_1685),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1779),
.B(n_1726),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1765),
.Y(n_1789)
);

NOR2x1_ASAP7_75t_L g1790 ( 
.A(n_1745),
.B(n_1726),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1756),
.B(n_1753),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1757),
.B(n_1714),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1778),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1746),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1785),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1747),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1749),
.B(n_1714),
.Y(n_1797)
);

NAND3xp33_ASAP7_75t_SL g1798 ( 
.A(n_1748),
.B(n_1695),
.C(n_1688),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1770),
.B(n_1760),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1786),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1769),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1779),
.B(n_1729),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1759),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1751),
.B(n_1715),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1763),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1744),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1780),
.Y(n_1807)
);

INVxp67_ASAP7_75t_L g1808 ( 
.A(n_1780),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1755),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1754),
.B(n_1715),
.Y(n_1810)
);

OR2x6_ASAP7_75t_L g1811 ( 
.A(n_1761),
.B(n_1750),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1783),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1766),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1774),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1758),
.B(n_1720),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1783),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1764),
.B(n_1316),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1777),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1782),
.B(n_1729),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1752),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1746),
.A2(n_1695),
.B1(n_1688),
.B2(n_1724),
.Y(n_1821)
);

CKINVDCx16_ASAP7_75t_R g1822 ( 
.A(n_1754),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1784),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1799),
.B(n_1781),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1789),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_SL g1826 ( 
.A1(n_1811),
.A2(n_1754),
.B(n_1408),
.Y(n_1826)
);

AOI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1790),
.A2(n_1771),
.B(n_1764),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1820),
.B(n_1775),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1798),
.A2(n_1784),
.B1(n_1772),
.B2(n_1617),
.Y(n_1829)
);

OAI322xp33_ASAP7_75t_L g1830 ( 
.A1(n_1791),
.A2(n_1762),
.A3(n_1775),
.B1(n_1773),
.B2(n_1730),
.C1(n_1776),
.C2(n_1768),
.Y(n_1830)
);

NOR2xp67_ASAP7_75t_L g1831 ( 
.A(n_1806),
.B(n_1744),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1806),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1812),
.B(n_1317),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1793),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1820),
.B(n_1782),
.Y(n_1835)
);

NAND2x1_ASAP7_75t_L g1836 ( 
.A(n_1811),
.B(n_1810),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1822),
.A2(n_1767),
.B1(n_1787),
.B2(n_1741),
.Y(n_1837)
);

AOI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1792),
.A2(n_1796),
.B1(n_1821),
.B2(n_1799),
.C(n_1809),
.Y(n_1838)
);

OAI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1821),
.A2(n_1740),
.B1(n_1717),
.B2(n_1675),
.C(n_1620),
.Y(n_1839)
);

NOR4xp25_ASAP7_75t_L g1840 ( 
.A(n_1807),
.B(n_1741),
.C(n_1739),
.D(n_1733),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1795),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1813),
.B(n_1733),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1814),
.B(n_1739),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1818),
.B(n_1687),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1788),
.B(n_1689),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1808),
.B(n_1689),
.Y(n_1846)
);

A2O1A1Ixp33_ASAP7_75t_L g1847 ( 
.A1(n_1817),
.A2(n_1644),
.B(n_1740),
.C(n_1717),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1800),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1817),
.A2(n_1801),
.B1(n_1788),
.B2(n_1823),
.Y(n_1849)
);

OAI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1815),
.A2(n_1646),
.B1(n_1621),
.B2(n_1622),
.C(n_1652),
.Y(n_1850)
);

INVx2_ASAP7_75t_SL g1851 ( 
.A(n_1836),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1833),
.B(n_1816),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1824),
.Y(n_1853)
);

AND2x2_ASAP7_75t_SL g1854 ( 
.A(n_1840),
.B(n_1838),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1827),
.A2(n_1823),
.B1(n_1794),
.B2(n_1803),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1835),
.B(n_1805),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1832),
.B(n_1819),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1843),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1832),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1831),
.B(n_1811),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1842),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1828),
.B(n_1819),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1833),
.B(n_1811),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1845),
.B(n_1815),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1825),
.B(n_1797),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1834),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_R g1867 ( 
.A1(n_1830),
.A2(n_1794),
.B1(n_1408),
.B2(n_1395),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1829),
.A2(n_1804),
.B1(n_1810),
.B2(n_1802),
.Y(n_1868)
);

CKINVDCx16_ASAP7_75t_R g1869 ( 
.A(n_1849),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1841),
.B(n_1810),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_SL g1871 ( 
.A1(n_1855),
.A2(n_1837),
.B(n_1847),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1851),
.B(n_1826),
.Y(n_1872)
);

AOI21xp33_ASAP7_75t_L g1873 ( 
.A1(n_1854),
.A2(n_1848),
.B(n_1847),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1854),
.A2(n_1839),
.B1(n_1850),
.B2(n_1846),
.Y(n_1874)
);

AOI32xp33_ASAP7_75t_L g1875 ( 
.A1(n_1855),
.A2(n_1844),
.A3(n_1802),
.B1(n_1652),
.B2(n_1395),
.Y(n_1875)
);

AOI222xp33_ASAP7_75t_L g1876 ( 
.A1(n_1868),
.A2(n_1639),
.B1(n_1584),
.B2(n_1585),
.C1(n_1567),
.C2(n_1569),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1868),
.A2(n_1615),
.B1(n_1618),
.B2(n_1569),
.C(n_1567),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1869),
.A2(n_1659),
.B1(n_1679),
.B2(n_1670),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_R g1879 ( 
.A(n_1852),
.B(n_1317),
.Y(n_1879)
);

OAI211xp5_ASAP7_75t_L g1880 ( 
.A1(n_1863),
.A2(n_1317),
.B(n_1662),
.C(n_1660),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1857),
.A2(n_1599),
.B(n_1668),
.Y(n_1881)
);

OAI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1867),
.A2(n_1381),
.B1(n_1390),
.B2(n_1623),
.C(n_1402),
.Y(n_1882)
);

NAND2x1p5_ASAP7_75t_L g1883 ( 
.A(n_1872),
.B(n_1860),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1879),
.B(n_1863),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_SL g1885 ( 
.A1(n_1871),
.A2(n_1852),
.B(n_1853),
.Y(n_1885)
);

NAND3xp33_ASAP7_75t_L g1886 ( 
.A(n_1873),
.B(n_1859),
.C(n_1866),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1874),
.A2(n_1870),
.B(n_1862),
.Y(n_1887)
);

NAND3xp33_ASAP7_75t_L g1888 ( 
.A(n_1875),
.B(n_1859),
.C(n_1858),
.Y(n_1888)
);

NAND5xp2_ASAP7_75t_L g1889 ( 
.A(n_1880),
.B(n_1861),
.C(n_1856),
.D(n_1864),
.E(n_1865),
.Y(n_1889)
);

OAI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1882),
.A2(n_1878),
.B1(n_1877),
.B2(n_1881),
.Y(n_1890)
);

NAND4xp75_ASAP7_75t_SL g1891 ( 
.A(n_1876),
.B(n_1660),
.C(n_1662),
.D(n_1682),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_L g1892 ( 
.A(n_1873),
.B(n_1500),
.C(n_1467),
.Y(n_1892)
);

AOI211x1_ASAP7_75t_L g1893 ( 
.A1(n_1886),
.A2(n_1684),
.B(n_1682),
.C(n_1678),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1885),
.B(n_1683),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1887),
.A2(n_1670),
.B(n_1668),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1889),
.B(n_1367),
.Y(n_1896)
);

NAND3xp33_ASAP7_75t_SL g1897 ( 
.A(n_1883),
.B(n_1884),
.C(n_1888),
.Y(n_1897)
);

NOR2x1_ASAP7_75t_L g1898 ( 
.A(n_1891),
.B(n_1678),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1896),
.B(n_1664),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1893),
.B(n_1890),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1894),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1897),
.A2(n_1892),
.B1(n_1608),
.B2(n_1664),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1895),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1898),
.A2(n_1684),
.B1(n_1588),
.B2(n_1591),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1894),
.Y(n_1905)
);

AO22x1_ASAP7_75t_L g1906 ( 
.A1(n_1901),
.A2(n_1466),
.B1(n_1548),
.B2(n_1555),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1905),
.Y(n_1907)
);

NOR2x1_ASAP7_75t_L g1908 ( 
.A(n_1903),
.B(n_1577),
.Y(n_1908)
);

NAND4xp75_ASAP7_75t_L g1909 ( 
.A(n_1900),
.B(n_1634),
.C(n_1633),
.D(n_1584),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1899),
.B(n_1548),
.Y(n_1910)
);

NOR2xp67_ASAP7_75t_L g1911 ( 
.A(n_1902),
.B(n_1904),
.Y(n_1911)
);

AND2x2_ASAP7_75t_SL g1912 ( 
.A(n_1907),
.B(n_1399),
.Y(n_1912)
);

OR2x6_ASAP7_75t_L g1913 ( 
.A(n_1908),
.B(n_1326),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1911),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1914),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_SL g1916 ( 
.A(n_1915),
.B(n_1912),
.C(n_1913),
.Y(n_1916)
);

OAI22x1_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1910),
.B1(n_1913),
.B2(n_1909),
.Y(n_1917)
);

OAI221xp5_ASAP7_75t_L g1918 ( 
.A1(n_1916),
.A2(n_1906),
.B1(n_1590),
.B2(n_1580),
.C(n_1576),
.Y(n_1918)
);

AOI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1917),
.A2(n_1576),
.B(n_1543),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1918),
.A2(n_1571),
.B(n_1553),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1919),
.A2(n_1556),
.B(n_1570),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1920),
.A2(n_1532),
.B1(n_1556),
.B2(n_1570),
.C(n_1575),
.Y(n_1922)
);

NAND3xp33_ASAP7_75t_L g1923 ( 
.A(n_1922),
.B(n_1468),
.C(n_1466),
.Y(n_1923)
);

AOI222xp33_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1921),
.B1(n_1585),
.B2(n_1584),
.C1(n_1532),
.C2(n_1570),
.Y(n_1924)
);

OAI221xp5_ASAP7_75t_R g1925 ( 
.A1(n_1924),
.A2(n_1410),
.B1(n_1555),
.B2(n_1548),
.C(n_1577),
.Y(n_1925)
);

AOI211xp5_ASAP7_75t_L g1926 ( 
.A1(n_1925),
.A2(n_1475),
.B(n_1450),
.C(n_1487),
.Y(n_1926)
);


endmodule