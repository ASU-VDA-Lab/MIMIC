module real_jpeg_6563_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_2),
.A2(n_107),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_2),
.A2(n_107),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_2),
.A2(n_35),
.B1(n_107),
.B2(n_297),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_3),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_3),
.A2(n_42),
.B1(n_71),
.B2(n_73),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_42),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_3),
.A2(n_42),
.B1(n_92),
.B2(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_4),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_4),
.A2(n_63),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_4),
.A2(n_63),
.B1(n_221),
.B2(n_382),
.Y(n_381)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_5),
.Y(n_128)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_6),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_6),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_6),
.Y(n_312)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_7),
.Y(n_212)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_8),
.Y(n_99)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_9),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_10),
.A2(n_28),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_10),
.A2(n_28),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_10),
.B(n_93),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_10),
.A2(n_127),
.B(n_257),
.C(n_264),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_10),
.B(n_287),
.C(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_10),
.B(n_125),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_10),
.B(n_175),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_10),
.B(n_48),
.Y(n_324)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_11),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_363),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_224),
.B(n_361),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_190),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_15),
.B(n_190),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_15),
.B(n_365),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_15),
.B(n_365),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_155),
.CI(n_164),
.CON(n_15),
.SN(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_83),
.B2(n_84),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_17),
.B(n_85),
.C(n_116),
.Y(n_386)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_19),
.B(n_46),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_20),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_22),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_24),
.A2(n_34),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_24),
.B(n_34),
.Y(n_235)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_27),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_28),
.A2(n_88),
.B(n_90),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_28),
.B(n_91),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_28),
.A2(n_258),
.B(n_261),
.Y(n_257)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_30),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_31),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_32),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_33),
.A2(n_167),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_34),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_34),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_38),
.B(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_40),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_40),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_58),
.B(n_69),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_47),
.A2(n_161),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_47),
.B(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_48),
.B(n_70),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_48),
.B(n_272),
.Y(n_291)
);

AO22x2_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_58),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_61),
.Y(n_263)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_62),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_62),
.Y(n_285)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_69),
.B(n_291),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_69),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_75),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_75),
.B(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_116),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_104),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_93),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_87),
.B(n_110),
.Y(n_240)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_87),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_108),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_90),
.Y(n_206)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_93),
.B(n_105),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_93),
.B(n_186),
.Y(n_196)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_93),
.Y(n_376)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_100),
.B2(n_102),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_101),
.Y(n_209)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_104),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.Y(n_104)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_110),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_110),
.Y(n_375)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_136),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_117),
.B(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_118),
.Y(n_245)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_120),
.Y(n_266)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_125),
.A2(n_137),
.B(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_125),
.B(n_218),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_125),
.A2(n_244),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_126),
.B(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_129),
.Y(n_273)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_136),
.B(n_246),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_149),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_137),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_138),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_142),
.B1(n_144),
.B2(n_146),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_141),
.Y(n_260)
);

AOI32xp33_ASAP7_75t_L g201 ( 
.A1(n_142),
.A2(n_202),
.A3(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_201)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_147),
.Y(n_382)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_149),
.Y(n_216)
);

INVx6_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_163),
.Y(n_155)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_156),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_156),
.A2(n_163),
.B1(n_256),
.B2(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_156),
.B(n_160),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_156),
.A2(n_163),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_162),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_162),
.B(n_271),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_182),
.C(n_184),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_176),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_166),
.B(n_176),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_172),
.B(n_173),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_173),
.B(n_295),
.Y(n_323)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_177),
.B(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_189),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.C(n_223),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_191),
.B(n_223),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_194),
.B(n_356),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.C(n_213),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_195),
.B(n_213),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_197),
.B(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_201),
.Y(n_237)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_345),
.B(n_358),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_277),
.B(n_344),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_251),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_227),
.B(n_251),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_238),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_236),
.B2(n_237),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_230),
.B(n_236),
.C(n_238),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.C(n_234),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_235),
.B(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_239),
.B(n_242),
.C(n_248),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_267),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_252),
.B(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_255),
.A2(n_267),
.B1(n_268),
.B2(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_255),
.Y(n_341)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_256),
.Y(n_336)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_270),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_338),
.B(n_343),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_328),
.B(n_337),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_304),
.B(n_327),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_292),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_292),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_290),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_282),
.A2(n_283),
.B1(n_290),
.B2(n_307),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_299),
.Y(n_292)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_300),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_302),
.C(n_330),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_313),
.B(n_326),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_308),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_322),
.B(n_325),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_321),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_331),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_334),
.C(n_335),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_342),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_354),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_348),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_351),
.C(n_352),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_354),
.A2(n_359),
.B(n_360),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_357),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_357),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_387),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_386),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_378),
.B2(n_379),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_371),
.B2(n_372),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B(n_377),
.Y(n_374)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_383),
.B(n_385),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_380),
.B(n_383),
.Y(n_385)
);


endmodule