module real_aes_7619_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_792;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_766;
wire n_329;
wire n_852;
wire n_857;
wire n_461;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_860;
wire n_748;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_898;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_385;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_0), .A2(n_249), .B1(n_690), .B2(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_1), .A2(n_115), .B1(n_477), .B2(n_578), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_2), .A2(n_95), .B1(n_386), .B2(n_472), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_3), .B(n_438), .Y(n_705) );
AOI22xp5_ASAP7_75t_SL g774 ( .A1(n_4), .A2(n_64), .B1(n_382), .B2(n_469), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_5), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_6), .A2(n_25), .B1(n_600), .B2(n_826), .Y(n_825) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_7), .A2(n_158), .B1(n_432), .B2(n_436), .C(n_439), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_8), .A2(n_217), .B1(n_465), .B2(n_469), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_9), .A2(n_105), .B1(n_335), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_10), .A2(n_177), .B1(n_390), .B2(n_392), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_11), .A2(n_176), .B1(n_472), .B2(n_651), .Y(n_786) );
AOI211xp5_ASAP7_75t_L g573 ( .A1(n_12), .A2(n_574), .B(n_575), .C(n_579), .Y(n_573) );
XOR2x2_ASAP7_75t_L g528 ( .A(n_13), .B(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_14), .Y(n_666) );
OA22x2_ASAP7_75t_L g456 ( .A1(n_15), .A2(n_457), .B1(n_458), .B2(n_498), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_15), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_16), .A2(n_193), .B1(n_421), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g564 ( .A1(n_17), .A2(n_269), .B1(n_491), .B2(n_494), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g712 ( .A1(n_18), .A2(n_128), .B1(n_390), .B2(n_628), .Y(n_712) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_19), .A2(n_246), .B1(n_392), .B2(n_462), .Y(n_461) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_20), .A2(n_134), .B1(n_170), .B2(n_446), .C1(n_449), .C2(n_450), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_21), .A2(n_149), .B1(n_504), .B2(n_586), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_22), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_23), .A2(n_229), .B1(n_467), .B2(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_24), .A2(n_201), .B1(n_518), .B2(n_586), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_26), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_27), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_28), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_29), .A2(n_40), .B1(n_377), .B2(n_684), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_30), .A2(n_274), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_31), .A2(n_80), .B1(n_426), .B2(n_532), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_32), .Y(n_620) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_33), .A2(n_87), .B1(n_310), .B2(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g847 ( .A(n_33), .Y(n_847) );
AOI22xp5_ASAP7_75t_SL g772 ( .A1(n_34), .A2(n_278), .B1(n_571), .B2(n_773), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_35), .A2(n_41), .B1(n_451), .B2(n_494), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_36), .Y(n_871) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_37), .A2(n_287), .B(n_295), .C(n_849), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_38), .A2(n_102), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_39), .A2(n_42), .B1(n_436), .B2(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_43), .A2(n_781), .B1(n_805), .B2(n_806), .Y(n_780) );
INVx1_ASAP7_75t_L g805 ( .A(n_43), .Y(n_805) );
AOI22xp5_ASAP7_75t_SL g768 ( .A1(n_44), .A2(n_152), .B1(n_574), .B2(n_626), .Y(n_768) );
AOI222xp33_ASAP7_75t_L g827 ( .A1(n_45), .A2(n_136), .B1(n_208), .B2(n_483), .C1(n_828), .C2(n_829), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_46), .A2(n_277), .B1(n_449), .B2(n_492), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_47), .A2(n_60), .B1(n_828), .B2(n_829), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_48), .A2(n_130), .B1(n_477), .B2(n_479), .Y(n_476) );
AO22x2_ASAP7_75t_L g313 ( .A1(n_49), .A2(n_91), .B1(n_310), .B2(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g848 ( .A(n_49), .Y(n_848) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_50), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_51), .A2(n_203), .B1(n_382), .B2(n_386), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_52), .A2(n_107), .B1(n_372), .B2(n_377), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_53), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_54), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_55), .B(n_801), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_56), .A2(n_285), .B1(n_387), .B2(n_540), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_57), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_58), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_59), .Y(n_863) );
INVx1_ASAP7_75t_L g889 ( .A(n_61), .Y(n_889) );
XNOR2xp5_ASAP7_75t_L g555 ( .A(n_62), .B(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_63), .A2(n_253), .B1(n_626), .B2(n_785), .Y(n_824) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_65), .A2(n_153), .B1(n_492), .B2(n_510), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_66), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_67), .A2(n_256), .B1(n_426), .B2(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_68), .A2(n_138), .B1(n_624), .B2(n_626), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_69), .A2(n_202), .B1(n_364), .B2(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_70), .B(n_433), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_71), .A2(n_121), .B1(n_535), .B2(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g550 ( .A(n_72), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_73), .A2(n_174), .B1(n_540), .B2(n_789), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g765 ( .A1(n_74), .A2(n_262), .B1(n_546), .B2(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_75), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_76), .A2(n_165), .B1(n_475), .B2(n_504), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_77), .A2(n_268), .B1(n_336), .B2(n_552), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_78), .A2(n_397), .B1(n_452), .B2(n_453), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_78), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_79), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_81), .A2(n_155), .B1(n_785), .B2(n_908), .Y(n_907) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_82), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_83), .A2(n_221), .B1(n_495), .B2(n_546), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_84), .A2(n_135), .B1(n_403), .B2(n_540), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_85), .A2(n_168), .B1(n_684), .B2(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_86), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_88), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_89), .A2(n_141), .B1(n_382), .B2(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_90), .A2(n_147), .B1(n_414), .B2(n_534), .Y(n_905) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_92), .A2(n_192), .B1(n_362), .B2(n_367), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_93), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_94), .A2(n_223), .B1(n_518), .B2(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g764 ( .A(n_96), .B(n_432), .Y(n_764) );
AOI22xp33_ASAP7_75t_SL g572 ( .A1(n_97), .A2(n_267), .B1(n_402), .B2(n_462), .Y(n_572) );
INVx1_ASAP7_75t_L g293 ( .A(n_98), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_99), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_100), .A2(n_151), .B1(n_342), .B2(n_451), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_101), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_103), .A2(n_200), .B1(n_475), .B2(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g290 ( .A(n_104), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_106), .A2(n_120), .B1(n_814), .B2(n_815), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_108), .B(n_578), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_109), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_110), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_111), .A2(n_178), .B1(n_433), .B2(n_566), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_112), .Y(n_897) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_113), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_114), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g647 ( .A1(n_116), .A2(n_143), .B1(n_491), .B2(n_494), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_117), .A2(n_166), .B1(n_451), .B2(n_552), .Y(n_898) );
OA22x2_ASAP7_75t_L g607 ( .A1(n_118), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_118), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_119), .A2(n_142), .B1(n_492), .B2(n_552), .Y(n_706) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_122), .A2(n_154), .B1(n_491), .B2(n_494), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_123), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_124), .A2(n_245), .B1(n_570), .B2(n_688), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_125), .A2(n_226), .B1(n_624), .B2(n_814), .Y(n_867) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_126), .A2(n_183), .B1(n_451), .B2(n_759), .Y(n_758) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_127), .A2(n_233), .B1(n_433), .B2(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_129), .A2(n_173), .B1(n_586), .B2(n_817), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_131), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_132), .A2(n_227), .B1(n_373), .B2(n_391), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_133), .A2(n_190), .B1(n_402), .B2(n_624), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_137), .B(n_644), .Y(n_667) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_139), .A2(n_231), .B1(n_569), .B2(n_651), .Y(n_650) );
XOR2x2_ASAP7_75t_L g299 ( .A(n_140), .B(n_300), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_144), .A2(n_228), .B1(n_386), .B2(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_145), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_146), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_148), .Y(n_757) );
INVx2_ASAP7_75t_L g294 ( .A(n_150), .Y(n_294) );
INVx1_ASAP7_75t_L g714 ( .A(n_156), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_157), .B(n_549), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_159), .B(n_438), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_160), .B(n_543), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_161), .A2(n_279), .B1(n_372), .B2(n_826), .Y(n_868) );
AND2x6_ASAP7_75t_L g289 ( .A(n_162), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_162), .Y(n_841) );
AO22x2_ASAP7_75t_L g319 ( .A1(n_163), .A2(n_237), .B1(n_310), .B2(n_314), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_164), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_167), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_169), .A2(n_265), .B1(n_509), .B2(n_510), .Y(n_591) );
AOI22xp5_ASAP7_75t_SL g769 ( .A1(n_171), .A2(n_234), .B1(n_535), .B2(n_770), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_172), .A2(n_238), .B1(n_403), .B2(n_773), .Y(n_909) );
AOI22xp33_ASAP7_75t_SL g630 ( .A1(n_175), .A2(n_252), .B1(n_540), .B2(n_571), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_179), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_180), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_181), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_182), .A2(n_225), .B1(n_343), .B2(n_492), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_184), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_185), .B(n_704), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_186), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_187), .A2(n_284), .B1(n_543), .B2(n_544), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g631 ( .A1(n_188), .A2(n_197), .B1(n_538), .B2(n_569), .Y(n_631) );
AO22x2_ASAP7_75t_L g317 ( .A1(n_189), .A2(n_255), .B1(n_310), .B2(n_311), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_191), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_194), .A2(n_282), .B1(n_364), .B2(n_600), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_195), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_196), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_198), .A2(n_266), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_199), .A2(n_232), .B1(n_364), .B2(n_467), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_204), .Y(n_400) );
INVx1_ASAP7_75t_L g775 ( .A(n_205), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_206), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_207), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_209), .A2(n_851), .B1(n_877), .B2(n_878), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_209), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_210), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_211), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_212), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_213), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_214), .A2(n_250), .B1(n_569), .B2(n_570), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g597 ( .A1(n_215), .A2(n_280), .B1(n_390), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_216), .A2(n_219), .B1(n_413), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_218), .A2(n_251), .B1(n_382), .B2(n_785), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_220), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_222), .B(n_438), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_224), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_230), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_235), .Y(n_856) );
AOI22x1_ASAP7_75t_L g661 ( .A1(n_236), .A2(n_662), .B1(n_691), .B2(n_692), .Y(n_661) );
INVx1_ASAP7_75t_L g691 ( .A(n_236), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g845 ( .A(n_237), .B(n_846), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_239), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g303 ( .A(n_240), .Y(n_303) );
OA22x2_ASAP7_75t_L g634 ( .A1(n_241), .A2(n_635), .B1(n_636), .B2(n_659), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_241), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_242), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_243), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_244), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_247), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_248), .A2(n_283), .B1(n_384), .B2(n_393), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_254), .Y(n_507) );
INVx1_ASAP7_75t_L g844 ( .A(n_255), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_257), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_258), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_259), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_260), .B(n_432), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_261), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_263), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_264), .Y(n_728) );
INVx1_ASAP7_75t_L g310 ( .A(n_270), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_270), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_271), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_272), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_273), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_275), .B(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_276), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_281), .Y(n_639) );
INVx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_290), .Y(n_840) );
OA21x2_ASAP7_75t_L g887 ( .A1(n_291), .A2(n_839), .B(n_888), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_720), .B1(n_834), .B2(n_835), .C(n_836), .Y(n_295) );
INVxp67_ASAP7_75t_L g834 ( .A(n_296), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B1(n_525), .B2(n_719), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_395), .B1(n_523), .B2(n_524), .Y(n_298) );
INVx2_ASAP7_75t_L g523 ( .A(n_299), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_359), .Y(n_300) );
NOR3xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_326), .C(n_346), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B1(n_320), .B2(n_321), .Y(n_302) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g614 ( .A(n_306), .Y(n_614) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_306), .Y(n_727) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_315), .Y(n_306) );
INVx2_ASAP7_75t_L g385 ( .A(n_307), .Y(n_385) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_313), .Y(n_307) );
AND2x2_ASAP7_75t_L g325 ( .A(n_308), .B(n_313), .Y(n_325) );
AND2x2_ASAP7_75t_L g366 ( .A(n_308), .B(n_345), .Y(n_366) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g329 ( .A(n_309), .B(n_313), .Y(n_329) );
AND2x2_ASAP7_75t_L g339 ( .A(n_309), .B(n_319), .Y(n_339) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_312), .Y(n_314) );
INVx2_ASAP7_75t_L g345 ( .A(n_313), .Y(n_345) );
INVx1_ASAP7_75t_L g379 ( .A(n_313), .Y(n_379) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_316), .B(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g388 ( .A(n_316), .B(n_366), .Y(n_388) );
AND2x4_ASAP7_75t_L g435 ( .A(n_316), .B(n_385), .Y(n_435) );
AND2x6_ASAP7_75t_L g438 ( .A(n_316), .B(n_325), .Y(n_438) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g331 ( .A(n_317), .Y(n_331) );
INVx1_ASAP7_75t_L g338 ( .A(n_317), .Y(n_338) );
INVx1_ASAP7_75t_L g358 ( .A(n_317), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_317), .B(n_319), .Y(n_370) );
AND2x2_ASAP7_75t_L g330 ( .A(n_318), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g376 ( .A(n_319), .B(n_358), .Y(n_376) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_323), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_612) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_323), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
BUFx3_ASAP7_75t_L g857 ( .A(n_323), .Y(n_857) );
BUFx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g672 ( .A(n_324), .Y(n_672) );
AND2x2_ASAP7_75t_L g375 ( .A(n_325), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g391 ( .A(n_325), .B(n_330), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_325), .B(n_376), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_332), .B1(n_333), .B2(n_340), .C(n_341), .Y(n_326) );
OAI221xp5_ASAP7_75t_L g664 ( .A1(n_327), .A2(n_640), .B1(n_665), .B2(n_666), .C(n_667), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_327), .A2(n_700), .B(n_701), .Y(n_699) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx4_ASAP7_75t_L g448 ( .A(n_328), .Y(n_448) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_328), .Y(n_483) );
BUFx3_ASAP7_75t_L g549 ( .A(n_328), .Y(n_549) );
INVx2_ASAP7_75t_SL g733 ( .A(n_328), .Y(n_733) );
AND2x6_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g355 ( .A(n_329), .Y(n_355) );
AND2x4_ASAP7_75t_L g495 ( .A(n_329), .B(n_357), .Y(n_495) );
AND2x2_ASAP7_75t_L g365 ( .A(n_330), .B(n_366), .Y(n_365) );
AND2x6_ASAP7_75t_L g384 ( .A(n_330), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g801 ( .A(n_335), .Y(n_801) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx12f_ASAP7_75t_L g451 ( .A(n_336), .Y(n_451) );
INVx1_ASAP7_75t_L g487 ( .A(n_336), .Y(n_487) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_336), .Y(n_509) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g344 ( .A(n_338), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g343 ( .A(n_339), .B(n_344), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g349 ( .A(n_339), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g492 ( .A(n_339), .B(n_493), .Y(n_492) );
INVx4_ASAP7_75t_L g760 ( .A(n_342), .Y(n_760) );
BUFx2_ASAP7_75t_L g828 ( .A(n_342), .Y(n_828) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx4f_ASAP7_75t_SL g449 ( .A(n_343), .Y(n_449) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_343), .Y(n_552) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_343), .Y(n_641) );
INVx1_ASAP7_75t_L g350 ( .A(n_345), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_351), .B2(n_352), .Y(n_346) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx4_ASAP7_75t_L g442 ( .A(n_349), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_349), .A2(n_354), .B1(n_620), .B2(n_621), .Y(n_619) );
BUFx3_ASAP7_75t_L g737 ( .A(n_349), .Y(n_737) );
OAI22xp33_ASAP7_75t_SL g862 ( .A1(n_349), .A2(n_352), .B1(n_863), .B2(n_864), .Y(n_862) );
AND2x2_ASAP7_75t_L g504 ( .A(n_350), .B(n_369), .Y(n_504) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_352), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_352), .A2(n_675), .B1(n_803), .B2(n_804), .Y(n_802) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g677 ( .A(n_353), .Y(n_677) );
CKINVDCx16_ASAP7_75t_R g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g444 ( .A(n_354), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g899 ( .A1(n_354), .A2(n_737), .B1(n_900), .B2(n_901), .Y(n_899) );
OR2x6_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_380), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_371), .Y(n_360) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g472 ( .A(n_364), .Y(n_472) );
BUFx3_ASAP7_75t_L g743 ( .A(n_364), .Y(n_743) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_SL g426 ( .A(n_365), .Y(n_426) );
BUFx2_ASAP7_75t_SL g574 ( .A(n_365), .Y(n_574) );
INVx2_ASAP7_75t_L g625 ( .A(n_365), .Y(n_625) );
AND2x4_ASAP7_75t_L g368 ( .A(n_366), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g394 ( .A(n_366), .B(n_376), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_366), .B(n_376), .Y(n_430) );
BUFx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g406 ( .A(n_368), .Y(n_406) );
INVx1_ASAP7_75t_L g463 ( .A(n_368), .Y(n_463) );
BUFx3_ASAP7_75t_L g518 ( .A(n_368), .Y(n_518) );
BUFx3_ASAP7_75t_L g540 ( .A(n_368), .Y(n_540) );
BUFx2_ASAP7_75t_SL g747 ( .A(n_368), .Y(n_747) );
BUFx2_ASAP7_75t_L g773 ( .A(n_368), .Y(n_773) );
BUFx3_ASAP7_75t_L g815 ( .A(n_368), .Y(n_815) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR2x6_ASAP7_75t_L g378 ( .A(n_370), .B(n_379), .Y(n_378) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g478 ( .A(n_373), .Y(n_478) );
BUFx2_ASAP7_75t_L g770 ( .A(n_373), .Y(n_770) );
INVx4_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g534 ( .A(n_374), .Y(n_534) );
INVx3_ASAP7_75t_L g600 ( .A(n_374), .Y(n_600) );
INVx5_ASAP7_75t_L g628 ( .A(n_374), .Y(n_628) );
INVx1_ASAP7_75t_L g654 ( .A(n_374), .Y(n_654) );
INVx8_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx6_ASAP7_75t_SL g414 ( .A(n_378), .Y(n_414) );
INVx1_ASAP7_75t_SL g479 ( .A(n_378), .Y(n_479) );
INVx1_ASAP7_75t_SL g578 ( .A(n_378), .Y(n_578) );
INVx1_ASAP7_75t_L g493 ( .A(n_379), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_389), .Y(n_380) );
INVx1_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
INVx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx4_ASAP7_75t_L g538 ( .A(n_383), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_383), .B(n_580), .Y(n_579) );
INVx11_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx11_ASAP7_75t_L g468 ( .A(n_384), .Y(n_468) );
BUFx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx3_ASAP7_75t_L g403 ( .A(n_388), .Y(n_403) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_388), .Y(n_475) );
BUFx3_ASAP7_75t_L g626 ( .A(n_388), .Y(n_626) );
INVx2_ASAP7_75t_L g790 ( .A(n_388), .Y(n_790) );
BUFx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx6_ASAP7_75t_L g422 ( .A(n_391), .Y(n_422) );
BUFx3_ASAP7_75t_L g569 ( .A(n_391), .Y(n_569) );
BUFx3_ASAP7_75t_L g690 ( .A(n_391), .Y(n_690) );
BUFx4f_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g750 ( .A(n_393), .Y(n_750) );
BUFx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx3_ASAP7_75t_L g532 ( .A(n_394), .Y(n_532) );
BUFx3_ASAP7_75t_L g571 ( .A(n_394), .Y(n_571) );
BUFx3_ASAP7_75t_L g586 ( .A(n_394), .Y(n_586) );
INVx1_ASAP7_75t_L g524 ( .A(n_395), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_454), .B1(n_521), .B2(n_522), .Y(n_395) );
INVx1_ASAP7_75t_L g522 ( .A(n_396), .Y(n_522) );
INVx1_ASAP7_75t_L g453 ( .A(n_397), .Y(n_453) );
AND4x1_ASAP7_75t_L g397 ( .A(n_398), .B(n_415), .C(n_431), .D(n_445), .Y(n_397) );
NOR2xp33_ASAP7_75t_SL g398 ( .A(n_399), .B(n_407), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_404), .B2(n_405), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_411), .B2(n_412), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g575 ( .A1(n_409), .A2(n_576), .B(n_577), .Y(n_575) );
BUFx2_ASAP7_75t_R g409 ( .A(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g535 ( .A(n_414), .Y(n_535) );
BUFx4f_ASAP7_75t_SL g792 ( .A(n_414), .Y(n_792) );
BUFx2_ASAP7_75t_L g826 ( .A(n_414), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_423), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_420), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_869) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g469 ( .A(n_422), .Y(n_469) );
INVx3_ASAP7_75t_L g785 ( .A(n_422), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_427), .B2(n_428), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g872 ( .A(n_429), .Y(n_872) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx5_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g497 ( .A(n_434), .Y(n_497) );
INVx2_ASAP7_75t_L g543 ( .A(n_434), .Y(n_543) );
INVx2_ASAP7_75t_L g704 ( .A(n_434), .Y(n_704) );
INVx4_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g763 ( .A(n_437), .Y(n_763) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_438), .Y(n_544) );
BUFx2_ASAP7_75t_L g566 ( .A(n_438), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_443), .B2(n_444), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_SL g675 ( .A(n_442), .Y(n_675) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI222xp33_ASAP7_75t_L g638 ( .A1(n_447), .A2(n_639), .B1(n_640), .B2(n_642), .C1(n_643), .C2(n_645), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g797 ( .A1(n_447), .A2(n_640), .B1(n_798), .B2(n_799), .C(n_800), .Y(n_797) );
BUFx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_448), .A2(n_507), .B(n_508), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_448), .A2(n_590), .B(n_591), .Y(n_589) );
OAI21xp5_ASAP7_75t_SL g756 ( .A1(n_448), .A2(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g485 ( .A(n_449), .Y(n_485) );
BUFx4f_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g830 ( .A(n_451), .Y(n_830) );
INVx2_ASAP7_75t_L g521 ( .A(n_454), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_499), .B2(n_520), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g498 ( .A(n_458), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_480), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_470), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_464), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_463), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_873) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx5_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g598 ( .A(n_468), .Y(n_598) );
INVx1_ASAP7_75t_L g657 ( .A(n_468), .Y(n_657) );
INVx2_ASAP7_75t_L g814 ( .A(n_468), .Y(n_814) );
INVx4_ASAP7_75t_L g908 ( .A(n_468), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_476), .Y(n_470) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_489), .Y(n_480) );
OAI222xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B1(n_485), .B2(n_486), .C1(n_487), .C2(n_488), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g559 ( .A(n_483), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_496), .Y(n_489) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx3_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
BUFx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_495), .Y(n_510) );
BUFx2_ASAP7_75t_SL g766 ( .A(n_495), .Y(n_766) );
INVx3_ASAP7_75t_L g520 ( .A(n_499), .Y(n_520) );
XOR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_519), .Y(n_499) );
NAND3x1_ASAP7_75t_SL g500 ( .A(n_501), .B(n_505), .C(n_515), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
NOR2x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
BUFx4f_ASAP7_75t_L g644 ( .A(n_509), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .C(n_514), .Y(n_511) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g682 ( .A(n_518), .Y(n_682) );
INVx1_ASAP7_75t_L g719 ( .A(n_525), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B1(n_605), .B2(n_718), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_553), .B1(n_554), .B2(n_604), .Y(n_527) );
INVx1_ASAP7_75t_SL g604 ( .A(n_528), .Y(n_604) );
NOR4xp75_ASAP7_75t_L g529 ( .A(n_530), .B(n_536), .C(n_541), .D(n_547), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_531), .B(n_533), .Y(n_530) );
BUFx3_ASAP7_75t_L g651 ( .A(n_532), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_537), .B(n_539), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_542), .B(n_545), .Y(n_541) );
OAI21xp5_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_550), .B(n_551), .Y(n_547) );
OAI21xp33_ASAP7_75t_SL g859 ( .A1(n_548), .A2(n_860), .B(n_861), .Y(n_859) );
OAI21xp33_ASAP7_75t_L g896 ( .A1(n_548), .A2(n_897), .B(n_898), .Y(n_896) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_552), .Y(n_562) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OAI22x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_581), .B1(n_602), .B2(n_603), .Y(n_554) );
INVx1_ASAP7_75t_L g602 ( .A(n_555), .Y(n_602) );
NAND3x1_ASAP7_75t_L g556 ( .A(n_557), .B(n_567), .C(n_573), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_563), .Y(n_557) );
OAI21xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_560), .B(n_561), .Y(n_558) );
INVx2_ASAP7_75t_SL g731 ( .A(n_562), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .Y(n_567) );
BUFx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g603 ( .A(n_581), .Y(n_603) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
XOR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_601), .Y(n_582) );
NAND3x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_588), .C(n_596), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .C(n_595), .Y(n_592) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g718 ( .A(n_605), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B1(n_632), .B2(n_717), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND3x1_ASAP7_75t_L g610 ( .A(n_611), .B(n_622), .C(n_629), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_616), .C(n_619), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_614), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_614), .A2(n_671), .B1(n_795), .B2(n_796), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_614), .A2(n_671), .B1(n_894), .B2(n_895), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_627), .Y(n_622) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx3_ASAP7_75t_L g817 ( .A(n_625), .Y(n_817) );
INVx1_ASAP7_75t_L g875 ( .A(n_626), .Y(n_875) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_628), .Y(n_684) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g717 ( .A(n_632), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B1(n_660), .B2(n_716), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g659 ( .A(n_636), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_649), .C(n_655), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_646), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_641), .Y(n_640) );
OAI222xp33_ASAP7_75t_L g730 ( .A1(n_643), .A2(n_731), .B1(n_732), .B2(n_733), .C1(n_734), .C2(n_735), .Y(n_730) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g716 ( .A(n_660), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_693), .B1(n_694), .B2(n_715), .Y(n_660) );
INVx1_ASAP7_75t_L g715 ( .A(n_661), .Y(n_715) );
INVx2_ASAP7_75t_SL g692 ( .A(n_662), .Y(n_692) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_678), .Y(n_662) );
NOR3xp33_ASAP7_75t_SL g663 ( .A(n_664), .B(n_668), .C(n_673), .Y(n_663) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g820 ( .A(n_672), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_673) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_685), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_683), .Y(n_679) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx3_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
XOR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_714), .Y(n_696) );
NAND2x1p5_ASAP7_75t_L g697 ( .A(n_698), .B(n_707), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .C(n_706), .Y(n_702) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g835 ( .A(n_720), .Y(n_835) );
AOI22xp5_ASAP7_75t_SL g720 ( .A1(n_721), .A2(n_777), .B1(n_778), .B2(n_833), .Y(n_720) );
INVx1_ASAP7_75t_L g833 ( .A(n_721), .Y(n_833) );
OAI22xp5_ASAP7_75t_SL g721 ( .A1(n_722), .A2(n_751), .B1(n_752), .B2(n_776), .Y(n_721) );
INVx2_ASAP7_75t_L g776 ( .A(n_722), .Y(n_776) );
XNOR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_740), .Y(n_724) );
NOR3xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_730), .C(n_736), .Y(n_725) );
INVx1_ASAP7_75t_L g855 ( .A(n_727), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_745), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_748), .Y(n_745) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
XOR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_775), .Y(n_753) );
NAND3x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_767), .C(n_771), .Y(n_754) );
NOR2x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_761), .Y(n_755) );
INVx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_764), .C(n_765), .Y(n_761) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_807), .B1(n_808), .B2(n_832), .Y(n_779) );
INVx1_ASAP7_75t_L g832 ( .A(n_780), .Y(n_832) );
INVx1_ASAP7_75t_SL g806 ( .A(n_781), .Y(n_806) );
AND2x2_ASAP7_75t_SL g781 ( .A(n_782), .B(n_793), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_787), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_786), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_791), .Y(n_787) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR3xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_797), .C(n_802), .Y(n_793) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
XOR2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_831), .Y(n_810) );
NAND4xp75_ASAP7_75t_L g811 ( .A(n_812), .B(n_818), .C(n_823), .D(n_827), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_816), .Y(n_812) );
OA211x2_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_820), .B(n_821), .C(n_822), .Y(n_818) );
AND2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
INVx3_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
NOR2x1_ASAP7_75t_L g837 ( .A(n_838), .B(n_842), .Y(n_837) );
OR2x2_ASAP7_75t_SL g910 ( .A(n_838), .B(n_843), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_841), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g881 ( .A(n_839), .Y(n_881) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_840), .B(n_884), .Y(n_888) );
CKINVDCx16_ASAP7_75t_R g884 ( .A(n_841), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_843), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
OAI322xp33_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_879), .A3(n_882), .B1(n_885), .B2(n_889), .C1(n_890), .C2(n_910), .Y(n_849) );
INVx2_ASAP7_75t_L g878 ( .A(n_851), .Y(n_878) );
AND2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_865), .Y(n_851) );
NOR3xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_859), .C(n_862), .Y(n_852) );
OAI22xp5_ASAP7_75t_SL g853 ( .A1(n_854), .A2(n_856), .B1(n_857), .B2(n_858), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NOR3xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_869), .C(n_873), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_886), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_887), .Y(n_886) );
XOR2x2_ASAP7_75t_L g890 ( .A(n_889), .B(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_902), .Y(n_891) );
NOR3xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_896), .C(n_899), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_906), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_904), .B(n_905), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_909), .Y(n_906) );
endmodule