module real_jpeg_17077_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_1),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_1),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_1),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_1),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_2),
.A2(n_196),
.B1(n_201),
.B2(n_205),
.Y(n_195)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_2),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_3),
.A2(n_136),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_3),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_4),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_4),
.A2(n_62),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_4),
.A2(n_62),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_4),
.A2(n_62),
.B1(n_412),
.B2(n_415),
.Y(n_411)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_5),
.A2(n_173),
.B1(n_178),
.B2(n_179),
.Y(n_172)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_5),
.A2(n_178),
.B1(n_213),
.B2(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_5),
.A2(n_178),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_6),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_6),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_6),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_7),
.Y(n_90)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_7),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_7),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_8),
.A2(n_141),
.B1(n_145),
.B2(n_147),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_8),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_8),
.A2(n_147),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_9),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_9),
.A2(n_52),
.B1(n_212),
.B2(n_217),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_9),
.A2(n_52),
.B1(n_362),
.B2(n_365),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_9),
.A2(n_52),
.B1(n_427),
.B2(n_430),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_10),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_10),
.A2(n_116),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_10),
.Y(n_304)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_10),
.A2(n_319),
.A3(n_328),
.B1(n_332),
.B2(n_334),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_10),
.A2(n_304),
.B1(n_374),
.B2(n_378),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_10),
.B(n_99),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_10),
.A2(n_120),
.B1(n_451),
.B2(n_459),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_11),
.A2(n_41),
.B1(n_45),
.B2(n_47),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_11),
.A2(n_47),
.B1(n_290),
.B2(n_294),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_11),
.A2(n_47),
.B1(n_189),
.B2(n_407),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_11),
.A2(n_47),
.B1(n_452),
.B2(n_455),
.Y(n_451)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_12),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_12),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_12),
.A2(n_134),
.B1(n_185),
.B2(n_189),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_13),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_15),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_15),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_15),
.A2(n_95),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_15),
.A2(n_95),
.B1(n_338),
.B2(n_342),
.Y(n_337)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_16),
.Y(n_128)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_16),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g204 ( 
.A(n_16),
.Y(n_204)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_17),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_238),
.CI(n_278),
.CON(n_18),
.SN(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_148),
.C(n_209),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_20),
.B(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_103),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_56),
.B1(n_101),
.B2(n_102),
.Y(n_21)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_40),
.B1(n_48),
.B2(n_49),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_23),
.A2(n_40),
.B1(n_48),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_23),
.A2(n_48),
.B1(n_49),
.B2(n_268),
.Y(n_267)
);

AO21x2_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_33),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_24),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_25),
.Y(n_228)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AO22x2_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_36),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_38),
.Y(n_295)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_43),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_46),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_48),
.B(n_304),
.Y(n_303)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_56),
.B(n_101),
.C(n_103),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_67),
.B1(n_92),
.B2(n_99),
.Y(n_56)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_57),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_60),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_61),
.Y(n_380)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g222 ( 
.A(n_67),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_75),
.B(n_81),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_74),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_75),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_79),
.Y(n_221)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_80),
.Y(n_293)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_80),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_88),
.B2(n_91),
.Y(n_81)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_87),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_87),
.Y(n_364)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_90),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g405 ( 
.A(n_90),
.Y(n_405)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_92),
.Y(n_273)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_100),
.A2(n_211),
.B1(n_222),
.B2(n_223),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_100),
.A2(n_222),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_100),
.A2(n_211),
.B1(n_222),
.B2(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_100),
.A2(n_222),
.B1(n_289),
.B2(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_119),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_104),
.B(n_119),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_111),
.B(n_116),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_129),
.B1(n_137),
.B2(n_140),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_120),
.A2(n_140),
.B1(n_195),
.B2(n_206),
.Y(n_194)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_120),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_120),
.A2(n_258),
.B1(n_411),
.B2(n_416),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_120),
.A2(n_426),
.B1(n_451),
.B2(n_463),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_121),
.A2(n_130),
.B1(n_255),
.B2(n_298),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_121),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_123),
.Y(n_465)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_124),
.Y(n_259)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_127),
.Y(n_429)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_128),
.Y(n_262)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_128),
.Y(n_302)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_128),
.Y(n_399)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_133),
.Y(n_433)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_139),
.Y(n_449)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_143),
.Y(n_300)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_143),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_148),
.B(n_209),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_193),
.B2(n_194),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_149),
.B(n_194),
.Y(n_265)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_172),
.B1(n_182),
.B2(n_184),
.Y(n_150)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_151),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_151),
.B(n_184),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_151),
.A2(n_182),
.B1(n_316),
.B2(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_151),
.A2(n_182),
.B1(n_402),
.B2(n_406),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_151),
.A2(n_182),
.B1(n_361),
.B2(n_406),
.Y(n_420)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_162),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_156),
.B1(n_157),
.B2(n_160),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_157),
.Y(n_344)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_158),
.Y(n_445)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_159),
.Y(n_389)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_159),
.Y(n_454)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_167),
.B2(n_171),
.Y(n_162)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_169),
.Y(n_391)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_175),
.Y(n_333)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_177),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_177),
.Y(n_408)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_182),
.B(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_183),
.A2(n_230),
.B1(n_231),
.B2(n_237),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_183),
.A2(n_230),
.B1(n_231),
.B2(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_183),
.B(n_304),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_200),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_203),
.Y(n_458)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_204),
.Y(n_414)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_224),
.C(n_229),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_210),
.B(n_229),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_224),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_264),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_254),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_253),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_260),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_255),
.A2(n_298),
.B1(n_337),
.B2(n_345),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_255),
.A2(n_425),
.B1(n_434),
.B2(n_435),
.Y(n_424)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

INVx3_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_305),
.B(n_478),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_281),
.B(n_283),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.C(n_287),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_287),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_296),
.C(n_303),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_288),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_297),
.B1(n_303),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_304),
.B(n_393),
.Y(n_392)
);

OAI21xp33_ASAP7_75t_SL g402 ( 
.A1(n_304),
.A2(n_392),
.B(n_403),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_304),
.B(n_447),
.Y(n_446)
);

AOI21x1_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_351),
.B(n_477),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_307),
.B(n_309),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.C(n_325),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_310),
.A2(n_311),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_314),
.A2(n_325),
.B1(n_326),
.B2(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_323),
.Y(n_387)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_335),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_327),
.A2(n_335),
.B1(n_336),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_350),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_381),
.B(n_476),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_353),
.B(n_357),
.Y(n_476)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.C(n_371),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_358),
.B(n_473),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_360),
.A2(n_371),
.B1(n_372),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_360),
.Y(n_474)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_369),
.Y(n_393)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI21x1_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_470),
.B(n_475),
.Y(n_381)
);

OAI21x1_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_422),
.B(n_469),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_409),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_384),
.B(n_409),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_400),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_385),
.A2(n_400),
.B1(n_401),
.B2(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_385),
.Y(n_437)
);

OAI32xp33_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_388),
.A3(n_390),
.B1(n_392),
.B2(n_394),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_390),
.Y(n_395)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_417),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_410),
.B(n_419),
.C(n_421),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_411),
.Y(n_435)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_417)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_418),
.Y(n_421)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_438),
.B(n_468),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_436),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_424),
.B(n_436),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_461),
.B(n_467),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_450),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_446),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_466),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_466),
.Y(n_467)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_SL g475 ( 
.A(n_471),
.B(n_472),
.Y(n_475)
);


endmodule