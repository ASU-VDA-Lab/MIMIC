module fake_jpeg_13046_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_13),
.B1(n_33),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_34),
.B1(n_31),
.B2(n_26),
.Y(n_51)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_1),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_21),
.B1(n_20),
.B2(n_15),
.Y(n_55)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_50),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_64),
.B1(n_56),
.B2(n_58),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_37),
.B(n_3),
.C(n_4),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_5),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_44),
.B(n_43),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_40),
.B1(n_44),
.B2(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_78),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_39),
.B(n_36),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_1),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_37),
.B1(n_11),
.B2(n_4),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_70),
.B1(n_6),
.B2(n_7),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_2),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_5),
.C(n_6),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_2),
.Y(n_88)
);

OAI221xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.C(n_8),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_82),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_70),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_98),
.Y(n_105)
);

XNOR2x1_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_7),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_85),
.Y(n_102)
);

AOI21x1_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_81),
.B(n_91),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_96),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_103),
.A2(n_104),
.B(n_93),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_107),
.B(n_105),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_99),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_104),
.B(n_97),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_93),
.B1(n_100),
.B2(n_94),
.C(n_80),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_8),
.Y(n_112)
);


endmodule