module fake_jpeg_821_n_714 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_714);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_714;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_60),
.Y(n_169)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_63),
.B(n_69),
.Y(n_148)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_20),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_70),
.B(n_75),
.Y(n_153)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_79),
.B(n_88),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_80),
.Y(n_201)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_42),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_82),
.A2(n_58),
.B1(n_28),
.B2(n_25),
.Y(n_178)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_83),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_55),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_84),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_29),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_87),
.Y(n_154)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_24),
.B(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_89),
.Y(n_212)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_91),
.B(n_92),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_38),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_94),
.Y(n_202)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_97),
.B(n_116),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_26),
.B(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_98),
.B(n_133),
.Y(n_220)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_100),
.Y(n_197)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_103),
.Y(n_171)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx6_ASAP7_75t_SL g106 ( 
.A(n_24),
.Y(n_106)
);

BUFx16f_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_44),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_112),
.Y(n_226)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_24),
.Y(n_113)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_52),
.Y(n_118)
);

NAND2x1_ASAP7_75t_SL g166 ( 
.A(n_118),
.B(n_23),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_47),
.Y(n_120)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_49),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_123),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_49),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_22),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_27),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_22),
.Y(n_127)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_31),
.Y(n_128)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_128),
.Y(n_228)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_31),
.Y(n_129)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_23),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_23),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_31),
.Y(n_132)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_26),
.B(n_50),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_135),
.B(n_182),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_65),
.A2(n_54),
.B1(n_53),
.B2(n_40),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_145),
.A2(n_184),
.B1(n_0),
.B2(n_3),
.Y(n_271)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_162),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_120),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_163),
.B(n_183),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_166),
.B(n_232),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_84),
.B(n_27),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_173),
.Y(n_315)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_177),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_178),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_290)
);

BUFx4f_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_179),
.Y(n_245)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_62),
.B(n_36),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_94),
.A2(n_101),
.B1(n_117),
.B2(n_118),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_62),
.B(n_36),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_187),
.B(n_189),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_93),
.B(n_41),
.Y(n_189)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_90),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g276 ( 
.A(n_190),
.Y(n_276)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_73),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_111),
.B(n_41),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_218),
.Y(n_243)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_90),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_205),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_126),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_208),
.B(n_0),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_81),
.Y(n_210)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_210),
.Y(n_310)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_96),
.Y(n_211)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

BUFx2_ASAP7_75t_R g214 ( 
.A(n_124),
.Y(n_214)
);

INVx5_ASAP7_75t_SL g246 ( 
.A(n_214),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_100),
.Y(n_216)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_216),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_67),
.B(n_43),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_82),
.A2(n_48),
.B(n_43),
.C(n_32),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_219),
.B(n_222),
.Y(n_280)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_131),
.B(n_48),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_66),
.Y(n_224)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_108),
.B(n_50),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_229),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_124),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_227),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_130),
.B(n_32),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_96),
.B(n_57),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_18),
.Y(n_269)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_68),
.Y(n_231)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_72),
.A2(n_57),
.B1(n_40),
.B2(n_54),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_74),
.Y(n_233)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_237),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_171),
.A2(n_25),
.B1(n_28),
.B2(n_58),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_238),
.A2(n_239),
.B1(n_256),
.B2(n_257),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_171),
.A2(n_25),
.B1(n_28),
.B2(n_58),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_240),
.Y(n_322)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_242),
.Y(n_366)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_244),
.Y(n_375)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_139),
.Y(n_247)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_247),
.Y(n_329)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_200),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_180),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_249),
.B(n_252),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_169),
.B(n_119),
.C(n_114),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_250),
.B(n_265),
.C(n_304),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_174),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_112),
.B1(n_109),
.B2(n_80),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_253),
.A2(n_255),
.B1(n_302),
.B2(n_319),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_145),
.A2(n_86),
.B1(n_102),
.B2(n_54),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_199),
.A2(n_102),
.B1(n_53),
.B2(n_40),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_199),
.A2(n_53),
.B1(n_35),
.B2(n_5),
.Y(n_257)
);

INVx3_ASAP7_75t_SL g261 ( 
.A(n_200),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_173),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_263),
.B(n_284),
.Y(n_359)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_139),
.Y(n_264)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_175),
.B(n_35),
.C(n_19),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_207),
.A2(n_35),
.B1(n_3),
.B2(n_5),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_266),
.A2(n_290),
.B1(n_292),
.B2(n_297),
.Y(n_351)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_186),
.Y(n_267)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_212),
.Y(n_268)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_269),
.B(n_295),
.Y(n_341)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_270),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_271),
.A2(n_150),
.B1(n_160),
.B2(n_158),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_206),
.B(n_17),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_273),
.B(n_307),
.Y(n_358)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_137),
.Y(n_275)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_161),
.Y(n_277)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_142),
.Y(n_279)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_142),
.Y(n_281)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g377 ( 
.A(n_282),
.Y(n_377)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_198),
.Y(n_283)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_283),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_148),
.B(n_3),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_153),
.B(n_5),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_R g321 ( 
.A(n_285),
.B(n_303),
.Y(n_321)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_164),
.Y(n_286)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_286),
.Y(n_361)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_167),
.Y(n_287)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_287),
.Y(n_367)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_147),
.Y(n_288)
);

INVx11_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_184),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_216),
.Y(n_293)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_293),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_154),
.B(n_8),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_161),
.Y(n_296)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_143),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_192),
.B(n_11),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_299),
.B(n_305),
.Y(n_365)
);

BUFx12f_ASAP7_75t_L g300 ( 
.A(n_147),
.Y(n_300)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

CKINVDCx12_ASAP7_75t_R g301 ( 
.A(n_190),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_144),
.A2(n_146),
.B1(n_203),
.B2(n_202),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_151),
.B(n_11),
.Y(n_303)
);

AND2x2_ASAP7_75t_SL g304 ( 
.A(n_215),
.B(n_12),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_213),
.B(n_15),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_210),
.Y(n_306)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_166),
.B(n_15),
.Y(n_307)
);

OR2x2_ASAP7_75t_SL g308 ( 
.A(n_228),
.B(n_16),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_308),
.B(n_191),
.C(n_141),
.Y(n_382)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_210),
.Y(n_311)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_311),
.Y(n_338)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_168),
.Y(n_312)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_217),
.B(n_157),
.Y(n_313)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_313),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_156),
.B(n_16),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_304),
.Y(n_323)
);

CKINVDCx12_ASAP7_75t_R g316 ( 
.A(n_149),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_316),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_193),
.B(n_136),
.Y(n_317)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_176),
.Y(n_318)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_318),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_202),
.A2(n_203),
.B1(n_172),
.B2(n_196),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_323),
.B(n_273),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_251),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_326),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_280),
.A2(n_172),
.B1(n_196),
.B2(n_152),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_328),
.A2(n_352),
.B1(n_360),
.B2(n_372),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_243),
.B(n_170),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_332),
.B(n_254),
.C(n_246),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_251),
.B(n_215),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_337),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_292),
.A2(n_204),
.B1(n_138),
.B2(n_209),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_342),
.A2(n_376),
.B1(n_246),
.B2(n_291),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_136),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_256),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_235),
.B(n_179),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_346),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_262),
.B(n_176),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_348),
.B(n_355),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_315),
.A2(n_152),
.B1(n_143),
.B2(n_226),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_272),
.B(n_197),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_274),
.B(n_197),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_258),
.A2(n_226),
.B1(n_223),
.B2(n_160),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_255),
.A2(n_223),
.B1(n_150),
.B2(n_201),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_362),
.A2(n_368),
.B1(n_279),
.B2(n_211),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_248),
.B(n_149),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_363),
.Y(n_415)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_245),
.Y(n_369)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_369),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_278),
.A2(n_201),
.B1(n_158),
.B2(n_204),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_241),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_379),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_250),
.A2(n_209),
.B1(n_191),
.B2(n_134),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_245),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_261),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_382),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_384),
.B(n_406),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_337),
.A2(n_291),
.B1(n_293),
.B2(n_242),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_332),
.B(n_308),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_386),
.B(n_390),
.Y(n_438)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_346),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_388),
.B(n_396),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_431),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_323),
.B(n_266),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_392),
.B(n_393),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_325),
.B(n_309),
.Y(n_393)
);

INVx13_ASAP7_75t_L g395 ( 
.A(n_345),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_395),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_346),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_397),
.A2(n_430),
.B1(n_363),
.B2(n_383),
.Y(n_454)
);

AND2x6_ASAP7_75t_L g398 ( 
.A(n_321),
.B(n_141),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_398),
.B(n_402),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_326),
.B(n_294),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_403),
.C(n_418),
.Y(n_445)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_377),
.Y(n_401)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_401),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_325),
.B(n_309),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_326),
.B(n_234),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_381),
.Y(n_404)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_365),
.B(n_240),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_336),
.B(n_318),
.Y(n_410)
);

NAND3xp33_ASAP7_75t_L g451 ( 
.A(n_410),
.B(n_411),
.C(n_414),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_350),
.B(n_282),
.Y(n_411)
);

INVx13_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_412),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_337),
.A2(n_239),
.B(n_238),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_413),
.A2(n_426),
.B(n_433),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_350),
.B(n_283),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_341),
.B(n_298),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_420),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_234),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_335),
.B(n_264),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_419),
.B(n_421),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_359),
.B(n_298),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_247),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_321),
.B(n_141),
.Y(n_422)
);

OA22x2_ASAP7_75t_L g469 ( 
.A1(n_422),
.A2(n_329),
.B1(n_333),
.B2(n_357),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_364),
.A2(n_236),
.B(n_257),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_423),
.A2(n_294),
.B(n_260),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_311),
.C(n_306),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_363),
.C(n_324),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_320),
.A2(n_275),
.B1(n_244),
.B2(n_281),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_425),
.A2(n_349),
.B1(n_375),
.B2(n_383),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_353),
.B(n_236),
.Y(n_426)
);

INVx13_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_427),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_358),
.B(n_289),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_428),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_344),
.B(n_259),
.Y(n_431)
);

CKINVDCx11_ASAP7_75t_R g432 ( 
.A(n_339),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_347),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_354),
.B(n_289),
.Y(n_433)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_394),
.Y(n_440)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_440),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_392),
.A2(n_320),
.B1(n_362),
.B2(n_351),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_441),
.A2(n_444),
.B1(n_472),
.B2(n_473),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_393),
.A2(n_358),
.B1(n_360),
.B2(n_328),
.Y(n_444)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_447),
.Y(n_499)
);

MAJx2_ASAP7_75t_L g448 ( 
.A(n_402),
.B(n_334),
.C(n_330),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_448),
.B(n_429),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_449),
.B(n_464),
.C(n_476),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_454),
.A2(n_409),
.B1(n_441),
.B2(n_429),
.Y(n_505)
);

OAI32xp33_ASAP7_75t_L g455 ( 
.A1(n_390),
.A2(n_357),
.A3(n_374),
.B1(n_370),
.B2(n_348),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_455),
.B(n_471),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_457),
.Y(n_481)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_460),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_421),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_462),
.B(n_420),
.Y(n_478)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_463),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_324),
.C(n_338),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_407),
.Y(n_466)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_426),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_469),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_468),
.Y(n_490)
);

OAI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_397),
.A2(n_329),
.B1(n_333),
.B2(n_374),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_470),
.A2(n_430),
.B1(n_425),
.B2(n_415),
.Y(n_495)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_405),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_434),
.A2(n_408),
.B1(n_422),
.B2(n_398),
.Y(n_472)
);

OAI22xp33_ASAP7_75t_L g473 ( 
.A1(n_434),
.A2(n_343),
.B1(n_375),
.B2(n_331),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_475),
.A2(n_436),
.B(n_413),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_400),
.B(n_338),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_478),
.B(n_483),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_435),
.B(n_389),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_482),
.B(n_507),
.C(n_448),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_465),
.B(n_417),
.Y(n_483)
);

NOR4xp25_ASAP7_75t_SL g484 ( 
.A(n_472),
.B(n_398),
.C(n_422),
.D(n_416),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_484),
.A2(n_503),
.B(n_509),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_461),
.B(n_391),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_485),
.B(n_493),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_457),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_486),
.B(n_508),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_435),
.B(n_403),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_487),
.B(n_482),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_465),
.Y(n_488)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_418),
.Y(n_492)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_492),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_456),
.B(n_391),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_406),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_494),
.B(n_496),
.Y(n_549)
);

OAI22x1_ASAP7_75t_L g521 ( 
.A1(n_495),
.A2(n_438),
.B1(n_469),
.B2(n_468),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_451),
.B(n_432),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_463),
.B(n_431),
.Y(n_497)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_497),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_437),
.B(n_419),
.Y(n_498)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_498),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_455),
.B(n_396),
.Y(n_500)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_500),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_457),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_502),
.B(n_506),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_505),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_458),
.A2(n_423),
.B1(n_416),
.B2(n_388),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_453),
.B(n_410),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_458),
.A2(n_428),
.B(n_405),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_442),
.B(n_386),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_510),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_444),
.A2(n_424),
.B1(n_429),
.B2(n_414),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_512),
.A2(n_459),
.B1(n_450),
.B2(n_477),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_460),
.B(n_411),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_513),
.B(n_439),
.Y(n_540)
);

MAJx2_ASAP7_75t_L g557 ( 
.A(n_514),
.B(n_356),
.C(n_348),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_464),
.B(n_384),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_517),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_471),
.A2(n_399),
.B1(n_405),
.B2(n_401),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_516),
.A2(n_401),
.B(n_427),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_452),
.B(n_404),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_518),
.B(n_520),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_503),
.A2(n_475),
.B(n_442),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_519),
.A2(n_554),
.B(n_555),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_521),
.A2(n_480),
.B1(n_490),
.B2(n_504),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_485),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_522),
.B(n_531),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_SL g530 ( 
.A1(n_490),
.A2(n_436),
.B1(n_446),
.B2(n_459),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_530),
.A2(n_552),
.B1(n_495),
.B2(n_516),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_481),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_487),
.B(n_445),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_533),
.B(n_535),
.C(n_543),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_445),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_534),
.B(n_506),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_438),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_513),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_538),
.Y(n_561)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_540),
.Y(n_559)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_500),
.A2(n_469),
.B(n_452),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_541),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_488),
.A2(n_509),
.B(n_510),
.Y(n_542)
);

XOR2x1_ASAP7_75t_L g582 ( 
.A(n_542),
.B(n_557),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_492),
.B(n_449),
.C(n_476),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_512),
.B(n_469),
.C(n_447),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_544),
.B(n_545),
.C(n_547),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_439),
.C(n_466),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_493),
.B(n_404),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_546),
.B(n_548),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_502),
.B(n_443),
.C(n_361),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_498),
.B(n_450),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_497),
.B(n_443),
.C(n_361),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_550),
.B(n_501),
.C(n_511),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_551),
.A2(n_521),
.B1(n_545),
.B2(n_553),
.Y(n_584)
);

NOR4xp25_ASAP7_75t_L g552 ( 
.A(n_504),
.B(n_473),
.C(n_427),
.D(n_477),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_501),
.Y(n_553)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_553),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_556),
.A2(n_479),
.B1(n_491),
.B2(n_480),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_558),
.A2(n_565),
.B1(n_577),
.B2(n_592),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_536),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_560),
.B(n_355),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_536),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_563),
.B(n_541),
.Y(n_601)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_564),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_556),
.A2(n_479),
.B1(n_491),
.B2(n_480),
.Y(n_565)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_532),
.Y(n_567)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_567),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_568),
.A2(n_573),
.B1(n_580),
.B2(n_584),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_571),
.B(n_576),
.Y(n_603)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_532),
.Y(n_572)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_572),
.Y(n_602)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_523),
.Y(n_574)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_574),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_538),
.A2(n_490),
.B1(n_484),
.B2(n_499),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_523),
.Y(n_578)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_578),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_518),
.B(n_499),
.C(n_511),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_579),
.B(n_581),
.C(n_591),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_528),
.A2(n_527),
.B1(n_549),
.B2(n_525),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_534),
.B(n_489),
.C(n_481),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_526),
.A2(n_555),
.B1(n_541),
.B2(n_542),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_585),
.A2(n_588),
.B1(n_412),
.B2(n_395),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_539),
.Y(n_598)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_550),
.Y(n_587)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_587),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_551),
.A2(n_489),
.B1(n_331),
.B2(n_322),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_520),
.B(n_322),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_590),
.B(n_327),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_533),
.B(n_543),
.C(n_524),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_529),
.A2(n_539),
.B1(n_524),
.B2(n_519),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_591),
.B(n_547),
.C(n_544),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_594),
.B(n_599),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_569),
.B(n_537),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_595),
.B(n_615),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_598),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_590),
.B(n_537),
.C(n_535),
.Y(n_599)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_601),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_583),
.A2(n_529),
.B(n_554),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_605),
.A2(n_586),
.B(n_592),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_579),
.B(n_557),
.C(n_381),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_606),
.B(n_613),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_607),
.B(n_616),
.Y(n_630)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_608),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_367),
.Y(n_610)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_610),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_566),
.B(n_367),
.Y(n_611)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_611),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_570),
.B(n_366),
.C(n_259),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_581),
.B(n_366),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_614),
.B(n_617),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_569),
.B(n_355),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_561),
.B(n_356),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_570),
.B(n_260),
.C(n_377),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_619),
.B(n_576),
.C(n_575),
.Y(n_624)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_560),
.Y(n_620)
);

NOR3xp33_ASAP7_75t_L g625 ( 
.A(n_620),
.B(n_563),
.C(n_562),
.Y(n_625)
);

BUFx12_ASAP7_75t_L g623 ( 
.A(n_605),
.Y(n_623)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_623),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_624),
.B(n_629),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_625),
.A2(n_628),
.B1(n_635),
.B2(n_644),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_593),
.B(n_575),
.C(n_571),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_627),
.B(n_631),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_612),
.A2(n_584),
.B1(n_573),
.B2(n_583),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_604),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_SL g631 ( 
.A(n_596),
.B(n_582),
.C(n_559),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_632),
.A2(n_639),
.B(n_602),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_618),
.B(n_593),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_633),
.B(n_636),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_612),
.A2(n_588),
.B1(n_558),
.B2(n_565),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_594),
.B(n_577),
.C(n_582),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_598),
.A2(n_412),
.B(n_395),
.Y(n_639)
);

BUFx12_ASAP7_75t_L g640 ( 
.A(n_617),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_640),
.B(n_606),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_603),
.B(n_343),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_624),
.B(n_603),
.C(n_615),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_645),
.B(n_646),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_627),
.B(n_613),
.C(n_595),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_621),
.A2(n_597),
.B(n_598),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_647),
.B(n_649),
.Y(n_668)
);

HAxp5_ASAP7_75t_L g650 ( 
.A(n_623),
.B(n_616),
.CON(n_650),
.SN(n_650)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_650),
.B(n_653),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_636),
.B(n_599),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_652),
.B(n_654),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_622),
.A2(n_600),
.B1(n_609),
.B2(n_619),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_634),
.B(n_377),
.C(n_340),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_655),
.B(n_658),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_632),
.A2(n_310),
.B(n_140),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_656),
.A2(n_629),
.B(n_300),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_638),
.A2(n_340),
.B1(n_140),
.B2(n_162),
.Y(n_658)
);

FAx1_ASAP7_75t_SL g659 ( 
.A(n_631),
.B(n_310),
.CI(n_177),
.CON(n_659),
.SN(n_659)
);

OAI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_659),
.A2(n_639),
.B1(n_630),
.B2(n_637),
.Y(n_667)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_626),
.B(n_628),
.Y(n_661)
);

XNOR2xp5_ASAP7_75t_L g673 ( 
.A(n_661),
.B(n_663),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_641),
.B(n_276),
.C(n_188),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_662),
.B(n_641),
.C(n_637),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_635),
.B(n_300),
.Y(n_663)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_665),
.Y(n_682)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_667),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_660),
.B(n_643),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_669),
.B(n_670),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_SL g670 ( 
.A1(n_664),
.A2(n_630),
.B1(n_623),
.B2(n_642),
.Y(n_670)
);

NOR3xp33_ASAP7_75t_L g683 ( 
.A(n_674),
.B(n_662),
.C(n_659),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_661),
.B(n_629),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_676),
.B(n_678),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_SL g677 ( 
.A1(n_650),
.A2(n_629),
.B(n_640),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_677),
.A2(n_656),
.B(n_663),
.Y(n_691)
);

MAJIxp5_ASAP7_75t_L g678 ( 
.A(n_648),
.B(n_645),
.C(n_646),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_648),
.Y(n_679)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_679),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_657),
.B(n_640),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_680),
.B(n_666),
.Y(n_690)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_683),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_671),
.A2(n_653),
.B(n_651),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_685),
.B(n_689),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_675),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_686),
.B(n_690),
.Y(n_693)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_670),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_691),
.A2(n_674),
.B(n_672),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_678),
.B(n_655),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_692),
.B(n_673),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_SL g695 ( 
.A1(n_687),
.A2(n_675),
.B(n_667),
.C(n_668),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_SL g701 ( 
.A(n_695),
.B(n_699),
.C(n_681),
.Y(n_701)
);

XOR2xp5_ASAP7_75t_L g696 ( 
.A(n_684),
.B(n_652),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_696),
.B(n_697),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_682),
.B(n_677),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_SL g705 ( 
.A(n_698),
.B(n_673),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_701),
.A2(n_705),
.B1(n_288),
.B2(n_276),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_694),
.B(n_688),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_702),
.Y(n_708)
);

BUFx24_ASAP7_75t_SL g703 ( 
.A(n_693),
.Y(n_703)
);

AOI322xp5_ASAP7_75t_L g706 ( 
.A1(n_703),
.A2(n_695),
.A3(n_683),
.B1(n_700),
.B2(n_691),
.C1(n_665),
.C2(n_276),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_706),
.B(n_188),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_707),
.A2(n_288),
.B(n_704),
.Y(n_709)
);

OAI321xp33_ASAP7_75t_L g711 ( 
.A1(n_709),
.A2(n_710),
.A3(n_708),
.B1(n_188),
.B2(n_205),
.C(n_149),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_711),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_SL g713 ( 
.A(n_712),
.B(n_185),
.Y(n_713)
);

AOI21x1_ASAP7_75t_L g714 ( 
.A1(n_713),
.A2(n_205),
.B(n_155),
.Y(n_714)
);


endmodule