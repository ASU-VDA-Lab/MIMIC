module fake_jpeg_18480_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_4),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_12),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_66),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx10_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_0),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_61),
.Y(n_75)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_77),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_52),
.B1(n_51),
.B2(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_58),
.B1(n_41),
.B2(n_50),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

HAxp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_60),
.CON(n_81),
.SN(n_81)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_54),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_5),
.B1(n_55),
.B2(n_14),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_2),
.Y(n_98)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_1),
.C(n_2),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_53),
.B1(n_44),
.B2(n_48),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_42),
.B1(n_63),
.B2(n_47),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_56),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_104),
.B(n_28),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_103),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_49),
.C(n_43),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_98),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_5),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_106),
.A2(n_108),
.B1(n_8),
.B2(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_115),
.Y(n_118)
);

INVxp33_ASAP7_75t_SL g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_21),
.B1(n_23),
.B2(n_26),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_114),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_101),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_111),
.C(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_107),
.C(n_115),
.Y(n_122)
);

NAND4xp25_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_120),
.C(n_122),
.D(n_105),
.Y(n_124)
);

OAI21x1_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_105),
.B(n_119),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_116),
.B(n_30),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_29),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_31),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_32),
.C(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_35),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_36),
.Y(n_131)
);


endmodule