module fake_aes_12663_n_719 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_719);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_719;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g107 ( .A(n_50), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_85), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_22), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_97), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_5), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_51), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_63), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_17), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_64), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_79), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_57), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_10), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_69), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_20), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_16), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_59), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_43), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_62), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_32), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_84), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_30), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_103), .Y(n_130) );
CKINVDCx14_ASAP7_75t_R g131 ( .A(n_81), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_41), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_17), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_9), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_36), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_90), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_8), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_49), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_94), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_44), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_95), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_3), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_60), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_12), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_101), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_91), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_19), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_56), .Y(n_149) );
INVxp67_ASAP7_75t_SL g150 ( .A(n_21), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_129), .B(n_0), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_144), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_113), .B(n_0), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_107), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_114), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_114), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_107), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_108), .Y(n_159) );
NAND2xp33_ASAP7_75t_L g160 ( .A(n_114), .B(n_27), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_108), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_112), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g163 ( .A1(n_145), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_112), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_116), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_114), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_113), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_120), .B(n_1), .Y(n_168) );
NAND2xp33_ASAP7_75t_L g169 ( .A(n_114), .B(n_106), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_118), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_157), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_157), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_162), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_162), .Y(n_174) );
BUFx10_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_167), .B(n_140), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_155), .B(n_130), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_162), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_162), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_158), .B(n_132), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_158), .B(n_118), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_170), .Y(n_185) );
NAND3xp33_ASAP7_75t_L g186 ( .A(n_159), .B(n_135), .C(n_116), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_157), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_159), .B(n_121), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_170), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_170), .Y(n_192) );
INVx4_ASAP7_75t_SL g193 ( .A(n_161), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_163), .B(n_117), .Y(n_194) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_152), .B(n_119), .Y(n_195) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_161), .B(n_119), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_173), .A2(n_165), .B(n_164), .Y(n_197) );
NAND2xp33_ASAP7_75t_L g198 ( .A(n_196), .B(n_164), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_179), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_175), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_175), .B(n_167), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_175), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_181), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_181), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_175), .B(n_165), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_185), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_179), .B(n_152), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_195), .B(n_168), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_181), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_185), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_179), .B(n_154), .Y(n_211) );
OR2x2_ASAP7_75t_SL g212 ( .A(n_194), .B(n_115), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_173), .A2(n_169), .B(n_160), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_179), .B(n_154), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_181), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_195), .A2(n_196), .B1(n_186), .B2(n_182), .Y(n_216) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_177), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_177), .B(n_150), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_177), .B(n_168), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_174), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_195), .B(n_126), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_185), .Y(n_222) );
INVxp67_ASAP7_75t_SL g223 ( .A(n_196), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_196), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_186), .A2(n_178), .B1(n_192), .B2(n_191), .Y(n_225) );
O2A1O1Ixp5_ASAP7_75t_L g226 ( .A1(n_184), .A2(n_143), .B(n_135), .C(n_124), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_174), .B(n_131), .Y(n_227) );
OR2x6_ASAP7_75t_L g228 ( .A(n_194), .B(n_163), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_194), .A2(n_137), .B1(n_142), .B2(n_117), .Y(n_229) );
AOI22xp33_ASAP7_75t_SL g230 ( .A1(n_194), .A2(n_137), .B1(n_142), .B2(n_134), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_223), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_220), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_199), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_202), .B(n_193), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_226), .A2(n_180), .B(n_184), .C(n_188), .Y(n_235) );
OR2x6_ASAP7_75t_L g236 ( .A(n_200), .B(n_194), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_205), .A2(n_180), .B(n_188), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_208), .A2(n_194), .B1(n_191), .B2(n_192), .Y(n_238) );
BUFx12f_ASAP7_75t_L g239 ( .A(n_212), .Y(n_239) );
BUFx12f_ASAP7_75t_L g240 ( .A(n_212), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_201), .B(n_109), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_220), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_205), .A2(n_176), .B(n_190), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_223), .A2(n_110), .B1(n_136), .B2(n_123), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_217), .B(n_111), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_202), .Y(n_246) );
NOR2xp33_ASAP7_75t_SL g247 ( .A(n_202), .B(n_193), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_200), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_224), .Y(n_249) );
NAND3xp33_ASAP7_75t_L g250 ( .A(n_226), .B(n_148), .C(n_123), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_217), .A2(n_148), .B(n_133), .C(n_134), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_199), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_224), .B(n_193), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_224), .Y(n_254) );
CKINVDCx6p67_ASAP7_75t_R g255 ( .A(n_201), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_198), .A2(n_176), .B(n_190), .Y(n_256) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_224), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_200), .B(n_193), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_200), .B(n_193), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_219), .A2(n_133), .B(n_122), .C(n_144), .Y(n_260) );
NOR3xp33_ASAP7_75t_SL g261 ( .A(n_208), .B(n_141), .C(n_147), .Y(n_261) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_250), .A2(n_213), .B(n_197), .Y(n_262) );
BUFx10_ASAP7_75t_L g263 ( .A(n_259), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_232), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_256), .A2(n_213), .B(n_197), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_231), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_236), .B(n_219), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_232), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_243), .A2(n_227), .B(n_216), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_242), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_231), .A2(n_216), .B1(n_229), .B2(n_230), .Y(n_271) );
NAND2x1p5_ASAP7_75t_L g272 ( .A(n_248), .B(n_206), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_250), .A2(n_242), .B(n_237), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_246), .Y(n_274) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_235), .A2(n_143), .B(n_146), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_246), .Y(n_276) );
CKINVDCx8_ASAP7_75t_R g277 ( .A(n_248), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_SL g278 ( .A1(n_258), .A2(n_227), .B(n_124), .C(n_146), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_233), .Y(n_279) );
OR2x6_ASAP7_75t_L g280 ( .A(n_236), .B(n_207), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_233), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_238), .A2(n_228), .B1(n_219), .B2(n_230), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_241), .A2(n_207), .B(n_214), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_252), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_234), .A2(n_225), .B(n_121), .Y(n_285) );
AO31x2_ASAP7_75t_L g286 ( .A1(n_252), .A2(n_166), .A3(n_156), .B(n_125), .Y(n_286) );
NAND2x1_ASAP7_75t_L g287 ( .A(n_264), .B(n_246), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_282), .A2(n_228), .B1(n_240), .B2(n_239), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_264), .B(n_255), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_282), .A2(n_228), .B1(n_240), .B2(n_239), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_271), .A2(n_255), .B1(n_236), .B2(n_229), .Y(n_291) );
OAI22xp33_ASAP7_75t_L g292 ( .A1(n_271), .A2(n_228), .B1(n_244), .B2(n_236), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_264), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_266), .B(n_236), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_266), .A2(n_228), .B1(n_249), .B2(n_254), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_270), .Y(n_296) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_285), .A2(n_166), .B(n_156), .Y(n_297) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_285), .A2(n_125), .B(n_138), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_270), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_266), .B(n_218), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_263), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_267), .B(n_218), .Y(n_302) );
NAND2x1p5_ASAP7_75t_L g303 ( .A(n_270), .B(n_246), .Y(n_303) );
OAI22xp33_ASAP7_75t_L g304 ( .A1(n_277), .A2(n_228), .B1(n_249), .B2(n_247), .Y(n_304) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_277), .A2(n_247), .B1(n_254), .B2(n_257), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_279), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_268), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_268), .B(n_218), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_299), .B(n_275), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_293), .B(n_275), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_293), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_289), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_292), .A2(n_283), .B(n_269), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_293), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_296), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_296), .B(n_275), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_296), .B(n_274), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_307), .B(n_267), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_306), .B(n_275), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_307), .B(n_275), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_306), .B(n_279), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_306), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_303), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_289), .B(n_281), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_289), .B(n_281), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_291), .B(n_284), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_301), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_292), .B(n_284), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_303), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_291), .B(n_286), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_298), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_298), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_316), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_316), .B(n_295), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_323), .B(n_295), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_322), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_333), .A2(n_288), .B1(n_290), .B2(n_304), .Y(n_340) );
INVxp67_ASAP7_75t_SL g341 ( .A(n_323), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_328), .Y(n_342) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_323), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_311), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_325), .B(n_298), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_322), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_335), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_335), .A2(n_269), .B(n_283), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_330), .B(n_294), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_325), .B(n_326), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_325), .B(n_298), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_330), .B(n_294), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_334), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_313), .A2(n_285), .B(n_305), .Y(n_355) );
INVx5_ASAP7_75t_SL g356 ( .A(n_318), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_334), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_311), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_309), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_319), .B(n_218), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_327), .B(n_308), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_329), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_309), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_309), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_321), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_326), .B(n_286), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_326), .B(n_286), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_329), .B(n_294), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_314), .Y(n_371) );
AO21x2_ASAP7_75t_L g372 ( .A1(n_313), .A2(n_305), .B(n_304), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
OAI211xp5_ASAP7_75t_L g374 ( .A1(n_312), .A2(n_277), .B(n_260), .C(n_261), .Y(n_374) );
INVx5_ASAP7_75t_L g375 ( .A(n_329), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_319), .B(n_218), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_320), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g378 ( .A1(n_327), .A2(n_302), .B1(n_308), .B2(n_301), .C1(n_245), .C2(n_153), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_320), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_373), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_350), .B(n_333), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
INVx2_ASAP7_75t_SL g383 ( .A(n_375), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_375), .B(n_333), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_375), .B(n_329), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_336), .Y(n_386) );
AND2x4_ASAP7_75t_SL g387 ( .A(n_346), .B(n_324), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_344), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_350), .B(n_327), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_377), .B(n_310), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_339), .B(n_322), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_344), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_347), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_339), .B(n_312), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_368), .B(n_369), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_368), .B(n_314), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_340), .A2(n_330), .B1(n_280), .B2(n_328), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_344), .Y(n_398) );
AOI221x1_ASAP7_75t_L g399 ( .A1(n_348), .A2(n_332), .B1(n_331), .B2(n_324), .C(n_328), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_347), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_354), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_373), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_369), .B(n_315), .Y(n_403) );
NAND2x1_ASAP7_75t_L g404 ( .A(n_363), .B(n_331), .Y(n_404) );
OAI33xp33_ASAP7_75t_L g405 ( .A1(n_354), .A2(n_138), .A3(n_149), .B1(n_151), .B2(n_139), .B3(n_320), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_375), .B(n_332), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_360), .B(n_310), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_377), .B(n_310), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_378), .B(n_149), .C(n_315), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_379), .B(n_315), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_379), .B(n_317), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_360), .B(n_317), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_352), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_364), .B(n_317), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_364), .B(n_318), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_365), .B(n_318), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_357), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_365), .B(n_318), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_345), .B(n_318), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_358), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_358), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_345), .B(n_328), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_366), .B(n_308), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_351), .B(n_286), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_351), .B(n_300), .Y(n_425) );
NAND4xp25_ASAP7_75t_L g426 ( .A(n_378), .B(n_251), .C(n_153), .D(n_139), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_352), .B(n_286), .Y(n_427) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_371), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_358), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_375), .B(n_287), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_349), .B(n_286), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_371), .B(n_286), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_359), .Y(n_433) );
INVx4_ASAP7_75t_L g434 ( .A(n_375), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_363), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_362), .B(n_300), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_359), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g438 ( .A(n_374), .B(n_153), .C(n_221), .Y(n_438) );
INVx3_ASAP7_75t_SL g439 ( .A(n_375), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_366), .B(n_286), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_367), .B(n_297), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_349), .B(n_300), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_367), .B(n_297), .Y(n_443) );
NAND2x1_ASAP7_75t_L g444 ( .A(n_363), .B(n_297), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_357), .B(n_337), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_342), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_382), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_395), .B(n_353), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_439), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_434), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_381), .B(n_337), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_396), .B(n_353), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_403), .B(n_341), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_387), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_389), .B(n_370), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_382), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_389), .B(n_370), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_386), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_391), .B(n_341), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_435), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_381), .B(n_362), .Y(n_461) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_434), .B(n_342), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_422), .B(n_370), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_409), .B(n_374), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_404), .A2(n_343), .B(n_372), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_386), .B(n_343), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_425), .B(n_359), .Y(n_467) );
OR2x6_ASAP7_75t_L g468 ( .A(n_404), .B(n_342), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_393), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_445), .B(n_338), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_393), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_431), .B(n_370), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_409), .B(n_2), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_387), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_422), .B(n_356), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_419), .B(n_356), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_387), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_431), .B(n_338), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_426), .B(n_4), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_413), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_419), .B(n_356), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_400), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_400), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_439), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_439), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_380), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_407), .B(n_356), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_401), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_401), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_445), .B(n_348), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_407), .B(n_356), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_380), .B(n_372), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_402), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_426), .A2(n_376), .B(n_361), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_390), .B(n_372), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_390), .B(n_372), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_417), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_417), .B(n_355), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_408), .B(n_355), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_394), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_408), .B(n_355), .Y(n_502) );
AOI221xp5_ASAP7_75t_SL g503 ( .A1(n_397), .A2(n_153), .B1(n_156), .B2(n_166), .C(n_7), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_428), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_438), .A2(n_301), .B1(n_355), .B2(n_280), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_414), .B(n_297), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_424), .B(n_4), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_402), .Y(n_508) );
AOI211xp5_ASAP7_75t_L g509 ( .A1(n_383), .A2(n_278), .B(n_6), .C(n_7), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_412), .B(n_5), .Y(n_510) );
AOI221xp5_ASAP7_75t_L g511 ( .A1(n_405), .A2(n_278), .B1(n_128), .B2(n_127), .C(n_225), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_412), .B(n_6), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_414), .B(n_297), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_424), .B(n_9), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_415), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_415), .B(n_287), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_416), .B(n_10), .Y(n_517) );
XNOR2xp5_ASAP7_75t_L g518 ( .A(n_384), .B(n_11), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_427), .B(n_11), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_416), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_427), .B(n_12), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_432), .B(n_14), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_418), .B(n_14), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_418), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_411), .B(n_15), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_411), .B(n_15), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_423), .B(n_16), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_410), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_434), .A2(n_280), .B1(n_276), .B2(n_263), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_464), .A2(n_384), .B1(n_383), .B2(n_423), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_455), .B(n_384), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_450), .B(n_385), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_457), .B(n_384), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_463), .B(n_406), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_447), .Y(n_535) );
INVx2_ASAP7_75t_SL g536 ( .A(n_474), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_494), .A2(n_436), .B1(n_432), .B2(n_440), .C1(n_410), .C2(n_385), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_515), .B(n_406), .Y(n_538) );
AOI222xp33_ASAP7_75t_L g539 ( .A1(n_494), .A2(n_440), .B1(n_385), .B2(n_441), .C1(n_406), .C2(n_446), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_507), .B(n_446), .C(n_444), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_485), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_453), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_496), .B(n_441), .Y(n_543) );
AOI322xp5_ASAP7_75t_L g544 ( .A1(n_497), .A2(n_385), .A3(n_406), .B1(n_444), .B2(n_446), .C1(n_443), .C2(n_430), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_456), .Y(n_545) );
INVxp67_ASAP7_75t_L g546 ( .A(n_480), .Y(n_546) );
OAI33xp33_ASAP7_75t_L g547 ( .A1(n_501), .A2(n_442), .A3(n_443), .B1(n_392), .B2(n_398), .B3(n_420), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g548 ( .A(n_462), .B(n_446), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_527), .A2(n_442), .B1(n_437), .B2(n_433), .C(n_388), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_458), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_469), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_471), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_503), .A2(n_399), .B(n_430), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_450), .Y(n_554) );
AOI222xp33_ASAP7_75t_L g555 ( .A1(n_473), .A2(n_421), .B1(n_433), .B2(n_392), .C1(n_429), .C2(n_388), .Y(n_555) );
OAI31xp33_ASAP7_75t_L g556 ( .A1(n_518), .A2(n_430), .A3(n_433), .B(n_437), .Y(n_556) );
OAI21xp33_ASAP7_75t_SL g557 ( .A1(n_468), .A2(n_437), .B(n_388), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_482), .Y(n_558) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_468), .A2(n_399), .B1(n_430), .B2(n_421), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_448), .B(n_392), .Y(n_560) );
AOI322xp5_ASAP7_75t_L g561 ( .A1(n_461), .A2(n_421), .A3(n_420), .B1(n_398), .B2(n_429), .C1(n_22), .C2(n_23), .Y(n_561) );
OAI221xp5_ASAP7_75t_L g562 ( .A1(n_503), .A2(n_429), .B1(n_420), .B2(n_398), .C(n_280), .Y(n_562) );
AOI322xp5_ASAP7_75t_L g563 ( .A1(n_451), .A2(n_18), .A3(n_19), .B1(n_20), .B2(n_21), .C1(n_23), .C2(n_24), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_452), .B(n_18), .Y(n_564) );
AO22x1_ASAP7_75t_L g565 ( .A1(n_449), .A2(n_276), .B1(n_274), .B2(n_26), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_525), .B(n_24), .Y(n_566) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_449), .B(n_274), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_519), .B(n_269), .C(n_273), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_483), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_484), .A2(n_280), .B1(n_272), .B2(n_276), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_520), .B(n_25), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_524), .B(n_25), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_488), .Y(n_573) );
OAI321xp33_ASAP7_75t_L g574 ( .A1(n_468), .A2(n_505), .A3(n_479), .B1(n_521), .B2(n_522), .C(n_514), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_470), .A2(n_171), .B1(n_176), .B2(n_183), .C(n_190), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_486), .Y(n_576) );
AOI32xp33_ASAP7_75t_L g577 ( .A1(n_484), .A2(n_273), .A3(n_26), .B1(n_265), .B2(n_253), .Y(n_577) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_526), .A2(n_280), .B1(n_214), .B2(n_211), .C(n_263), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_478), .B(n_273), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_470), .B(n_262), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_489), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_510), .B(n_280), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_498), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_500), .B(n_262), .Y(n_584) );
NOR2xp33_ASAP7_75t_SL g585 ( .A(n_495), .B(n_274), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_486), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_459), .Y(n_587) );
OAI311xp33_ASAP7_75t_L g588 ( .A1(n_512), .A2(n_28), .A3(n_29), .B1(n_31), .C1(n_33), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_502), .B(n_262), .Y(n_589) );
OAI22xp33_ASAP7_75t_SL g590 ( .A1(n_495), .A2(n_272), .B1(n_259), .B2(n_263), .Y(n_590) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_472), .A2(n_272), .B1(n_274), .B2(n_246), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_504), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_517), .A2(n_262), .B1(n_272), .B2(n_263), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_528), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_SL g595 ( .A1(n_509), .A2(n_171), .B(n_183), .C(n_210), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_467), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_490), .B(n_262), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_466), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_509), .A2(n_274), .B1(n_259), .B2(n_211), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_490), .B(n_265), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_465), .A2(n_265), .B(n_259), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_460), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_487), .Y(n_603) );
AOI21xp5_ASAP7_75t_SL g604 ( .A1(n_454), .A2(n_274), .B(n_253), .Y(n_604) );
OAI322xp33_ASAP7_75t_L g605 ( .A1(n_492), .A2(n_171), .A3(n_183), .B1(n_187), .B2(n_172), .C1(n_189), .C2(n_204), .Y(n_605) );
OAI31xp33_ASAP7_75t_L g606 ( .A1(n_556), .A2(n_508), .A3(n_493), .B(n_523), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_598), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_L g608 ( .A1(n_544), .A2(n_477), .B(n_476), .C(n_481), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_574), .A2(n_499), .B1(n_508), .B2(n_493), .C(n_475), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_576), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_592), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_595), .A2(n_499), .B(n_491), .C(n_511), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_537), .B(n_516), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_535), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_545), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_536), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_550), .Y(n_617) );
XNOR2xp5_ASAP7_75t_L g618 ( .A(n_603), .B(n_529), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_543), .B(n_513), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_562), .A2(n_506), .B1(n_513), .B2(n_253), .Y(n_620) );
OA211x2_ASAP7_75t_L g621 ( .A1(n_553), .A2(n_506), .B(n_35), .C(n_37), .Y(n_621) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_557), .A2(n_253), .B(n_222), .C(n_206), .Y(n_622) );
AOI32xp33_ASAP7_75t_L g623 ( .A1(n_574), .A2(n_222), .A3(n_210), .B1(n_206), .B2(n_40), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_SL g624 ( .A1(n_566), .A2(n_222), .B(n_210), .C(n_206), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_551), .Y(n_625) );
CKINVDCx16_ASAP7_75t_R g626 ( .A(n_564), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_586), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_531), .B(n_34), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_560), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_552), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_587), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_558), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_549), .A2(n_204), .B1(n_215), .B2(n_209), .C1(n_203), .C2(n_187), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_577), .A2(n_222), .B(n_210), .C(n_215), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_599), .A2(n_209), .B1(n_203), .B2(n_189), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_569), .Y(n_636) );
OAI22xp33_ASAP7_75t_SL g637 ( .A1(n_554), .A2(n_38), .B1(n_39), .B2(n_42), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_540), .B(n_45), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_539), .B(n_189), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_573), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_581), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_542), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_537), .B(n_46), .Y(n_643) );
AO22x2_ASAP7_75t_L g644 ( .A1(n_602), .A2(n_47), .B1(n_48), .B2(n_52), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_583), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_534), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_594), .Y(n_647) );
OAI211xp5_ASAP7_75t_SL g648 ( .A1(n_539), .A2(n_53), .B(n_54), .C(n_55), .Y(n_648) );
XOR2x2_ASAP7_75t_L g649 ( .A(n_578), .B(n_58), .Y(n_649) );
OAI21xp33_ASAP7_75t_L g650 ( .A1(n_553), .A2(n_189), .B(n_172), .Y(n_650) );
INVx6_ASAP7_75t_L g651 ( .A(n_571), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_555), .B(n_61), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_559), .A2(n_189), .B(n_172), .C(n_187), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_533), .B(n_65), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_596), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g656 ( .A1(n_606), .A2(n_530), .B1(n_546), .B2(n_555), .C(n_548), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_614), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_609), .B(n_561), .C(n_563), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_608), .A2(n_548), .B1(n_532), .B2(n_593), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_623), .A2(n_572), .B(n_570), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_613), .A2(n_547), .B1(n_582), .B2(n_589), .C(n_584), .Y(n_661) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_648), .B(n_604), .Y(n_662) );
OA22x2_ASAP7_75t_L g663 ( .A1(n_616), .A2(n_541), .B1(n_538), .B2(n_601), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g664 ( .A1(n_620), .A2(n_588), .B(n_590), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_607), .A2(n_580), .B1(n_565), .B2(n_601), .C(n_597), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_653), .B(n_585), .Y(n_666) );
BUFx2_ASAP7_75t_SL g667 ( .A(n_627), .Y(n_667) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_639), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_642), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_610), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_650), .A2(n_567), .B(n_585), .C(n_579), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g672 ( .A1(n_643), .A2(n_600), .B(n_591), .Y(n_672) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_638), .B(n_605), .Y(n_673) );
INVx2_ASAP7_75t_SL g674 ( .A(n_651), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g675 ( .A1(n_650), .A2(n_568), .B1(n_575), .B2(n_68), .C(n_70), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_621), .A2(n_189), .B1(n_172), .B2(n_187), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_626), .A2(n_172), .B1(n_187), .B2(n_71), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_637), .A2(n_172), .B(n_187), .Y(n_678) );
XNOR2x1_ASAP7_75t_L g679 ( .A(n_618), .B(n_66), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_615), .Y(n_680) );
OA22x2_ASAP7_75t_L g681 ( .A1(n_646), .A2(n_67), .B1(n_72), .B2(n_73), .Y(n_681) );
AOI211xp5_ASAP7_75t_L g682 ( .A1(n_637), .A2(n_187), .B(n_75), .C(n_76), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_655), .B(n_74), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_669), .Y(n_684) );
O2A1O1Ixp33_ASAP7_75t_L g685 ( .A1(n_668), .A2(n_624), .B(n_652), .C(n_634), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_656), .A2(n_621), .B1(n_651), .B2(n_649), .Y(n_686) );
XNOR2x1_ASAP7_75t_L g687 ( .A(n_679), .B(n_644), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_661), .B(n_647), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_657), .B(n_632), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_659), .A2(n_612), .B1(n_611), .B2(n_635), .C(n_640), .Y(n_690) );
INVx1_ASAP7_75t_SL g691 ( .A(n_667), .Y(n_691) );
NAND4xp25_ASAP7_75t_L g692 ( .A(n_664), .B(n_633), .C(n_635), .D(n_638), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_658), .B(n_628), .C(n_654), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_665), .A2(n_645), .B1(n_617), .B2(n_641), .C(n_636), .Y(n_694) );
OAI221xp5_ASAP7_75t_SL g695 ( .A1(n_660), .A2(n_619), .B1(n_622), .B2(n_631), .C(n_625), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_672), .A2(n_630), .B1(n_629), .B2(n_644), .C(n_82), .Y(n_696) );
OAI221xp5_ASAP7_75t_SL g697 ( .A1(n_674), .A2(n_77), .B1(n_78), .B2(n_80), .C(n_83), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_691), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_690), .A2(n_666), .B(n_675), .C(n_671), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_687), .B(n_695), .Y(n_700) );
NOR2xp33_ASAP7_75t_R g701 ( .A(n_686), .B(n_683), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_692), .B(n_673), .C(n_662), .Y(n_702) );
NOR2xp67_ASAP7_75t_L g703 ( .A(n_684), .B(n_670), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_688), .A2(n_663), .B(n_682), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_702), .A2(n_693), .B1(n_696), .B2(n_694), .Y(n_705) );
OR3x1_ASAP7_75t_L g706 ( .A(n_700), .B(n_685), .C(n_680), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_704), .A2(n_682), .B(n_681), .Y(n_707) );
OR4x2_ASAP7_75t_L g708 ( .A(n_701), .B(n_699), .C(n_698), .D(n_703), .Y(n_708) );
XNOR2x1_ASAP7_75t_L g709 ( .A(n_707), .B(n_677), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_705), .B(n_689), .Y(n_710) );
INVx2_ASAP7_75t_SL g711 ( .A(n_708), .Y(n_711) );
OAI22xp5_ASAP7_75t_SL g712 ( .A1(n_711), .A2(n_706), .B1(n_707), .B2(n_677), .Y(n_712) );
XNOR2xp5_ASAP7_75t_L g713 ( .A(n_709), .B(n_683), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_712), .A2(n_710), .B1(n_689), .B2(n_676), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_713), .A2(n_678), .B1(n_697), .B2(n_199), .Y(n_715) );
AOI222xp33_ASAP7_75t_SL g716 ( .A1(n_714), .A2(n_86), .B1(n_87), .B2(n_88), .C1(n_89), .C2(n_93), .Y(n_716) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_715), .A2(n_96), .B(n_98), .Y(n_717) );
OAI221xp5_ASAP7_75t_R g718 ( .A1(n_716), .A2(n_99), .B1(n_100), .B2(n_102), .C(n_104), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_717), .B(n_105), .Y(n_719) );
endmodule