module real_aes_6295_n_239 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_239);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_239;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_763;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_725;
wire n_504;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_751;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_741;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_639;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp5_ASAP7_75t_SL g527 ( .A1(n_0), .A2(n_206), .B1(n_528), .B2(n_529), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_1), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_2), .A2(n_200), .B1(n_280), .B2(n_283), .Y(n_279) );
AOI222xp33_ASAP7_75t_L g559 ( .A1(n_3), .A2(n_78), .B1(n_222), .B2(n_324), .C1(n_331), .C2(n_445), .Y(n_559) );
INVx1_ASAP7_75t_L g622 ( .A(n_4), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_5), .A2(n_17), .B1(n_651), .B2(n_652), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_6), .B(n_480), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_7), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_8), .A2(n_111), .B1(n_466), .B2(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g619 ( .A(n_9), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_10), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_11), .A2(n_113), .B1(n_421), .B2(n_456), .Y(n_473) );
AOI222xp33_ASAP7_75t_L g507 ( .A1(n_12), .A2(n_110), .B1(n_188), .B2(n_327), .C1(n_451), .C2(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_13), .A2(n_47), .B1(n_651), .B2(n_659), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_14), .A2(n_721), .B1(n_747), .B2(n_748), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_14), .Y(n_747) );
AOI22xp33_ASAP7_75t_SL g407 ( .A1(n_15), .A2(n_51), .B1(n_408), .B2(n_410), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_16), .A2(n_123), .B1(n_308), .B2(n_311), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_18), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_19), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_20), .A2(n_79), .B1(n_125), .B2(n_380), .C1(n_669), .C2(n_670), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_21), .B(n_311), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_22), .A2(n_109), .B1(n_297), .B2(n_363), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_23), .Y(n_597) );
AO22x2_ASAP7_75t_L g260 ( .A1(n_24), .A2(n_80), .B1(n_261), .B2(n_262), .Y(n_260) );
INVx1_ASAP7_75t_L g717 ( .A(n_24), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_25), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_26), .A2(n_176), .B1(n_456), .B2(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_27), .A2(n_129), .B1(n_291), .B2(n_486), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_28), .A2(n_184), .B1(n_445), .B2(n_446), .Y(n_537) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_29), .A2(n_121), .B1(n_465), .B2(n_529), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_30), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_31), .A2(n_238), .B1(n_458), .B2(n_460), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_32), .A2(n_141), .B1(n_347), .B2(n_417), .Y(n_693) );
INVx1_ASAP7_75t_L g725 ( .A(n_33), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_34), .Y(n_727) );
AOI222xp33_ASAP7_75t_L g323 ( .A1(n_35), .A2(n_173), .B1(n_218), .B2(n_324), .C1(n_327), .C2(n_331), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_36), .A2(n_214), .B1(n_360), .B2(n_465), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_37), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_38), .B(n_308), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_39), .A2(n_168), .B1(n_405), .B2(n_406), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_40), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_41), .Y(n_381) );
AO22x2_ASAP7_75t_L g264 ( .A1(n_42), .A2(n_83), .B1(n_261), .B2(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g718 ( .A(n_42), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_43), .A2(n_118), .B1(n_320), .B2(n_332), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_44), .A2(n_128), .B1(n_350), .B2(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g569 ( .A(n_45), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_46), .A2(n_142), .B1(n_417), .B2(n_420), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_48), .A2(n_77), .B1(n_658), .B2(n_659), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_49), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_50), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_52), .A2(n_55), .B1(n_415), .B2(n_416), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_53), .Y(n_358) );
AOI222xp33_ASAP7_75t_L g487 ( .A1(n_54), .A2(n_166), .B1(n_223), .B2(n_324), .C1(n_445), .C2(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_56), .A2(n_64), .B1(n_465), .B2(n_466), .Y(n_464) );
AOI22xp5_ASAP7_75t_SL g525 ( .A1(n_57), .A2(n_137), .B1(n_289), .B2(n_347), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_58), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_59), .A2(n_195), .B1(n_293), .B2(n_343), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_60), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_61), .A2(n_233), .B1(n_280), .B2(n_495), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_62), .A2(n_131), .B1(n_319), .B2(n_446), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_63), .A2(n_160), .B1(n_420), .B2(n_458), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_65), .A2(n_172), .B1(n_314), .B2(n_376), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_66), .Y(n_633) );
AOI22xp5_ASAP7_75t_SL g523 ( .A1(n_67), .A2(n_124), .B1(n_475), .B2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_68), .A2(n_194), .B1(n_312), .B2(n_409), .Y(n_538) );
XNOR2x2_ASAP7_75t_L g541 ( .A(n_69), .B(n_542), .Y(n_541) );
AO22x2_ASAP7_75t_L g673 ( .A1(n_70), .A2(n_674), .B1(n_698), .B2(n_699), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_70), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_71), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_72), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_73), .A2(n_96), .B1(n_419), .B2(n_421), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_74), .A2(n_203), .B1(n_486), .B2(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_75), .A2(n_199), .B1(n_408), .B2(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_SL g625 ( .A1(n_76), .A2(n_130), .B1(n_417), .B2(n_524), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_81), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_82), .A2(n_231), .B1(n_289), .B2(n_291), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_84), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_85), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_86), .Y(n_490) );
INVx1_ASAP7_75t_L g247 ( .A(n_87), .Y(n_247) );
INVx1_ASAP7_75t_L g758 ( .A(n_88), .Y(n_758) );
AOI22xp5_ASAP7_75t_SL g762 ( .A1(n_88), .A2(n_721), .B1(n_748), .B2(n_758), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_89), .A2(n_226), .B1(n_297), .B2(n_302), .Y(n_296) );
INVx1_ASAP7_75t_L g467 ( .A(n_90), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_91), .A2(n_114), .B1(n_351), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_92), .A2(n_122), .B1(n_661), .B2(n_663), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_93), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_94), .A2(n_163), .B1(n_319), .B2(n_331), .Y(n_639) );
INVx1_ASAP7_75t_L g243 ( .A(n_95), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_97), .Y(n_432) );
XOR2x2_ASAP7_75t_L g250 ( .A(n_98), .B(n_251), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_99), .A2(n_165), .B1(n_550), .B2(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g596 ( .A(n_100), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_101), .A2(n_136), .B1(n_406), .B2(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_102), .A2(n_212), .B1(n_421), .B2(n_502), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g422 ( .A1(n_103), .A2(n_423), .B(n_424), .C(n_431), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_104), .A2(n_190), .B1(n_445), .B2(n_446), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_105), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_106), .A2(n_149), .B1(n_294), .B2(n_495), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_107), .B(n_308), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_108), .A2(n_155), .B1(n_455), .B2(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g449 ( .A(n_112), .Y(n_449) );
INVx1_ASAP7_75t_L g620 ( .A(n_115), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_116), .A2(n_204), .B1(n_303), .B2(n_463), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_117), .A2(n_207), .B1(n_314), .B2(n_319), .Y(n_313) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_119), .A2(n_232), .B1(n_496), .B2(n_548), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_120), .A2(n_159), .B1(n_320), .B2(n_451), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_126), .Y(n_509) );
AND2x2_ASAP7_75t_L g246 ( .A(n_127), .B(n_247), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_132), .Y(n_396) );
INVx1_ASAP7_75t_L g577 ( .A(n_133), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_134), .A2(n_202), .B1(n_320), .B2(n_405), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_135), .A2(n_182), .B1(n_314), .B2(n_558), .Y(n_557) );
AND2x6_ASAP7_75t_L g242 ( .A(n_138), .B(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_138), .Y(n_711) );
AO22x2_ASAP7_75t_L g268 ( .A1(n_139), .A2(n_201), .B1(n_261), .B2(n_265), .Y(n_268) );
INVx1_ASAP7_75t_L g579 ( .A(n_140), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_143), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_144), .A2(n_220), .B1(n_495), .B2(n_496), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_145), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_146), .A2(n_180), .B1(n_475), .B2(n_476), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_147), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_148), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_150), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_151), .Y(n_504) );
OA22x2_ASAP7_75t_L g563 ( .A1(n_152), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_152), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_153), .A2(n_236), .B1(n_280), .B2(n_551), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_154), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_156), .A2(n_339), .B1(n_387), .B2(n_388), .Y(n_338) );
INVx1_ASAP7_75t_L g387 ( .A(n_156), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_157), .A2(n_177), .B1(n_415), .B2(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_158), .A2(n_164), .B1(n_398), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_161), .A2(n_187), .B1(n_738), .B2(n_739), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_162), .A2(n_224), .B1(n_421), .B2(n_455), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_167), .A2(n_191), .B1(n_319), .B2(n_331), .Y(n_575) );
AO22x2_ASAP7_75t_L g270 ( .A1(n_169), .A2(n_216), .B1(n_261), .B2(n_262), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_170), .A2(n_230), .B1(n_406), .B2(n_451), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_171), .A2(n_193), .B1(n_283), .B2(n_423), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_174), .A2(n_192), .B1(n_548), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_175), .A2(n_219), .B1(n_488), .B2(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g593 ( .A(n_178), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_179), .A2(n_185), .B1(n_429), .B2(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g724 ( .A(n_181), .Y(n_724) );
INVx1_ASAP7_75t_L g616 ( .A(n_183), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_186), .B(n_529), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_189), .A2(n_217), .B1(n_303), .B2(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_196), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_197), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g239 ( .A1(n_198), .A2(n_240), .B(n_248), .C(n_719), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_201), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g573 ( .A(n_205), .Y(n_573) );
AOI22xp5_ASAP7_75t_SL g628 ( .A1(n_208), .A2(n_237), .B1(n_434), .B2(n_460), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_209), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_210), .A2(n_221), .B1(n_412), .B2(n_480), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_211), .Y(n_679) );
INVx1_ASAP7_75t_L g571 ( .A(n_213), .Y(n_571) );
XNOR2xp5_ASAP7_75t_L g391 ( .A(n_215), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g714 ( .A(n_216), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_225), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_227), .A2(n_229), .B1(n_254), .B2(n_271), .Y(n_253) );
INVx1_ASAP7_75t_L g261 ( .A(n_228), .Y(n_261) );
INVx1_ASAP7_75t_L g263 ( .A(n_228), .Y(n_263) );
OA22x2_ASAP7_75t_L g646 ( .A1(n_234), .A2(n_647), .B1(n_648), .B2(n_671), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_234), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_235), .Y(n_402) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_243), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_244), .A2(n_709), .B(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_245), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_515), .B1(n_704), .B2(n_705), .C(n_706), .Y(n_248) );
INVx1_ASAP7_75t_L g704 ( .A(n_249), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_334), .B1(n_513), .B2(n_514), .Y(n_249) );
INVx1_ASAP7_75t_L g513 ( .A(n_250), .Y(n_513) );
NAND4xp75_ASAP7_75t_L g251 ( .A(n_252), .B(n_287), .C(n_306), .D(n_323), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_279), .Y(n_252) );
INVx4_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx4_ASAP7_75t_L g434 ( .A(n_255), .Y(n_434) );
INVx3_ASAP7_75t_L g475 ( .A(n_255), .Y(n_475) );
INVx2_ASAP7_75t_SL g659 ( .A(n_255), .Y(n_659) );
INVx11_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx11_ASAP7_75t_L g344 ( .A(n_256), .Y(n_344) );
AND2x6_ASAP7_75t_L g256 ( .A(n_257), .B(n_266), .Y(n_256) );
AND2x4_ASAP7_75t_L g310 ( .A(n_257), .B(n_282), .Y(n_310) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g368 ( .A(n_258), .B(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_264), .Y(n_258) );
AND2x2_ASAP7_75t_L g277 ( .A(n_259), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g295 ( .A(n_259), .B(n_264), .Y(n_295) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g318 ( .A(n_260), .B(n_268), .Y(n_318) );
AND2x2_ASAP7_75t_L g322 ( .A(n_260), .B(n_264), .Y(n_322) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g265 ( .A(n_263), .Y(n_265) );
INVx2_ASAP7_75t_L g278 ( .A(n_264), .Y(n_278) );
INVx1_ASAP7_75t_L g305 ( .A(n_264), .Y(n_305) );
AND2x2_ASAP7_75t_L g290 ( .A(n_266), .B(n_277), .Y(n_290) );
AND2x4_ASAP7_75t_L g294 ( .A(n_266), .B(n_295), .Y(n_294) );
AND2x6_ASAP7_75t_L g326 ( .A(n_266), .B(n_322), .Y(n_326) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
AND2x2_ASAP7_75t_L g282 ( .A(n_267), .B(n_270), .Y(n_282) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g275 ( .A(n_268), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_268), .B(n_270), .Y(n_286) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g276 ( .A(n_270), .Y(n_276) );
INVx1_ASAP7_75t_L g330 ( .A(n_270), .Y(n_330) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx3_ASAP7_75t_L g354 ( .A(n_274), .Y(n_354) );
BUFx3_ASAP7_75t_L g417 ( .A(n_274), .Y(n_417) );
BUFx3_ASAP7_75t_L g456 ( .A(n_274), .Y(n_456) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
AND2x2_ASAP7_75t_L g301 ( .A(n_275), .B(n_295), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_275), .B(n_295), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_275), .B(n_277), .Y(n_617) );
INVx1_ASAP7_75t_L g321 ( .A(n_276), .Y(n_321) );
AND2x4_ASAP7_75t_L g281 ( .A(n_277), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g284 ( .A(n_277), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g329 ( .A(n_278), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g530 ( .A(n_278), .Y(n_530) );
BUFx2_ASAP7_75t_L g357 ( .A(n_280), .Y(n_357) );
BUFx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx3_ASAP7_75t_L g420 ( .A(n_281), .Y(n_420) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_281), .Y(n_465) );
BUFx3_ASAP7_75t_L g502 ( .A(n_281), .Y(n_502) );
INVx2_ASAP7_75t_L g604 ( .A(n_281), .Y(n_604) );
AND2x6_ASAP7_75t_L g312 ( .A(n_282), .B(n_295), .Y(n_312) );
INVx1_ASAP7_75t_L g369 ( .A(n_282), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g373 ( .A(n_282), .B(n_295), .Y(n_373) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_SL g360 ( .A(n_284), .Y(n_360) );
BUFx3_ASAP7_75t_L g421 ( .A(n_284), .Y(n_421) );
BUFx3_ASAP7_75t_L g460 ( .A(n_284), .Y(n_460) );
BUFx3_ASAP7_75t_L g528 ( .A(n_284), .Y(n_528) );
INVx1_ASAP7_75t_L g613 ( .A(n_284), .Y(n_613) );
BUFx2_ASAP7_75t_L g663 ( .A(n_284), .Y(n_663) );
BUFx2_ASAP7_75t_SL g739 ( .A(n_284), .Y(n_739) );
AND2x2_ASAP7_75t_L g529 ( .A(n_285), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x6_ASAP7_75t_L g304 ( .A(n_286), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_296), .Y(n_287) );
BUFx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_290), .Y(n_351) );
BUFx2_ASAP7_75t_SL g423 ( .A(n_290), .Y(n_423) );
INVx2_ASAP7_75t_L g459 ( .A(n_290), .Y(n_459) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx3_ASAP7_75t_L g347 ( .A(n_294), .Y(n_347) );
BUFx3_ASAP7_75t_L g415 ( .A(n_294), .Y(n_415) );
INVx6_ASAP7_75t_L g477 ( .A(n_294), .Y(n_477) );
INVx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx2_ASAP7_75t_L g655 ( .A(n_299), .Y(n_655) );
INVx4_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx5_ASAP7_75t_L g463 ( .A(n_300), .Y(n_463) );
INVx2_ASAP7_75t_L g486 ( .A(n_300), .Y(n_486) );
INVx3_ASAP7_75t_L g524 ( .A(n_300), .Y(n_524) );
INVx1_ASAP7_75t_L g550 ( .A(n_300), .Y(n_550) );
BUFx3_ASAP7_75t_L g742 ( .A(n_300), .Y(n_742) );
INVx8_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx2_ASAP7_75t_L g429 ( .A(n_303), .Y(n_429) );
BUFx2_ASAP7_75t_L g695 ( .A(n_303), .Y(n_695) );
INVx6_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g363 ( .A(n_304), .Y(n_363) );
INVx1_ASAP7_75t_SL g466 ( .A(n_304), .Y(n_466) );
INVx1_ASAP7_75t_L g551 ( .A(n_304), .Y(n_551) );
INVx1_ASAP7_75t_L g317 ( .A(n_305), .Y(n_317) );
AND2x2_ASAP7_75t_SL g306 ( .A(n_307), .B(n_313), .Y(n_306) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx5_ASAP7_75t_L g409 ( .A(n_309), .Y(n_409) );
INVx2_ASAP7_75t_L g480 ( .A(n_309), .Y(n_480) );
INVx4_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx4f_ASAP7_75t_L g412 ( .A(n_312), .Y(n_412) );
BUFx2_ASAP7_75t_L g666 ( .A(n_312), .Y(n_666) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g405 ( .A(n_316), .Y(n_405) );
BUFx3_ASAP7_75t_L g446 ( .A(n_316), .Y(n_446) );
BUFx2_ASAP7_75t_L g482 ( .A(n_316), .Y(n_482) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x4_ASAP7_75t_L g328 ( .A(n_318), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g332 ( .A(n_318), .B(n_333), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_318), .B(n_530), .Y(n_580) );
INVx1_ASAP7_75t_SL g377 ( .A(n_319), .Y(n_377) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx3_ASAP7_75t_L g406 ( .A(n_320), .Y(n_406) );
BUFx2_ASAP7_75t_SL g558 ( .A(n_320), .Y(n_558) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g691 ( .A(n_321), .Y(n_691) );
INVx1_ASAP7_75t_L g690 ( .A(n_322), .Y(n_690) );
INVx4_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI22xp5_ASAP7_75t_SL g640 ( .A1(n_325), .A2(n_641), .B1(n_642), .B2(n_643), .Y(n_640) );
INVx4_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_SL g382 ( .A(n_326), .Y(n_382) );
INVx2_ASAP7_75t_L g395 ( .A(n_326), .Y(n_395) );
INVx2_ASAP7_75t_L g448 ( .A(n_326), .Y(n_448) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_326), .Y(n_508) );
BUFx3_ASAP7_75t_L g669 ( .A(n_326), .Y(n_669) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx4f_ASAP7_75t_SL g380 ( .A(n_328), .Y(n_380) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_328), .Y(n_399) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_328), .Y(n_445) );
BUFx2_ASAP7_75t_L g684 ( .A(n_328), .Y(n_684) );
INVx1_ASAP7_75t_L g333 ( .A(n_330), .Y(n_333) );
INVx1_ASAP7_75t_L g401 ( .A(n_331), .Y(n_401) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_332), .Y(n_385) );
BUFx12f_ASAP7_75t_L g451 ( .A(n_332), .Y(n_451) );
INVx1_ASAP7_75t_L g514 ( .A(n_334), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_435), .B2(n_512), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI22xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_338), .B1(n_389), .B2(n_390), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g388 ( .A(n_339), .Y(n_388) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_364), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_355), .Y(n_340) );
OAI221xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_345), .B1(n_346), .B2(n_348), .C(n_349), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_SL g455 ( .A(n_344), .Y(n_455) );
INVx5_ASAP7_75t_SL g496 ( .A(n_344), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_344), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g658 ( .A(n_351), .Y(n_658) );
INVx3_ASAP7_75t_L g746 ( .A(n_351), .Y(n_746) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx4f_ASAP7_75t_SL g548 ( .A(n_354), .Y(n_548) );
OAI221xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_358), .B1(n_359), .B2(n_361), .C(n_362), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_378), .Y(n_364) );
OAI221xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_370), .B1(n_371), .B2(n_374), .C(n_375), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_366), .A2(n_372), .B1(n_724), .B2(n_725), .Y(n_723) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g678 ( .A(n_367), .Y(n_678) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_368), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_368), .A2(n_593), .B(n_594), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_371), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OA211x2_ASAP7_75t_L g503 ( .A1(n_372), .A2(n_504), .B(n_505), .C(n_506), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_372), .A2(n_580), .B1(n_596), .B2(n_597), .Y(n_595) );
BUFx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g555 ( .A(n_373), .Y(n_555) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI222xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B1(n_382), .B2(n_383), .C1(n_384), .C2(n_386), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_382), .A2(n_599), .B1(n_600), .B2(n_601), .Y(n_598) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g729 ( .A(n_385), .Y(n_729) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND3x1_ASAP7_75t_L g392 ( .A(n_393), .B(n_413), .C(n_422), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_403), .Y(n_393) );
OAI222xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_397), .B2(n_400), .C1(n_401), .C2(n_402), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_395), .A2(n_534), .B(n_535), .Y(n_533) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g578 ( .A(n_399), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_418), .Y(n_413) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g653 ( .A(n_417), .Y(n_653) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_427), .B1(n_428), .B2(n_430), .Y(n_424) );
BUFx2_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_426), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g512 ( .A(n_435), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_437), .B1(n_468), .B2(n_469), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
XOR2x2_ASAP7_75t_SL g438 ( .A(n_439), .B(n_467), .Y(n_438) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_440), .B(n_452), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_447), .Y(n_440) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .C(n_444), .Y(n_441) );
INVx4_ASAP7_75t_L g601 ( .A(n_445), .Y(n_601) );
INVx2_ASAP7_75t_L g642 ( .A(n_445), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_449), .B(n_450), .Y(n_447) );
INVx2_ASAP7_75t_L g489 ( .A(n_451), .Y(n_489) );
BUFx4f_ASAP7_75t_SL g670 ( .A(n_451), .Y(n_670) );
NOR2x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_461), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_457), .Y(n_453) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g607 ( .A1(n_459), .A2(n_477), .B1(n_608), .B2(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx4_ASAP7_75t_L g662 ( .A(n_465), .Y(n_662) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AO22x1_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_491), .B1(n_510), .B2(n_511), .Y(n_469) );
INVx2_ASAP7_75t_SL g510 ( .A(n_470), .Y(n_510) );
XOR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_490), .Y(n_470) );
NAND4xp75_ASAP7_75t_L g471 ( .A(n_472), .B(n_478), .C(n_483), .D(n_487), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx3_ASAP7_75t_L g500 ( .A(n_477), .Y(n_500) );
INVx2_ASAP7_75t_L g651 ( .A(n_477), .Y(n_651) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_479), .B(n_481), .Y(n_478) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g511 ( .A(n_491), .Y(n_511) );
XOR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_509), .Y(n_491) );
NAND4xp75_ASAP7_75t_L g492 ( .A(n_493), .B(n_498), .C(n_503), .D(n_507), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .Y(n_493) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
INVx2_ASAP7_75t_SL g574 ( .A(n_508), .Y(n_574) );
INVx1_ASAP7_75t_L g705 ( .A(n_515), .Y(n_705) );
AOI22xp5_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_645), .B1(n_702), .B2(n_703), .Y(n_515) );
INVx1_ASAP7_75t_L g702 ( .A(n_516), .Y(n_702) );
XOR2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_560), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B1(n_540), .B2(n_541), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
XOR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_539), .Y(n_521) );
NAND4xp75_ASAP7_75t_SL g522 ( .A(n_523), .B(n_525), .C(n_526), .D(n_532), .Y(n_522) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_531), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_536), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND4xp75_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .C(n_552), .D(n_559), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
OA211x2_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B(n_556), .C(n_557), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g632 ( .A(n_555), .Y(n_632) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AO22x2_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_588), .B2(n_644), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_581), .Y(n_566) );
NOR3xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .C(n_576), .Y(n_567) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_570), .A2(n_638), .B(n_639), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B(n_575), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_576) );
INVx4_ASAP7_75t_L g635 ( .A(n_580), .Y(n_635) );
BUFx3_ASAP7_75t_L g732 ( .A(n_580), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx2_ASAP7_75t_L g644 ( .A(n_588), .Y(n_644) );
XOR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_621), .Y(n_588) );
XNOR2x1_ASAP7_75t_L g589 ( .A(n_590), .B(n_620), .Y(n_589) );
AND3x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_602), .C(n_610), .Y(n_590) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .C(n_598), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_607), .Y(n_602) );
OAI21xp5_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B(n_606), .Y(n_603) );
INVx2_ASAP7_75t_L g738 ( .A(n_604), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_615), .C(n_618), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
XNOR2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND3x1_ASAP7_75t_SL g623 ( .A(n_624), .B(n_627), .C(n_630), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NOR3xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_637), .C(n_640), .Y(n_630) );
OAI22xp5_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_633), .B1(n_634), .B2(n_636), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_632), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_676) );
INVx3_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g687 ( .A(n_635), .Y(n_687) );
INVx1_ASAP7_75t_L g703 ( .A(n_645), .Y(n_703) );
AOI22x1_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_672), .B1(n_700), .B2(n_701), .Y(n_645) );
INVx1_ASAP7_75t_L g700 ( .A(n_646), .Y(n_700) );
INVx1_ASAP7_75t_SL g671 ( .A(n_648), .Y(n_671) );
NAND4xp75_ASAP7_75t_L g648 ( .A(n_649), .B(n_656), .C(n_664), .D(n_668), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_654), .Y(n_649) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_660), .Y(n_656) );
INVx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_SL g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx3_ASAP7_75t_L g682 ( .A(n_669), .Y(n_682) );
INVx1_ASAP7_75t_L g701 ( .A(n_672), .Y(n_701) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g698 ( .A(n_674), .Y(n_698) );
AND2x2_ASAP7_75t_SL g674 ( .A(n_675), .B(n_692), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_680), .C(n_685), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B(n_683), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g726 ( .A1(n_682), .A2(n_727), .B(n_728), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_685) );
CKINVDCx16_ASAP7_75t_R g735 ( .A(n_689), .Y(n_735) );
OR2x6_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
AND4x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .C(n_696), .D(n_697), .Y(n_692) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_712), .Y(n_707) );
OR2x2_ASAP7_75t_SL g765 ( .A(n_708), .B(n_713), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_709), .Y(n_750) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_710), .B(n_754), .Y(n_757) );
CKINVDCx16_ASAP7_75t_R g754 ( .A(n_711), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
OAI322xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_749), .A3(n_751), .B1(n_755), .B2(n_758), .C1(n_759), .C2(n_763), .Y(n_719) );
INVx2_ASAP7_75t_SL g748 ( .A(n_721), .Y(n_748) );
AND2x2_ASAP7_75t_SL g721 ( .A(n_722), .B(n_736), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_726), .C(n_730), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_730) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND4x1_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .C(n_743), .D(n_744), .Y(n_736) );
INVx3_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
BUFx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
CKINVDCx16_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
endmodule