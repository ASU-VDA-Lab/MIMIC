module fake_jpeg_17809_n_384 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_384);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_384;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_6),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_39),
.B(n_56),
.Y(n_89)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_31),
.B1(n_35),
.B2(n_26),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_5),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_5),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_14),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_14),
.B(n_32),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_69),
.Y(n_80)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_55),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_83),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_86),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_22),
.B1(n_34),
.B2(n_20),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_75),
.A2(n_104),
.B1(n_105),
.B2(n_21),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_14),
.B1(n_35),
.B2(n_26),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_76),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_36),
.C(n_15),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_77),
.B(n_36),
.C(n_46),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_57),
.B1(n_59),
.B2(n_42),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_38),
.B(n_19),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_108),
.Y(n_161)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_40),
.A2(n_34),
.B1(n_20),
.B2(n_30),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_34),
.B1(n_30),
.B2(n_17),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_39),
.B(n_29),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_29),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_116),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_40),
.A2(n_17),
.B1(n_35),
.B2(n_32),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_21),
.B1(n_45),
.B2(n_63),
.Y(n_148)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_61),
.B(n_25),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_25),
.Y(n_117)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_123),
.A2(n_148),
.B1(n_82),
.B2(n_85),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_70),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_125),
.A2(n_126),
.B1(n_135),
.B2(n_106),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_89),
.B(n_21),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_128),
.B(n_157),
.Y(n_195)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_131),
.A2(n_135),
.B(n_125),
.Y(n_179)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_31),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_142),
.B(n_4),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_143),
.B(n_172),
.Y(n_186)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_76),
.A2(n_57),
.B1(n_59),
.B2(n_42),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_99),
.B1(n_113),
.B2(n_118),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_156),
.Y(n_178)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_104),
.B(n_45),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_88),
.A2(n_48),
.B1(n_64),
.B2(n_49),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_114),
.B1(n_79),
.B2(n_85),
.Y(n_181)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_171),
.Y(n_215)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_163),
.Y(n_196)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_168),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_96),
.B(n_51),
.C(n_44),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_69),
.C(n_53),
.Y(n_176)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_170),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_92),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_10),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_174),
.B(n_192),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_175),
.A2(n_184),
.B1(n_193),
.B2(n_202),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_165),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_156),
.B(n_113),
.C(n_118),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_177),
.A2(n_188),
.B(n_207),
.C(n_197),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_SL g218 ( 
.A1(n_179),
.A2(n_181),
.B(n_191),
.C(n_124),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_182),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_140),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_82),
.B(n_72),
.C(n_114),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_125),
.A2(n_79),
.B1(n_36),
.B2(n_53),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_126),
.A2(n_10),
.B(n_13),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_126),
.A2(n_43),
.B1(n_74),
.B2(n_86),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_43),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_208),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_143),
.A2(n_62),
.B1(n_8),
.B2(n_9),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_211),
.B1(n_8),
.B2(n_12),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_166),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_205),
.B(n_201),
.Y(n_253)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_127),
.B(n_0),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_210),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_142),
.A2(n_8),
.B1(n_10),
.B2(n_9),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_3),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_191),
.C(n_196),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

AO22x1_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_159),
.B1(n_144),
.B2(n_138),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_249),
.B(n_224),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_218),
.A2(n_223),
.B(n_253),
.Y(n_273)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_137),
.C(n_150),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_222),
.C(n_230),
.Y(n_259)
);

AO22x1_ASAP7_75t_SL g224 ( 
.A1(n_177),
.A2(n_141),
.B1(n_147),
.B2(n_140),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_224),
.A2(n_181),
.B1(n_177),
.B2(n_165),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_137),
.B1(n_153),
.B2(n_154),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_232),
.B1(n_234),
.B2(n_237),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_167),
.C(n_139),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_227),
.A2(n_231),
.B1(n_238),
.B2(n_254),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_170),
.B(n_134),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_229),
.B(n_250),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_10),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_173),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_136),
.B1(n_163),
.B2(n_3),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_176),
.B(n_12),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_245),
.C(n_223),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_202),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_198),
.A2(n_212),
.B1(n_175),
.B2(n_174),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_189),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_193),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_178),
.A2(n_0),
.B1(n_2),
.B2(n_195),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_194),
.A2(n_192),
.B1(n_180),
.B2(n_199),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_230),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_194),
.A2(n_180),
.B1(n_173),
.B2(n_188),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_251),
.B1(n_252),
.B2(n_239),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_248),
.B(n_225),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_197),
.A2(n_190),
.B(n_209),
.C(n_206),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_190),
.A2(n_187),
.B1(n_203),
.B2(n_200),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_187),
.A2(n_203),
.B1(n_200),
.B2(n_201),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_263),
.C(n_260),
.Y(n_289)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_258),
.A2(n_261),
.B1(n_285),
.B2(n_271),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_259),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_233),
.C(n_226),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_266),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_265),
.B(n_261),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_217),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_272),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_236),
.A2(n_220),
.B1(n_218),
.B2(n_216),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_277),
.B(n_284),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

AO22x1_ASAP7_75t_SL g271 ( 
.A1(n_224),
.A2(n_221),
.B1(n_237),
.B2(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_219),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g274 ( 
.A(n_229),
.B(n_232),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_269),
.B(n_273),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_236),
.A2(n_221),
.B1(n_218),
.B2(n_240),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_280),
.B1(n_274),
.B2(n_279),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_218),
.A2(n_235),
.B(n_242),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_241),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_234),
.A2(n_246),
.B1(n_231),
.B2(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_238),
.Y(n_281)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_226),
.B(n_222),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_286),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_239),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_257),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_218),
.A2(n_253),
.B(n_205),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_226),
.B(n_222),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_294),
.C(n_296),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_291),
.A2(n_305),
.B1(n_311),
.B2(n_271),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_258),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_286),
.C(n_263),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_256),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_297),
.B(n_303),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_259),
.C(n_284),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_308),
.C(n_289),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_299),
.A2(n_292),
.B(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_256),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_262),
.A2(n_274),
.B1(n_278),
.B2(n_275),
.Y(n_305)
);

OAI32xp33_ASAP7_75t_L g307 ( 
.A1(n_262),
.A2(n_271),
.A3(n_258),
.B1(n_275),
.B2(n_274),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_269),
.B(n_273),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_277),
.B(n_258),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_281),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_301),
.Y(n_316)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_326),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_318),
.A2(n_306),
.B1(n_290),
.B2(n_307),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_276),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_298),
.C(n_296),
.Y(n_333)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_300),
.Y(n_323)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_313),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_293),
.A2(n_267),
.B1(n_272),
.B2(n_283),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_328),
.B(n_330),
.Y(n_346)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_331),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_312),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_320),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_R g334 ( 
.A(n_326),
.B(n_299),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_334),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_337),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_323),
.A2(n_290),
.B1(n_291),
.B2(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_339),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_329),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_331),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_344),
.B(n_345),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_314),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_325),
.A2(n_304),
.B1(n_292),
.B2(n_308),
.Y(n_347)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_347),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_315),
.C(n_346),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_348),
.B(n_353),
.C(n_354),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_343),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_334),
.A2(n_324),
.B(n_328),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_351),
.A2(n_338),
.B1(n_337),
.B2(n_324),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_314),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_315),
.C(n_330),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_347),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_297),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_359),
.B(n_338),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_362),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_339),
.Y(n_362)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_358),
.Y(n_363)
);

NOR2x1_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_336),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_364),
.A2(n_366),
.B(n_367),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_349),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_343),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_372),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_371),
.B(n_295),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_364),
.A2(n_357),
.B1(n_355),
.B2(n_350),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_375),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_360),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_369),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_377),
.A2(n_374),
.B(n_352),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_365),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_379),
.A2(n_376),
.B(n_368),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_317),
.B(n_340),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_340),
.C(n_341),
.Y(n_382)
);

O2A1O1Ixp33_ASAP7_75t_SL g383 ( 
.A1(n_382),
.A2(n_341),
.B(n_322),
.C(n_321),
.Y(n_383)
);

OAI311xp33_ASAP7_75t_L g384 ( 
.A1(n_383),
.A2(n_335),
.A3(n_332),
.B1(n_327),
.C1(n_351),
.Y(n_384)
);


endmodule