module fake_aes_7794_n_21 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_21;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
BUFx2_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_3), .B(n_4), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
AOI22xp33_ASAP7_75t_SL g15 ( .A1(n_10), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
AO32x1_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_11), .A3(n_15), .B1(n_12), .B2(n_6), .Y(n_18) );
AOI221x1_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_9), .B1(n_12), .B2(n_15), .C(n_1), .Y(n_19) );
OAI22x1_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_16), .B1(n_18), .B2(n_9), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_5), .B(n_3), .Y(n_21) );
endmodule