module fake_netlist_1_12346_n_708 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_708);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_708;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g93 ( .A(n_65), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_18), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_49), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_72), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_48), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_0), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_25), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_22), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_51), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_50), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_69), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_68), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_91), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_78), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_58), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_56), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_18), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_88), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_26), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_11), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_13), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_62), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_59), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_11), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_10), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_0), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_27), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_67), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_10), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_1), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_43), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_66), .Y(n_127) );
CKINVDCx14_ASAP7_75t_R g128 ( .A(n_37), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_24), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_15), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_94), .B(n_1), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_94), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_94), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_113), .Y(n_136) );
XOR2xp5_ASAP7_75t_L g137 ( .A(n_98), .B(n_2), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_110), .B(n_2), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_97), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_93), .B(n_3), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_97), .Y(n_141) );
INVx2_ASAP7_75t_SL g142 ( .A(n_104), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_113), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_113), .B(n_3), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_118), .B(n_4), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_118), .B(n_4), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_109), .Y(n_147) );
AND2x6_ASAP7_75t_L g148 ( .A(n_104), .B(n_20), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_97), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_101), .B(n_5), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_101), .Y(n_151) );
INVxp33_ASAP7_75t_SL g152 ( .A(n_151), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_144), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_151), .B(n_99), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
NAND3xp33_ASAP7_75t_L g156 ( .A(n_144), .B(n_93), .C(n_100), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_139), .Y(n_157) );
XNOR2xp5_ASAP7_75t_L g158 ( .A(n_137), .B(n_109), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_142), .B(n_128), .Y(n_159) );
INVx4_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
INVxp33_ASAP7_75t_L g162 ( .A(n_150), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_144), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_132), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_147), .B(n_102), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
BUFx6f_ASAP7_75t_SL g167 ( .A(n_133), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_142), .B(n_115), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_134), .B(n_115), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_144), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_150), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_133), .A2(n_116), .B1(n_112), .B2(n_119), .Y(n_177) );
OAI22xp33_ASAP7_75t_L g178 ( .A1(n_138), .A2(n_116), .B1(n_112), .B2(n_119), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_135), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_133), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_136), .B(n_95), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
INVx1_ASAP7_75t_SL g184 ( .A(n_176), .Y(n_184) );
NAND3xp33_ASAP7_75t_SL g185 ( .A(n_162), .B(n_137), .C(n_96), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_156), .A2(n_148), .B(n_133), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_165), .B(n_145), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_160), .B(n_145), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_181), .A2(n_146), .B(n_145), .C(n_140), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_153), .Y(n_190) );
O2A1O1Ixp5_ASAP7_75t_L g191 ( .A1(n_160), .A2(n_145), .B(n_146), .C(n_100), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_153), .B(n_146), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_183), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_177), .A2(n_146), .B1(n_148), .B2(n_120), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_159), .B(n_148), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_183), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_164), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_164), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_160), .B(n_107), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_182), .B(n_148), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_181), .A2(n_114), .B(n_126), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_166), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_160), .B(n_136), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_153), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_153), .B(n_148), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_163), .B(n_148), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_163), .B(n_123), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_163), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_167), .A2(n_120), .B1(n_124), .B2(n_125), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_154), .B(n_103), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_163), .B(n_143), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_173), .B(n_143), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_178), .A2(n_125), .B(n_124), .C(n_106), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_173), .B(n_131), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_167), .Y(n_215) );
BUFx8_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_173), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_173), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_158), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_156), .A2(n_131), .B1(n_117), .B2(n_103), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_152), .B(n_105), .Y(n_221) );
BUFx12f_ASAP7_75t_L g222 ( .A(n_158), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_175), .B(n_105), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_175), .A2(n_132), .B1(n_131), .B2(n_115), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_200), .A2(n_180), .B(n_179), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_205), .A2(n_180), .B(n_179), .Y(n_226) );
NOR3xp33_ASAP7_75t_L g227 ( .A(n_185), .B(n_106), .C(n_121), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_206), .A2(n_169), .B(n_170), .Y(n_228) );
OA22x2_ASAP7_75t_L g229 ( .A1(n_184), .A2(n_157), .B1(n_172), .B2(n_171), .Y(n_229) );
INVx2_ASAP7_75t_SL g230 ( .A(n_184), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_210), .B(n_155), .Y(n_231) );
NAND2xp33_ASAP7_75t_L g232 ( .A(n_194), .B(n_155), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_221), .B(n_157), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_194), .B(n_161), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_216), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_195), .A2(n_172), .B(n_171), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_192), .A2(n_168), .B1(n_161), .B2(n_131), .Y(n_237) );
NAND2x1_ASAP7_75t_L g238 ( .A(n_215), .B(n_168), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_187), .B(n_131), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_192), .A2(n_131), .B1(n_117), .B2(n_108), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_222), .B(n_5), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_186), .A2(n_174), .B(n_166), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_219), .B(n_108), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_215), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_188), .A2(n_174), .B(n_114), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_190), .A2(n_114), .B(n_111), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_190), .A2(n_111), .B(n_121), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_216), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_192), .A2(n_126), .B1(n_129), .B2(n_127), .Y(n_249) );
AND2x6_ASAP7_75t_L g250 ( .A(n_192), .B(n_122), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_209), .B(n_122), .Y(n_251) );
OR2x6_ASAP7_75t_L g252 ( .A(n_222), .B(n_219), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_204), .A2(n_130), .B(n_129), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_189), .A2(n_130), .B1(n_127), .B2(n_110), .Y(n_254) );
OAI21xp33_ASAP7_75t_L g255 ( .A1(n_203), .A2(n_122), .B(n_7), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_215), .B(n_6), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_191), .A2(n_6), .B(n_7), .C(n_8), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_229), .A2(n_201), .B(n_214), .Y(n_258) );
AO22x2_ASAP7_75t_L g259 ( .A1(n_254), .A2(n_215), .B1(n_220), .B2(n_214), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_242), .A2(n_212), .B(n_193), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_234), .A2(n_211), .B1(n_208), .B2(n_218), .Y(n_261) );
INVx4_ASAP7_75t_L g262 ( .A(n_244), .Y(n_262) );
AOI21x1_ASAP7_75t_L g263 ( .A1(n_239), .A2(n_193), .B(n_196), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_244), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_230), .B(n_211), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_257), .A2(n_213), .B(n_223), .C(n_207), .Y(n_266) );
AOI221x1_ASAP7_75t_L g267 ( .A1(n_255), .A2(n_218), .B1(n_217), .B2(n_208), .C(n_204), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_231), .A2(n_237), .B1(n_249), .B2(n_256), .Y(n_268) );
AOI221x1_ASAP7_75t_L g269 ( .A1(n_227), .A2(n_217), .B1(n_203), .B2(n_193), .C(n_202), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_228), .A2(n_199), .B(n_202), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_233), .Y(n_271) );
AOI21xp33_ASAP7_75t_L g272 ( .A1(n_243), .A2(n_216), .B(n_222), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_250), .B(n_216), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_244), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_248), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_225), .A2(n_202), .B(n_198), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_226), .A2(n_198), .B(n_197), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_250), .B(n_224), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_232), .A2(n_198), .B(n_197), .Y(n_279) );
NOR4xp25_ASAP7_75t_L g280 ( .A(n_240), .B(n_251), .C(n_235), .D(n_241), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_260), .Y(n_281) );
INVx6_ASAP7_75t_L g282 ( .A(n_262), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_260), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_262), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_265), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_263), .A2(n_253), .B(n_236), .Y(n_286) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_280), .A2(n_246), .B(n_247), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_265), .B(n_250), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_258), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_275), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_270), .A2(n_245), .B(n_238), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_262), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_274), .B(n_250), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_263), .A2(n_196), .B(n_197), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_271), .B(n_196), .Y(n_295) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_267), .A2(n_52), .B(n_92), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_276), .A2(n_252), .B(n_47), .Y(n_297) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_266), .A2(n_252), .B(n_9), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_274), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_258), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_264), .Y(n_302) );
INVxp67_ASAP7_75t_SL g303 ( .A(n_261), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_281), .A2(n_279), .B(n_268), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_285), .B(n_274), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_285), .B(n_273), .Y(n_306) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_281), .A2(n_277), .B(n_278), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_301), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_284), .B(n_292), .Y(n_309) );
INVx5_ASAP7_75t_SL g310 ( .A(n_293), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_301), .Y(n_311) );
OAI221xp5_ASAP7_75t_L g312 ( .A1(n_298), .A2(n_272), .B1(n_275), .B2(n_259), .C(n_269), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_301), .Y(n_313) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_281), .A2(n_267), .B(n_259), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_284), .B(n_259), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_293), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_301), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_284), .B(n_8), .Y(n_319) );
OR2x6_ASAP7_75t_L g320 ( .A(n_298), .B(n_259), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_292), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_289), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_281), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_292), .B(n_269), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_289), .Y(n_325) );
OA21x2_ASAP7_75t_L g326 ( .A1(n_283), .A2(n_53), .B(n_90), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_283), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_288), .B(n_12), .Y(n_328) );
OA21x2_ASAP7_75t_L g329 ( .A1(n_283), .A2(n_46), .B(n_89), .Y(n_329) );
AO21x1_ASAP7_75t_SL g330 ( .A1(n_302), .A2(n_45), .B(n_86), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_282), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_302), .B(n_12), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_303), .B(n_13), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_288), .B(n_14), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_295), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_323), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_322), .B(n_300), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_322), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_325), .B(n_300), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_316), .B(n_300), .Y(n_341) );
BUFx2_ASAP7_75t_SL g342 ( .A(n_331), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_320), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_325), .B(n_300), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_283), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_308), .B(n_303), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_311), .B(n_296), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_316), .B(n_291), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_311), .B(n_296), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_323), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_313), .B(n_296), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_313), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_320), .B(n_287), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_327), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_318), .B(n_296), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_306), .B(n_288), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_327), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_318), .B(n_296), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_307), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_309), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_324), .Y(n_362) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_304), .A2(n_291), .B(n_297), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_307), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_324), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_320), .B(n_296), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_307), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_324), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_320), .B(n_287), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_309), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_332), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_314), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_320), .B(n_287), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_304), .B(n_287), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_336), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_331), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_333), .B(n_287), .Y(n_379) );
OR2x2_ASAP7_75t_SL g380 ( .A(n_333), .B(n_282), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_304), .B(n_294), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_314), .A2(n_297), .B(n_294), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_306), .B(n_290), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_321), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_336), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_314), .B(n_294), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_326), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_319), .B(n_299), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_317), .Y(n_389) );
INVx5_ASAP7_75t_L g390 ( .A(n_310), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_326), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_326), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_319), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_339), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_374), .B(n_305), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_379), .B(n_332), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_369), .B(n_317), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_383), .B(n_315), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_379), .B(n_305), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_369), .B(n_317), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_369), .B(n_317), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_374), .B(n_328), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_360), .B(n_317), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_337), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_379), .B(n_334), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_375), .B(n_334), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_390), .B(n_328), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_373), .B(n_310), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_373), .B(n_341), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_378), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_343), .A2(n_312), .B1(n_293), .B2(n_310), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_375), .B(n_310), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_377), .B(n_299), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_357), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_339), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_341), .B(n_330), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_337), .Y(n_417) );
INVx1_ASAP7_75t_SL g418 ( .A(n_342), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_341), .B(n_330), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_341), .B(n_329), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_383), .B(n_14), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_341), .B(n_329), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_354), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_377), .B(n_299), .Y(n_424) );
NOR2xp67_ASAP7_75t_L g425 ( .A(n_390), .B(n_15), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_378), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_360), .B(n_362), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_370), .B(n_329), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_362), .B(n_329), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_365), .B(n_326), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_393), .B(n_282), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_370), .B(n_286), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_365), .B(n_286), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_361), .B(n_286), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_393), .B(n_282), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_384), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_352), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_384), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_368), .B(n_16), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_368), .B(n_16), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_352), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_348), .B(n_17), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_348), .B(n_17), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_348), .B(n_19), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_354), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_348), .B(n_19), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_361), .B(n_293), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_348), .B(n_293), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_385), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_343), .B(n_293), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_371), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_371), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_390), .B(n_282), .Y(n_453) );
NAND2x1_ASAP7_75t_L g454 ( .A(n_357), .B(n_282), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_346), .B(n_21), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_361), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_346), .B(n_23), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_388), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_353), .B(n_28), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_378), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_338), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_338), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_346), .B(n_29), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_356), .B(n_30), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_343), .B(n_31), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_366), .B(n_32), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_338), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_356), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_340), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_380), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_366), .B(n_36), .Y(n_471) );
AND2x4_ASAP7_75t_SL g472 ( .A(n_345), .B(n_38), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_436), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_409), .B(n_397), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_409), .B(n_389), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_405), .B(n_380), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_394), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_394), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_415), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_470), .B(n_353), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_417), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_417), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_400), .B(n_389), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_400), .B(n_353), .Y(n_485) );
INVx3_ASAP7_75t_SL g486 ( .A(n_418), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_404), .Y(n_487) );
BUFx3_ASAP7_75t_L g488 ( .A(n_410), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_415), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_401), .B(n_345), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_401), .B(n_366), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_470), .B(n_342), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_437), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_398), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_408), .B(n_340), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_437), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_451), .B(n_376), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_452), .B(n_376), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_441), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_404), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_461), .B(n_376), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_423), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_445), .Y(n_503) );
INVxp67_ASAP7_75t_SL g504 ( .A(n_445), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_461), .B(n_344), .Y(n_505) );
OR2x6_ASAP7_75t_L g506 ( .A(n_410), .B(n_388), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_462), .B(n_344), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_449), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_449), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_448), .B(n_344), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_421), .B(n_388), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_427), .B(n_390), .Y(n_512) );
AND2x4_ASAP7_75t_L g513 ( .A(n_427), .B(n_390), .Y(n_513) );
NOR2x1p5_ASAP7_75t_L g514 ( .A(n_454), .B(n_392), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_448), .B(n_357), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_399), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_426), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_399), .B(n_396), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_462), .B(n_386), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_442), .B(n_357), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_396), .B(n_467), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_426), .B(n_460), .Y(n_522) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_453), .B(n_390), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_442), .B(n_357), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_395), .B(n_390), .Y(n_525) );
NAND2x1_ASAP7_75t_L g526 ( .A(n_416), .B(n_350), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_443), .B(n_350), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_467), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_469), .B(n_367), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_443), .B(n_386), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_469), .B(n_367), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_444), .A2(n_390), .B1(n_349), .B2(n_347), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_458), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_460), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_444), .B(n_386), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_456), .B(n_364), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_413), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_402), .B(n_39), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_416), .B(n_419), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_446), .B(n_347), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_406), .B(n_364), .Y(n_541) );
INVxp67_ASAP7_75t_SL g542 ( .A(n_428), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_424), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_446), .B(n_364), .C(n_359), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_432), .B(n_359), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_432), .B(n_359), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_431), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_435), .Y(n_548) );
AND3x1_ASAP7_75t_L g549 ( .A(n_465), .B(n_372), .C(n_349), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_419), .B(n_367), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_447), .B(n_372), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_433), .B(n_372), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_447), .B(n_347), .Y(n_553) );
NAND4xp25_ASAP7_75t_L g554 ( .A(n_411), .B(n_381), .C(n_351), .D(n_355), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_450), .B(n_381), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_516), .B(n_433), .Y(n_556) );
OAI22xp5_ASAP7_75t_SL g557 ( .A1(n_549), .A2(n_459), .B1(n_450), .B2(n_412), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_521), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_547), .B(n_440), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_486), .B(n_464), .Y(n_560) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_482), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_475), .B(n_450), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_518), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_548), .B(n_440), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_473), .Y(n_565) );
BUFx2_ASAP7_75t_L g566 ( .A(n_488), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_474), .Y(n_567) );
AOI21xp33_ASAP7_75t_L g568 ( .A1(n_538), .A2(n_439), .B(n_459), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_537), .B(n_439), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_476), .B(n_403), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_517), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_545), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_485), .B(n_403), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_542), .B(n_429), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_508), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_509), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_543), .B(n_429), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_499), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_490), .B(n_471), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_542), .B(n_430), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_534), .Y(n_581) );
OAI32xp33_ASAP7_75t_L g582 ( .A1(n_477), .A2(n_407), .A3(n_428), .B1(n_465), .B2(n_434), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_519), .B(n_434), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_478), .Y(n_584) );
OR2x6_ASAP7_75t_L g585 ( .A(n_492), .B(n_471), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_491), .B(n_466), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_495), .B(n_466), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_479), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_519), .B(n_414), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_511), .A2(n_425), .B1(n_463), .B2(n_457), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_501), .B(n_414), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_480), .Y(n_592) );
NAND2x1_ASAP7_75t_L g593 ( .A(n_492), .B(n_414), .Y(n_593) );
AOI32xp33_ASAP7_75t_L g594 ( .A1(n_549), .A2(n_472), .A3(n_455), .B1(n_463), .B2(n_457), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_526), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_489), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_554), .A2(n_455), .B1(n_472), .B2(n_422), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_497), .B(n_422), .Y(n_598) );
NOR2xp33_ASAP7_75t_R g599 ( .A(n_494), .B(n_420), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_522), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_493), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_553), .B(n_420), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_546), .Y(n_603) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_539), .B(n_392), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_528), .B(n_349), .Y(n_605) );
AOI21xp33_ASAP7_75t_SL g606 ( .A1(n_492), .A2(n_468), .B(n_392), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_496), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_555), .B(n_358), .Y(n_608) );
AOI32xp33_ASAP7_75t_L g609 ( .A1(n_539), .A2(n_358), .A3(n_355), .B1(n_351), .B2(n_391), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_555), .B(n_358), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_541), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_533), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_497), .B(n_382), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_498), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_484), .B(n_382), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_552), .B(n_363), .Y(n_616) );
NAND4xp75_ASAP7_75t_L g617 ( .A(n_525), .B(n_391), .C(n_387), .D(n_363), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_483), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_506), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_498), .B(n_382), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_552), .B(n_363), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_606), .B(n_554), .C(n_544), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_614), .B(n_530), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_557), .A2(n_481), .B1(n_544), .B2(n_506), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_574), .B(n_551), .Y(n_625) );
XNOR2xp5_ASAP7_75t_L g626 ( .A(n_566), .B(n_535), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_578), .Y(n_627) );
NAND2x1_ASAP7_75t_L g628 ( .A(n_585), .B(n_506), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_571), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_611), .B(n_510), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_567), .B(n_540), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_575), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_557), .A2(n_523), .B(n_504), .Y(n_633) );
OAI31xp33_ASAP7_75t_SL g634 ( .A1(n_600), .A2(n_512), .A3(n_513), .B(n_504), .Y(n_634) );
AO22x1_ASAP7_75t_L g635 ( .A1(n_595), .A2(n_513), .B1(n_512), .B2(n_550), .Y(n_635) );
OAI31xp33_ASAP7_75t_L g636 ( .A1(n_600), .A2(n_523), .A3(n_514), .B(n_550), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_576), .Y(n_637) );
CKINVDCx16_ASAP7_75t_R g638 ( .A(n_599), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_581), .B(n_503), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_573), .B(n_515), .Y(n_640) );
AOI32xp33_ASAP7_75t_L g641 ( .A1(n_561), .A2(n_520), .A3(n_524), .B1(n_527), .B2(n_507), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_612), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_563), .B(n_503), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_580), .B(n_558), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_562), .Y(n_645) );
OAI311xp33_ASAP7_75t_L g646 ( .A1(n_597), .A2(n_532), .A3(n_536), .B1(n_531), .C1(n_529), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g647 ( .A1(n_585), .A2(n_532), .B1(n_505), .B2(n_500), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_585), .A2(n_505), .B1(n_487), .B2(n_502), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_590), .A2(n_387), .B1(n_382), .B2(n_363), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_594), .B(n_604), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_565), .B(n_382), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_584), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_590), .A2(n_387), .B1(n_363), .B2(n_41), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_570), .B(n_40), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_619), .B(n_42), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g656 ( .A1(n_568), .A2(n_44), .B(n_54), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_588), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_592), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_622), .A2(n_582), .B1(n_609), .B2(n_615), .C(n_568), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_638), .A2(n_560), .B1(n_577), .B2(n_569), .Y(n_660) );
O2A1O1Ixp5_ASAP7_75t_L g661 ( .A1(n_650), .A2(n_593), .B(n_620), .C(n_613), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_633), .A2(n_617), .B(n_621), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_647), .A2(n_564), .B1(n_559), .B2(n_556), .Y(n_663) );
AO22x2_ASAP7_75t_L g664 ( .A1(n_629), .A2(n_596), .B1(n_601), .B2(n_607), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_634), .B(n_603), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_624), .A2(n_602), .B1(n_583), .B2(n_579), .Y(n_666) );
OAI21xp33_ASAP7_75t_SL g667 ( .A1(n_634), .A2(n_587), .B(n_586), .Y(n_667) );
NAND2xp33_ASAP7_75t_SL g668 ( .A(n_628), .B(n_589), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_644), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_635), .A2(n_620), .B(n_613), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_646), .A2(n_598), .B1(n_572), .B2(n_616), .C(n_618), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_639), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_626), .A2(n_591), .B1(n_610), .B2(n_608), .Y(n_673) );
AOI322xp5_ASAP7_75t_L g674 ( .A1(n_645), .A2(n_605), .A3(n_57), .B1(n_60), .B2(n_61), .C1(n_63), .C2(n_64), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_648), .A2(n_55), .B1(n_70), .B2(n_71), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_649), .A2(n_73), .B(n_75), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_641), .A2(n_76), .B(n_77), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_651), .B(n_79), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_636), .B(n_80), .C(n_81), .D(n_82), .Y(n_679) );
NAND3xp33_ASAP7_75t_SL g680 ( .A(n_656), .B(n_83), .C(n_85), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_625), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_653), .A2(n_642), .B(n_627), .C(n_658), .Y(n_682) );
AOI221xp5_ASAP7_75t_SL g683 ( .A1(n_631), .A2(n_643), .B1(n_630), .B2(n_623), .C(n_637), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_632), .A2(n_652), .B1(n_657), .B2(n_640), .C(n_654), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_655), .A2(n_634), .B1(n_624), .B2(n_650), .C(n_622), .Y(n_685) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_634), .A2(n_624), .B(n_650), .C(n_636), .Y(n_686) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_686), .B(n_679), .Y(n_687) );
AND4x1_ASAP7_75t_L g688 ( .A(n_659), .B(n_661), .C(n_677), .D(n_682), .Y(n_688) );
OA211x2_ASAP7_75t_L g689 ( .A1(n_662), .A2(n_672), .B(n_684), .C(n_671), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_685), .A2(n_667), .B(n_666), .C(n_675), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_683), .B(n_669), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_667), .B(n_660), .Y(n_692) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_687), .B(n_680), .Y(n_693) );
BUFx12f_ASAP7_75t_L g694 ( .A(n_689), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_690), .B(n_692), .C(n_691), .D(n_674), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_688), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_696), .B(n_664), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_693), .B(n_665), .Y(n_698) );
AND2x4_ASAP7_75t_L g699 ( .A(n_694), .B(n_681), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_699), .B(n_668), .Y(n_700) );
XNOR2xp5_ASAP7_75t_L g701 ( .A(n_699), .B(n_695), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_701), .Y(n_702) );
XNOR2xp5_ASAP7_75t_L g703 ( .A(n_700), .B(n_697), .Y(n_703) );
OAI21xp5_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_698), .B(n_673), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_704), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_705), .B(n_702), .Y(n_706) );
AO21x2_ASAP7_75t_L g707 ( .A1(n_706), .A2(n_663), .B(n_670), .Y(n_707) );
AO21x2_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_678), .B(n_676), .Y(n_708) );
endmodule