module real_aes_1644_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_0), .B(n_219), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_1), .A2(n_214), .B(n_261), .Y(n_260) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_2), .A2(n_54), .B1(n_92), .B2(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_3), .B(n_230), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_3), .A2(n_82), .B1(n_83), .B2(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_3), .Y(n_511) );
INVx1_ASAP7_75t_L g194 ( .A(n_4), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_5), .B(n_230), .Y(n_269) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_6), .A2(n_22), .B1(n_92), .B2(n_102), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_7), .B(n_228), .Y(n_281) );
INVx2_ASAP7_75t_L g211 ( .A(n_8), .Y(n_211) );
AOI221x1_ASAP7_75t_L g213 ( .A1(n_9), .A2(n_16), .B1(n_214), .B2(n_219), .C(n_226), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_10), .A2(n_51), .B1(n_123), .B2(n_126), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_11), .B(n_219), .Y(n_277) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_12), .A2(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_13), .B(n_209), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_14), .B(n_230), .Y(n_289) );
AO21x1_ASAP7_75t_L g300 ( .A1(n_15), .A2(n_219), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g532 ( .A(n_15), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g86 ( .A1(n_17), .A2(n_59), .B1(n_87), .B2(n_106), .Y(n_86) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_18), .A2(n_49), .B1(n_140), .B2(n_143), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_19), .A2(n_33), .B1(n_166), .B2(n_170), .Y(n_165) );
NAND2x1_ASAP7_75t_L g238 ( .A(n_20), .B(n_230), .Y(n_238) );
NAND2x1_ASAP7_75t_L g268 ( .A(n_21), .B(n_228), .Y(n_268) );
OAI221xp5_ASAP7_75t_L g186 ( .A1(n_22), .A2(n_54), .B1(n_60), .B2(n_187), .C(n_189), .Y(n_186) );
OR2x2_ASAP7_75t_L g212 ( .A(n_23), .B(n_67), .Y(n_212) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_23), .A2(n_67), .B(n_211), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_24), .B(n_228), .Y(n_263) );
INVx3_ASAP7_75t_L g92 ( .A(n_25), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_26), .B(n_230), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_27), .B(n_228), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_28), .A2(n_214), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_SL g97 ( .A(n_29), .Y(n_97) );
INVx1_ASAP7_75t_L g196 ( .A(n_30), .Y(n_196) );
AND2x2_ASAP7_75t_L g215 ( .A(n_30), .B(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g225 ( .A(n_30), .B(n_194), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_31), .B(n_219), .Y(n_252) );
OAI22xp5_ASAP7_75t_SL g180 ( .A1(n_32), .A2(n_45), .B1(n_181), .B2(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_32), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_34), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_35), .B(n_228), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_36), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_37), .A2(n_214), .B(n_267), .Y(n_266) );
AO22x2_ASAP7_75t_L g91 ( .A1(n_38), .A2(n_60), .B1(n_92), .B2(n_93), .Y(n_91) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_39), .A2(n_46), .B1(n_177), .B2(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g178 ( .A(n_39), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_40), .A2(n_82), .B1(n_83), .B2(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_40), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_41), .B(n_228), .Y(n_239) );
INVx1_ASAP7_75t_L g218 ( .A(n_42), .Y(n_218) );
INVx1_ASAP7_75t_L g222 ( .A(n_42), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g156 ( .A1(n_43), .A2(n_66), .B1(n_157), .B2(n_160), .Y(n_156) );
INVx1_ASAP7_75t_L g98 ( .A(n_44), .Y(n_98) );
INVx1_ASAP7_75t_L g181 ( .A(n_45), .Y(n_181) );
INVx1_ASAP7_75t_L g177 ( .A(n_46), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_46), .B(n_230), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_47), .A2(n_74), .B1(n_131), .B2(n_134), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_48), .A2(n_214), .B(n_237), .Y(n_236) );
AO21x1_ASAP7_75t_L g302 ( .A1(n_50), .A2(n_214), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_52), .B(n_219), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_53), .B(n_219), .Y(n_270) );
INVxp33_ASAP7_75t_L g191 ( .A(n_54), .Y(n_191) );
AND2x2_ASAP7_75t_L g253 ( .A(n_55), .B(n_210), .Y(n_253) );
INVx1_ASAP7_75t_L g216 ( .A(n_56), .Y(n_216) );
INVx1_ASAP7_75t_L g224 ( .A(n_56), .Y(n_224) );
AND2x2_ASAP7_75t_L g272 ( .A(n_57), .B(n_242), .Y(n_272) );
INVx1_ASAP7_75t_L g81 ( .A(n_58), .Y(n_81) );
INVxp67_ASAP7_75t_L g190 ( .A(n_60), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_61), .A2(n_63), .B1(n_114), .B2(n_118), .Y(n_113) );
AND2x2_ASAP7_75t_L g257 ( .A(n_62), .B(n_242), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_64), .B(n_219), .Y(n_291) );
AND2x2_ASAP7_75t_L g301 ( .A(n_65), .B(n_282), .Y(n_301) );
AND2x2_ASAP7_75t_L g245 ( .A(n_68), .B(n_242), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_69), .B(n_228), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_70), .B(n_230), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_71), .B(n_228), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_72), .A2(n_214), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_73), .B(n_230), .Y(n_262) );
BUFx2_ASAP7_75t_SL g188 ( .A(n_75), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_76), .A2(n_214), .B(n_279), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_183), .B1(n_197), .B2(n_505), .C(n_509), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_174), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NOR2x1_ASAP7_75t_L g84 ( .A(n_85), .B(n_138), .Y(n_84) );
NAND4xp25_ASAP7_75t_L g85 ( .A(n_86), .B(n_113), .C(n_122), .D(n_130), .Y(n_85) );
BUFx3_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
BUFx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_99), .Y(n_89) );
AND2x2_ASAP7_75t_L g125 ( .A(n_90), .B(n_111), .Y(n_125) );
AND2x4_ASAP7_75t_L g169 ( .A(n_90), .B(n_137), .Y(n_169) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_94), .Y(n_90) );
INVx2_ASAP7_75t_L g110 ( .A(n_91), .Y(n_110) );
BUFx2_ASAP7_75t_L g129 ( .A(n_91), .Y(n_129) );
AND2x2_ASAP7_75t_L g147 ( .A(n_91), .B(n_95), .Y(n_147) );
INVx1_ASAP7_75t_L g93 ( .A(n_92), .Y(n_93) );
OAI22x1_ASAP7_75t_L g95 ( .A1(n_92), .A2(n_96), .B1(n_97), .B2(n_98), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
INVx2_ASAP7_75t_L g102 ( .A(n_92), .Y(n_102) );
INVx1_ASAP7_75t_L g105 ( .A(n_92), .Y(n_105) );
AND2x4_ASAP7_75t_L g109 ( .A(n_94), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
AND2x2_ASAP7_75t_L g117 ( .A(n_95), .B(n_110), .Y(n_117) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_95), .Y(n_164) );
AND2x4_ASAP7_75t_L g116 ( .A(n_99), .B(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g133 ( .A(n_99), .B(n_109), .Y(n_133) );
AND2x2_ASAP7_75t_L g155 ( .A(n_99), .B(n_147), .Y(n_155) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_103), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g112 ( .A(n_101), .Y(n_112) );
AND2x2_ASAP7_75t_L g121 ( .A(n_101), .B(n_104), .Y(n_121) );
AND2x4_ASAP7_75t_L g137 ( .A(n_101), .B(n_103), .Y(n_137) );
INVxp67_ASAP7_75t_L g173 ( .A(n_103), .Y(n_173) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g111 ( .A(n_104), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx8_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND2x4_ASAP7_75t_L g120 ( .A(n_109), .B(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g136 ( .A(n_109), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g142 ( .A(n_111), .B(n_117), .Y(n_142) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_112), .Y(n_149) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx6_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g159 ( .A(n_117), .B(n_137), .Y(n_159) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g128 ( .A(n_121), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g163 ( .A(n_121), .B(n_164), .Y(n_163) );
BUFx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx5_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
INVx3_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
INVx8_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND4xp25_ASAP7_75t_L g138 ( .A(n_139), .B(n_150), .C(n_156), .D(n_165), .Y(n_138) );
BUFx6f_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g172 ( .A(n_147), .B(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_SL g153 ( .A(n_154), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx12f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx6_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B1(n_179), .B2(n_180), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
AND3x1_ASAP7_75t_SL g185 ( .A(n_186), .B(n_192), .C(n_195), .Y(n_185) );
INVxp67_ASAP7_75t_L g517 ( .A(n_186), .Y(n_517) );
CKINVDCx8_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_192), .Y(n_515) );
AO21x1_ASAP7_75t_SL g525 ( .A1(n_192), .A2(n_526), .B(n_530), .Y(n_525) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OR2x2_ASAP7_75t_SL g522 ( .A(n_193), .B(n_195), .Y(n_522) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g217 ( .A(n_194), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_195), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2x1p5_ASAP7_75t_L g527 ( .A(n_196), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_417), .Y(n_200) );
AND4x1_ASAP7_75t_L g201 ( .A(n_202), .B(n_329), .C(n_356), .D(n_391), .Y(n_201) );
AOI221xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_254), .B1(n_294), .B2(n_309), .C(n_313), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_233), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_205), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g370 ( .A(n_206), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g425 ( .A(n_206), .B(n_380), .Y(n_425) );
BUFx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g328 ( .A(n_207), .B(n_246), .Y(n_328) );
AND2x4_ASAP7_75t_L g364 ( .A(n_207), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g378 ( .A(n_207), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g295 ( .A(n_208), .Y(n_295) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_208), .Y(n_467) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_213), .B(n_232), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_209), .A2(n_259), .B(n_260), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_209), .Y(n_271) );
OA21x2_ASAP7_75t_L g341 ( .A1(n_209), .A2(n_213), .B(n_232), .Y(n_341) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AND2x4_ASAP7_75t_L g282 ( .A(n_211), .B(n_212), .Y(n_282) );
AND2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
AND2x6_ASAP7_75t_L g228 ( .A(n_216), .B(n_221), .Y(n_228) );
INVx2_ASAP7_75t_L g529 ( .A(n_216), .Y(n_529) );
AND2x4_ASAP7_75t_L g230 ( .A(n_218), .B(n_223), .Y(n_230) );
INVx2_ASAP7_75t_L g531 ( .A(n_218), .Y(n_531) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_219), .Y(n_508) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_225), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_223), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx5_ASAP7_75t_L g231 ( .A(n_225), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_229), .B(n_231), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_231), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_231), .A2(n_250), .B(n_251), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_231), .A2(n_262), .B(n_263), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_231), .A2(n_268), .B(n_269), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_231), .A2(n_280), .B(n_281), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_231), .A2(n_289), .B(n_290), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_231), .A2(n_304), .B(n_305), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_SL g322 ( .A1(n_233), .A2(n_295), .B(n_323), .C(n_327), .Y(n_322) );
AND2x2_ASAP7_75t_L g343 ( .A(n_233), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_233), .B(n_295), .Y(n_483) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_246), .Y(n_233) );
INVx2_ASAP7_75t_L g363 ( .A(n_234), .Y(n_363) );
BUFx3_ASAP7_75t_L g379 ( .A(n_234), .Y(n_379) );
INVxp67_ASAP7_75t_L g383 ( .A(n_234), .Y(n_383) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_241), .B(n_245), .Y(n_234) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_235), .A2(n_241), .B(n_245), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_240), .Y(n_235) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_241), .A2(n_247), .B(n_253), .Y(n_246) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_241), .A2(n_247), .B(n_253), .Y(n_308) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx4_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx4f_ASAP7_75t_L g275 ( .A(n_244), .Y(n_275) );
INVx2_ASAP7_75t_L g362 ( .A(n_246), .Y(n_362) );
AND2x2_ASAP7_75t_L g368 ( .A(n_246), .B(n_341), .Y(n_368) );
AND2x2_ASAP7_75t_L g394 ( .A(n_246), .B(n_363), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_248), .B(n_252), .Y(n_247) );
AOI211xp5_ASAP7_75t_L g391 ( .A1(n_254), .A2(n_392), .B(n_395), .C(n_405), .Y(n_391) );
AND2x2_ASAP7_75t_SL g254 ( .A(n_255), .B(n_273), .Y(n_254) );
OAI321xp33_ASAP7_75t_L g366 ( .A1(n_255), .A2(n_314), .A3(n_367), .B1(n_369), .B2(n_370), .C(n_372), .Y(n_366) );
AND2x2_ASAP7_75t_L g487 ( .A(n_255), .B(n_462), .Y(n_487) );
INVx1_ASAP7_75t_L g490 ( .A(n_255), .Y(n_490) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_264), .Y(n_255) );
INVx5_ASAP7_75t_L g312 ( .A(n_256), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_256), .B(n_326), .Y(n_325) );
NOR2x1_ASAP7_75t_SL g357 ( .A(n_256), .B(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g402 ( .A(n_256), .Y(n_402) );
AND2x2_ASAP7_75t_L g504 ( .A(n_256), .B(n_274), .Y(n_504) );
OR2x6_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g311 ( .A(n_264), .B(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_264), .Y(n_321) );
INVx4_ASAP7_75t_L g326 ( .A(n_264), .Y(n_326) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_271), .B(n_272), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_270), .Y(n_265) );
INVx1_ASAP7_75t_L g369 ( .A(n_273), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_R g472 ( .A1(n_273), .A2(n_311), .B(n_343), .C(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g492 ( .A(n_273), .B(n_317), .Y(n_492) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_283), .Y(n_273) );
INVx1_ASAP7_75t_L g310 ( .A(n_274), .Y(n_310) );
INVx2_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
OR2x2_ASAP7_75t_L g335 ( .A(n_274), .B(n_326), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_274), .B(n_358), .Y(n_404) );
BUFx3_ASAP7_75t_L g411 ( .A(n_274), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B(n_282), .Y(n_276) );
INVx1_ASAP7_75t_SL g285 ( .A(n_282), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_282), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g374 ( .A(n_283), .Y(n_374) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_283), .Y(n_387) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g320 ( .A(n_284), .Y(n_320) );
INVx1_ASAP7_75t_L g429 ( .A(n_284), .Y(n_429) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_292), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_285), .B(n_293), .Y(n_292) );
AO21x2_ASAP7_75t_L g358 ( .A1(n_285), .A2(n_286), .B(n_292), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
AND2x2_ASAP7_75t_L g330 ( .A(n_294), .B(n_331), .Y(n_330) );
OAI31xp33_ASAP7_75t_L g481 ( .A1(n_294), .A2(n_482), .A3(n_484), .B(n_487), .Y(n_481) );
INVx1_ASAP7_75t_SL g499 ( .A(n_294), .Y(n_499) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_295), .A2(n_314), .B(n_322), .Y(n_313) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_295), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g422 ( .A(n_295), .Y(n_422) );
INVx2_ASAP7_75t_L g371 ( .A(n_296), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_296), .B(n_354), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_296), .B(n_353), .Y(n_463) );
NOR2xp33_ASAP7_75t_SL g471 ( .A(n_296), .B(n_422), .Y(n_471) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_308), .Y(n_296) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_297), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g351 ( .A(n_297), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g380 ( .A(n_297), .B(n_362), .Y(n_380) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_L g344 ( .A(n_298), .Y(n_344) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g365 ( .A(n_299), .Y(n_365) );
OAI21x1_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .B(n_306), .Y(n_299) );
INVx1_ASAP7_75t_L g307 ( .A(n_301), .Y(n_307) );
INVx2_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_308), .Y(n_412) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g348 ( .A(n_310), .Y(n_348) );
AND2x2_ASAP7_75t_L g427 ( .A(n_310), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g338 ( .A(n_311), .B(n_332), .Y(n_338) );
INVx2_ASAP7_75t_SL g386 ( .A(n_311), .Y(n_386) );
INVx4_ASAP7_75t_L g317 ( .A(n_312), .Y(n_317) );
AND2x2_ASAP7_75t_L g415 ( .A(n_312), .B(n_358), .Y(n_415) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_312), .B(n_428), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g450 ( .A(n_312), .B(n_326), .Y(n_450) );
INVx1_ASAP7_75t_L g456 ( .A(n_314), .Y(n_456) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
INVx1_ASAP7_75t_L g375 ( .A(n_315), .Y(n_375) );
OR2x2_ASAP7_75t_L g388 ( .A(n_315), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
OR2x2_ASAP7_75t_L g440 ( .A(n_316), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g470 ( .A(n_316), .B(n_358), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_317), .B(n_320), .Y(n_346) );
AND2x2_ASAP7_75t_L g438 ( .A(n_317), .B(n_428), .Y(n_438) );
AND2x4_ASAP7_75t_L g500 ( .A(n_317), .B(n_379), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx2_ASAP7_75t_L g324 ( .A(n_319), .Y(n_324) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp67_ASAP7_75t_SL g323 ( .A(n_324), .B(n_325), .Y(n_323) );
OAI322xp33_ASAP7_75t_SL g336 ( .A1(n_324), .A2(n_337), .A3(n_339), .B1(n_342), .B2(n_345), .C1(n_347), .C2(n_349), .Y(n_336) );
INVx1_ASAP7_75t_L g494 ( .A(n_324), .Y(n_494) );
OR2x2_ASAP7_75t_L g347 ( .A(n_325), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g373 ( .A(n_326), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_326), .B(n_374), .Y(n_389) );
INVx2_ASAP7_75t_L g416 ( .A(n_326), .Y(n_416) );
AND2x4_ASAP7_75t_L g428 ( .A(n_326), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_328), .B(n_344), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_334), .B(n_336), .Y(n_329) );
AND2x2_ASAP7_75t_L g397 ( .A(n_331), .B(n_364), .Y(n_397) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_332), .B(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g355 ( .A(n_333), .Y(n_355) );
AND2x4_ASAP7_75t_SL g437 ( .A(n_333), .B(n_352), .Y(n_437) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g345 ( .A(n_335), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_338), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g473 ( .A(n_340), .B(n_437), .Y(n_473) );
NOR4xp25_ASAP7_75t_L g477 ( .A(n_340), .B(n_354), .C(n_394), .D(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g354 ( .A(n_341), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g390 ( .A(n_341), .B(n_365), .Y(n_390) );
AND2x4_ASAP7_75t_L g454 ( .A(n_341), .B(n_365), .Y(n_454) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_344), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
OR2x2_ASAP7_75t_L g443 ( .A(n_351), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g497 ( .A(n_351), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_352), .B(n_364), .Y(n_398) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AOI211xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_359), .B(n_366), .C(n_381), .Y(n_356) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_364), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_362), .B(n_365), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_363), .B(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g445 ( .A(n_363), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_364), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g460 ( .A(n_364), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_375), .B(n_376), .Y(n_372) );
AND2x4_ASAP7_75t_L g409 ( .A(n_373), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g503 ( .A(n_373), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_SL g407 ( .A(n_379), .Y(n_407) );
AND2x2_ASAP7_75t_L g466 ( .A(n_380), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g480 ( .A(n_380), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_384), .B(n_388), .C(n_390), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_382), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g458 ( .A(n_383), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g479 ( .A(n_383), .B(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
OR2x2_ASAP7_75t_L g468 ( .A(n_386), .B(n_410), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_389), .A2(n_396), .B1(n_398), .B2(n_399), .Y(n_395) );
INVx1_ASAP7_75t_SL g486 ( .A(n_390), .Y(n_486) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_401), .B(n_410), .Y(n_452) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_404), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B1(n_412), .B2(n_413), .Y(n_405) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI21xp5_ASAP7_75t_SL g419 ( .A1(n_410), .A2(n_420), .B(n_423), .Y(n_419) );
AND2x2_ASAP7_75t_L g448 ( .A(n_410), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND3x2_ASAP7_75t_L g414 ( .A(n_411), .B(n_415), .C(n_416), .Y(n_414) );
AND2x2_ASAP7_75t_L g476 ( .A(n_411), .B(n_433), .Y(n_476) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g461 ( .A(n_416), .B(n_462), .Y(n_461) );
NOR2xp67_ASAP7_75t_L g417 ( .A(n_418), .B(n_474), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_419), .B(n_434), .C(n_455), .D(n_472), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_430), .B2(n_432), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_426), .A2(n_440), .B1(n_460), .B2(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g441 ( .A(n_428), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_430), .A2(n_453), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx3_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_438), .B1(n_439), .B2(n_442), .C(n_446), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_451), .B1(n_452), .B2(n_453), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_449), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_449), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_461), .B2(n_463), .C(n_464), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_458), .B(n_460), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_468), .B1(n_469), .B2(n_471), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI211xp5_ASAP7_75t_SL g489 ( .A1(n_470), .A2(n_490), .B(n_491), .C(n_493), .Y(n_489) );
OAI211xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_477), .B(n_481), .C(n_488), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_495), .B1(n_498), .B2(n_500), .C(n_501), .Y(n_488) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI222xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_512), .B1(n_518), .B2(n_520), .C1(n_523), .C2(n_532), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
endmodule