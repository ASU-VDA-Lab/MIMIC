module real_jpeg_11236_n_16 (n_5, n_4, n_8, n_0, n_12, n_339, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_340, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_339;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_340;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_1),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_1),
.A2(n_48),
.B1(n_50),
.B2(n_60),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_60),
.Y(n_265)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_3),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_3),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_3),
.A2(n_48),
.B1(n_50),
.B2(n_62),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_4),
.A2(n_50),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_4),
.B(n_50),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_4),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_4),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_4),
.B(n_26),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_4),
.A2(n_28),
.B(n_30),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_4),
.A2(n_23),
.B1(n_25),
.B2(n_113),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_5),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_50),
.B(n_65),
.C(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_7),
.B(n_50),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_10),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_10),
.A2(n_24),
.B1(n_48),
.B2(n_50),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_24),
.B1(n_67),
.B2(n_68),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_34),
.B1(n_67),
.B2(n_68),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_11),
.A2(n_34),
.B1(n_48),
.B2(n_50),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_13),
.A2(n_48),
.B1(n_50),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_13),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_104),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_104),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_13),
.A2(n_23),
.B1(n_25),
.B2(n_104),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_14),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_14),
.A2(n_48),
.B1(n_50),
.B2(n_92),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_92),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_14),
.A2(n_23),
.B1(n_25),
.B2(n_92),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_15),
.A2(n_67),
.B1(n_68),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_15),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_15),
.A2(n_48),
.B1(n_50),
.B2(n_97),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_97),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_15),
.A2(n_23),
.B1(n_25),
.B2(n_97),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_337),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_79),
.B(n_335),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_20),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_21),
.A2(n_36),
.B(n_238),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_22),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_22),
.A2(n_26),
.B(n_35),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_27),
.B(n_31),
.C(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_31),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_23),
.A2(n_31),
.B(n_113),
.C(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_26),
.B(n_33),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_26),
.A2(n_35),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_27),
.A2(n_36),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_27),
.A2(n_36),
.B1(n_210),
.B2(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_27),
.A2(n_36),
.B1(n_219),
.B2(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_27),
.A2(n_32),
.B(n_59),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_45),
.B(n_46),
.C(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_46),
.Y(n_54)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_30),
.B(n_113),
.CON(n_143),
.SN(n_143)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_35),
.A2(n_74),
.B(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_36),
.A2(n_76),
.B(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_39),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_73),
.C(n_77),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_40),
.A2(n_41),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_57),
.C(n_63),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_42),
.A2(n_43),
.B1(n_63),
.B2(n_310),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_52),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_44),
.A2(n_162),
.B(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_51),
.B(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_45),
.A2(n_53),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_45),
.A2(n_53),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_46),
.B(n_50),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_48),
.A2(n_54),
.B1(n_143),
.B2(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_51),
.A2(n_53),
.B(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_52),
.A2(n_129),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_53),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_56),
.B(n_129),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_57),
.A2(n_58),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_63),
.A2(n_307),
.B1(n_310),
.B2(n_311),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_63),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_71),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_66),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_64),
.A2(n_66),
.B1(n_103),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_64),
.A2(n_66),
.B1(n_131),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_64),
.A2(n_141),
.B(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_64),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_64),
.A2(n_66),
.B1(n_225),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_64),
.A2(n_245),
.B(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_66),
.B(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_66),
.B(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_66),
.A2(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_67),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_67),
.B(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_67),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_72),
.B(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_72),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_73),
.A2(n_77),
.B1(n_78),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_73),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_328),
.B(n_334),
.Y(n_79)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_300),
.A3(n_321),
.B1(n_326),
.B2(n_327),
.C(n_339),
.Y(n_80)
);

AOI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_253),
.A3(n_275),
.B1(n_293),
.B2(n_299),
.C(n_340),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_212),
.C(n_249),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_183),
.B(n_211),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_156),
.B(n_182),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_136),
.B(n_155),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_124),
.B(n_135),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_110),
.B(n_123),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_98),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_89),
.B(n_98),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_93),
.B(n_153),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_94),
.B(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_96),
.A2(n_116),
.B(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_105),
.B2(n_109),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_109),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_102),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_105),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_118),
.B(n_122),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_116),
.A2(n_117),
.B1(n_168),
.B2(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_116),
.A2(n_152),
.B(n_193),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_116),
.A2(n_117),
.B(n_151),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_117),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_125),
.B(n_126),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_137),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.CI(n_132),
.CON(n_127),
.SN(n_127)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_129),
.A2(n_162),
.B1(n_164),
.B2(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_133),
.B(n_169),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_147),
.B2(n_154),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_140),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_146),
.C(n_154),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_147),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_150),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_157),
.B(n_158),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_174),
.B2(n_175),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_177),
.C(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_173),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_162),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_171),
.C(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_176),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_177),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_178),
.B(n_226),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_185),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_197),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_187),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_196),
.C(n_197),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_207),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_204),
.B2(n_205),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_204),
.C(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_202),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_231),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_213),
.B(n_231),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.C(n_229),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_217),
.C(n_221),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_223),
.B1(n_229),
.B2(n_230),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_228),
.Y(n_234)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_242),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_242),
.C(n_246),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_236),
.C(n_240),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_241),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_244),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_254),
.A2(n_294),
.B(n_298),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_255),
.B(n_256),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_274),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_267),
.B2(n_268),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_268),
.C(n_274),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_262),
.C(n_266),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_264),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_265),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_273),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_270),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_269),
.A2(n_282),
.B(n_285),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_271),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_271),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_276),
.B(n_277),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_277),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_286),
.CI(n_292),
.CON(n_277),
.SN(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_284),
.B2(n_285),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_290),
.B(n_291),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_290),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_289),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_291),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_291),
.A2(n_302),
.B1(n_312),
.B2(n_325),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B(n_297),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_314),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_314),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_312),
.C(n_313),
.Y(n_301)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_304),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_310),
.C(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_316),
.C(n_320),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_307),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_331),
.Y(n_333)
);


endmodule