module real_jpeg_12056_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx10_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_23),
.B1(n_27),
.B2(n_35),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_6),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_23),
.B1(n_27),
.B2(n_33),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_8),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_10),
.B(n_29),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_29),
.B(n_60),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_45),
.C(n_72),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_10),
.A2(n_23),
.B1(n_27),
.B2(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_10),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_10),
.B(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_11),
.A2(n_23),
.B1(n_27),
.B2(n_65),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_12),
.A2(n_23),
.B1(n_27),
.B2(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_12),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_78),
.Y(n_108)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_92),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_84),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_18),
.B(n_84),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_56),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_32),
.B2(n_34),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_21),
.A2(n_22),
.B1(n_32),
.B2(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

INVx5_ASAP7_75t_SL g27 ( 
.A(n_23),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_23),
.A2(n_26),
.B(n_59),
.C(n_61),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_23),
.A2(n_27),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_23),
.B(n_99),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_SL g61 ( 
.A(n_25),
.B(n_27),
.C(n_30),
.Y(n_61)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_43),
.B2(n_55),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B(n_50),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_46),
.B1(n_72),
.B2(n_73),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_46),
.B(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_49),
.A2(n_66),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_49),
.B(n_64),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_51),
.A2(n_52),
.B1(n_106),
.B2(n_114),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_51),
.A2(n_108),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_52),
.B(n_102),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_68),
.B1(n_82),
.B2(n_83),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_67),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_76),
.B(n_79),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_77),
.B1(n_80),
.B2(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_80),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_70),
.A2(n_80),
.B1(n_91),
.B2(n_103),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_102),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.C(n_90),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_132),
.B(n_137),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_120),
.B(n_131),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_109),
.B(n_119),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_104),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_104),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_100),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_115),
.B(n_118),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_117),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_122),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_126),
.C(n_130),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_136),
.Y(n_137)
);


endmodule