module real_jpeg_28486_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_342, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_342;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_22),
.B1(n_23),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_0),
.A2(n_26),
.B1(n_30),
.B2(n_36),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_0),
.A2(n_36),
.B1(n_57),
.B2(n_59),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_0),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_121)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_1),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_1),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_26),
.B1(n_30),
.B2(n_45),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_2),
.A2(n_45),
.B1(n_57),
.B2(n_59),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_3),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_3),
.A2(n_26),
.B1(n_30),
.B2(n_140),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_140),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_3),
.A2(n_57),
.B1(n_59),
.B2(n_140),
.Y(n_252)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_5),
.A2(n_47),
.B1(n_57),
.B2(n_59),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_5),
.A2(n_26),
.B1(n_30),
.B2(n_47),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_6),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_6),
.B(n_25),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_6),
.B(n_30),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_6),
.A2(n_30),
.B(n_212),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_173),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_6),
.A2(n_54),
.B(n_57),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_6),
.B(n_76),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_6),
.A2(n_95),
.B1(n_116),
.B2(n_260),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_8),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_8),
.A2(n_26),
.B1(n_30),
.B2(n_112),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_112),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_8),
.A2(n_57),
.B1(n_59),
.B2(n_112),
.Y(n_247)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_24),
.B1(n_52),
.B2(n_53),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_24),
.B1(n_57),
.B2(n_59),
.Y(n_101)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_12),
.A2(n_22),
.B1(n_23),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_12),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_12),
.A2(n_26),
.B1(n_30),
.B2(n_175),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_175),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_12),
.A2(n_57),
.B1(n_59),
.B2(n_175),
.Y(n_260)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_15),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_83),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_81),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_20),
.A2(n_43),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_21),
.A2(n_32),
.B(n_80),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_25),
.B(n_28),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_28),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g172 ( 
.A(n_22),
.B(n_173),
.CON(n_172),
.SN(n_172)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_25),
.A2(n_32),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_26),
.A2(n_30),
.B1(n_65),
.B2(n_67),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_26),
.A2(n_33),
.B1(n_172),
.B2(n_186),
.Y(n_185)
);

AOI32xp33_ASAP7_75t_L g210 ( 
.A1(n_26),
.A2(n_52),
.A3(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_210)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_28),
.B(n_30),
.Y(n_186)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_31),
.A2(n_44),
.B(n_48),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_32),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_48),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_73),
.C(n_78),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_39),
.A2(n_40),
.B1(n_337),
.B2(n_339),
.Y(n_336)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.C(n_62),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_41),
.A2(n_42),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_43),
.A2(n_48),
.B1(n_111),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_43),
.A2(n_48),
.B1(n_139),
.B2(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_49),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_49),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_49),
.A2(n_62),
.B1(n_309),
.B2(n_323),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_56),
.B(n_60),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_56),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_50),
.A2(n_104),
.B(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_50),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_50),
.A2(n_60),
.B(n_120),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_50),
.A2(n_56),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_50),
.A2(n_146),
.B(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_50),
.A2(n_56),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_50),
.A2(n_56),
.B1(n_219),
.B2(n_237),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_53),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g213 ( 
.A(n_53),
.B(n_65),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_53),
.A2(n_55),
.B(n_173),
.C(n_239),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_56),
.A2(n_103),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_56),
.B(n_173),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_57),
.Y(n_59)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_59),
.B(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_61),
.B(n_122),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_62),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_63),
.A2(n_75),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_64),
.B(n_70),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_64),
.A2(n_71),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_64),
.A2(n_71),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_64),
.A2(n_71),
.B1(n_169),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_64),
.A2(n_71),
.B1(n_198),
.B2(n_216),
.Y(n_215)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_65),
.Y(n_211)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_76),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_77),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_75),
.A2(n_77),
.B(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_75),
.A2(n_136),
.B(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_78),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_334),
.B(n_340),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_304),
.A3(n_326),
.B1(n_332),
.B2(n_333),
.C(n_342),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_158),
.B(n_303),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_141),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_87),
.B(n_141),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_113),
.C(n_124),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_88),
.A2(n_89),
.B1(n_113),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_105),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_107),
.C(n_109),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_102),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_91),
.B(n_102),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_92),
.A2(n_188),
.B(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_93),
.A2(n_101),
.B(n_129),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_93),
.A2(n_99),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_95),
.A2(n_116),
.B1(n_252),
.B2(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_95),
.B(n_173),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_98),
.A2(n_116),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g117 ( 
.A(n_99),
.Y(n_117)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_108),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_113),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_123),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_114),
.A2(n_115),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_119),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_115),
.A2(n_152),
.B(n_155),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_116),
.A2(n_127),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_124),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_135),
.C(n_137),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_125),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_132),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_135),
.A2(n_137),
.B1(n_138),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_135),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_156),
.B2(n_157),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_151),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_144),
.B(n_151),
.C(n_157),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_147),
.B(n_150),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_147),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_149),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_150),
.B(n_306),
.C(n_316),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_150),
.A2(n_306),
.B1(n_307),
.B2(n_331),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_150),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_156),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_297),
.B(n_302),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_202),
.B(n_283),
.C(n_296),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_190),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_161),
.B(n_190),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_176),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_163),
.B(n_164),
.C(n_176),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_171),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_174),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_184),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_178),
.B(n_182),
.C(n_184),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_187),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.C(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_191),
.A2(n_192),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_196),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.C(n_201),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_282),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_275),
.B(n_281),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_230),
.B(n_274),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_221),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_206),
.B(n_221),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.C(n_217),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_207),
.A2(n_208),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_210),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_228),
.C(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_268),
.B(n_273),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_248),
.B(n_267),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_233),
.B(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_235),
.B1(n_238),
.B2(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_247),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_256),
.B(n_266),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_254),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_261),
.B(n_265),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_259),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_285),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_294),
.B2(n_295),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_291),
.C(n_295),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_318),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_318),
.Y(n_333)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_307)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_308),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_311),
.C(n_313),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_313),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_315),
.B1(n_320),
.B2(n_324),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_324),
.C(n_325),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_316),
.A2(n_317),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_325),
.Y(n_318)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_336),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_337),
.Y(n_339)
);


endmodule