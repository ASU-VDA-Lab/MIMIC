module real_aes_8198_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g480 ( .A1(n_0), .A2(n_153), .B(n_481), .C(n_484), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_1), .B(n_475), .Y(n_485) );
INVx1_ASAP7_75t_L g429 ( .A(n_2), .Y(n_429) );
INVx1_ASAP7_75t_L g151 ( .A(n_3), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_4), .B(n_154), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_5), .A2(n_445), .B1(n_731), .B2(n_732), .C1(n_738), .C2(n_739), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_6), .A2(n_470), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_7), .B(n_435), .Y(n_434) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_8), .A2(n_176), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_9), .A2(n_41), .B1(n_141), .B2(n_199), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_10), .A2(n_11), .B1(n_735), .B2(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_10), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_11), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_12), .B(n_176), .Y(n_184) );
AND2x6_ASAP7_75t_L g156 ( .A(n_13), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_14), .A2(n_156), .B(n_461), .C(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_15), .B(n_42), .Y(n_430) );
INVx1_ASAP7_75t_L g135 ( .A(n_16), .Y(n_135) );
INVx1_ASAP7_75t_L g132 ( .A(n_17), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_18), .B(n_137), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_19), .B(n_154), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_20), .B(n_128), .Y(n_186) );
AO32x2_ASAP7_75t_L g237 ( .A1(n_21), .A2(n_127), .A3(n_170), .B1(n_176), .B2(n_238), .Y(n_237) );
OAI22xp5_ASAP7_75t_SL g116 ( .A1(n_22), .A2(n_33), .B1(n_117), .B2(n_118), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_22), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_23), .B(n_141), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_24), .B(n_128), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_25), .A2(n_56), .B1(n_141), .B2(n_199), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g201 ( .A1(n_26), .A2(n_82), .B1(n_137), .B2(n_141), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_27), .B(n_141), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_28), .A2(n_170), .B(n_461), .C(n_492), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_29), .A2(n_170), .B(n_461), .C(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_30), .Y(n_146) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_31), .A2(n_733), .B1(n_734), .B2(n_737), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_31), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_32), .B(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_33), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_33), .A2(n_118), .B1(n_119), .B2(n_120), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_34), .A2(n_470), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_35), .B(n_172), .Y(n_214) );
INVx2_ASAP7_75t_L g139 ( .A(n_36), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_37), .A2(n_467), .B(n_510), .C(n_511), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_38), .B(n_141), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_39), .B(n_172), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_40), .B(n_221), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_43), .B(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_44), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_45), .B(n_154), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_46), .B(n_470), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_47), .A2(n_467), .B(n_510), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_48), .B(n_141), .Y(n_179) );
INVx1_ASAP7_75t_L g482 ( .A(n_49), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_50), .A2(n_90), .B1(n_199), .B2(n_200), .Y(n_198) );
INVx1_ASAP7_75t_L g535 ( .A(n_51), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_52), .B(n_141), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_53), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_54), .B(n_470), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_55), .B(n_149), .Y(n_183) );
AOI22xp33_ASAP7_75t_SL g190 ( .A1(n_57), .A2(n_61), .B1(n_137), .B2(n_141), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_58), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_59), .B(n_141), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_60), .B(n_141), .Y(n_218) );
INVx1_ASAP7_75t_L g157 ( .A(n_62), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_63), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_64), .B(n_475), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_65), .A2(n_143), .B(n_149), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_66), .B(n_141), .Y(n_152) );
INVx1_ASAP7_75t_L g131 ( .A(n_67), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_68), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_69), .B(n_154), .Y(n_513) );
AO32x2_ASAP7_75t_L g196 ( .A1(n_70), .A2(n_170), .A3(n_176), .B1(n_197), .B2(n_202), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_71), .B(n_155), .Y(n_526) );
INVx1_ASAP7_75t_L g166 ( .A(n_72), .Y(n_166) );
INVx1_ASAP7_75t_L g209 ( .A(n_73), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_74), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_75), .B(n_494), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_76), .A2(n_461), .B(n_463), .C(n_467), .Y(n_460) );
AOI222xp33_ASAP7_75t_SL g103 ( .A1(n_77), .A2(n_104), .B1(n_113), .B2(n_436), .C1(n_438), .C2(n_443), .Y(n_103) );
OAI321xp33_ASAP7_75t_L g113 ( .A1(n_77), .A2(n_114), .A3(n_424), .B1(n_431), .B2(n_432), .C(n_434), .Y(n_113) );
INVx1_ASAP7_75t_L g431 ( .A(n_77), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_78), .B(n_137), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_79), .Y(n_544) );
INVx1_ASAP7_75t_L g112 ( .A(n_80), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_81), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_83), .B(n_199), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_84), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_85), .B(n_137), .Y(n_213) );
INVx2_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_87), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_88), .B(n_169), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_89), .B(n_137), .Y(n_180) );
OR2x2_ASAP7_75t_L g426 ( .A(n_91), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g448 ( .A(n_91), .B(n_428), .Y(n_448) );
INVx2_ASAP7_75t_L g452 ( .A(n_91), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_92), .A2(n_102), .B1(n_137), .B2(n_138), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_93), .B(n_470), .Y(n_508) );
INVx1_ASAP7_75t_L g512 ( .A(n_94), .Y(n_512) );
INVxp67_ASAP7_75t_L g547 ( .A(n_95), .Y(n_547) );
XNOR2xp5_ASAP7_75t_L g114 ( .A(n_96), .B(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_97), .B(n_137), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g464 ( .A(n_99), .Y(n_464) );
INVx1_ASAP7_75t_L g522 ( .A(n_100), .Y(n_522) );
AND2x2_ASAP7_75t_L g537 ( .A(n_101), .B(n_172), .Y(n_537) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
CKINVDCx6p67_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_109), .A2(n_110), .B(n_433), .Y(n_437) );
NOR2xp33_ASAP7_75t_SL g440 ( .A(n_109), .B(n_111), .Y(n_440) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_114), .B(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_119), .B1(n_120), .B2(n_423), .Y(n_115) );
INVx1_ASAP7_75t_L g423 ( .A(n_116), .Y(n_423) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR5x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_314), .C(n_372), .D(n_408), .E(n_415), .Y(n_120) );
NAND3xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_260), .C(n_284), .Y(n_121) );
AOI221xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_192), .B1(n_226), .B2(n_231), .C(n_241), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g394 ( .A1(n_123), .A2(n_395), .B(n_397), .Y(n_394) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_173), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_124), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_159), .Y(n_124) );
INVx2_ASAP7_75t_L g230 ( .A(n_125), .Y(n_230) );
AND2x2_ASAP7_75t_L g243 ( .A(n_125), .B(n_175), .Y(n_243) );
AND2x2_ASAP7_75t_L g297 ( .A(n_125), .B(n_174), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_125), .B(n_160), .Y(n_312) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_133), .B(n_158), .Y(n_125) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_126), .A2(n_161), .B(n_171), .Y(n_160) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_127), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_129), .B(n_130), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_147), .B(n_156), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_140), .C(n_143), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_136), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_136), .A2(n_555), .B(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g142 ( .A(n_139), .Y(n_142) );
INVx1_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
INVx3_ASAP7_75t_L g208 ( .A(n_141), .Y(n_208) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_141), .Y(n_466) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g199 ( .A(n_142), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_142), .Y(n_200) );
AND2x6_ASAP7_75t_L g461 ( .A(n_142), .B(n_462), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_143), .A2(n_464), .B(n_465), .C(n_466), .Y(n_463) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_144), .A2(n_212), .B(n_213), .Y(n_211) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g494 ( .A(n_145), .Y(n_494) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
INVx1_ASAP7_75t_L g221 ( .A(n_146), .Y(n_221) );
INVx1_ASAP7_75t_L g462 ( .A(n_146), .Y(n_462) );
AND2x2_ASAP7_75t_L g471 ( .A(n_146), .B(n_150), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B(n_152), .C(n_153), .Y(n_147) );
O2A1O1Ixp5_ASAP7_75t_L g165 ( .A1(n_148), .A2(n_166), .B(n_167), .C(n_168), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_148), .A2(n_493), .B(n_495), .Y(n_492) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_153), .A2(n_182), .B(n_183), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_153), .A2(n_169), .B1(n_189), .B2(n_190), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_153), .A2(n_169), .B1(n_239), .B2(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_154), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_154), .A2(n_179), .B(n_180), .Y(n_178) );
O2A1O1Ixp5_ASAP7_75t_SL g207 ( .A1(n_154), .A2(n_208), .B(n_209), .C(n_210), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_154), .B(n_547), .Y(n_546) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_155), .A2(n_169), .B1(n_198), .B2(n_201), .Y(n_197) );
BUFx3_ASAP7_75t_L g170 ( .A(n_156), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_156), .A2(n_178), .B(n_181), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_156), .A2(n_207), .B(n_211), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_156), .A2(n_217), .B(n_222), .Y(n_216) );
INVx4_ASAP7_75t_SL g468 ( .A(n_156), .Y(n_468) );
AND2x4_ASAP7_75t_L g470 ( .A(n_156), .B(n_471), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_156), .B(n_471), .Y(n_523) );
AND2x2_ASAP7_75t_L g330 ( .A(n_159), .B(n_271), .Y(n_330) );
AND2x2_ASAP7_75t_L g363 ( .A(n_159), .B(n_175), .Y(n_363) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OR2x2_ASAP7_75t_L g270 ( .A(n_160), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g283 ( .A(n_160), .B(n_175), .Y(n_283) );
AND2x2_ASAP7_75t_L g290 ( .A(n_160), .B(n_271), .Y(n_290) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_160), .Y(n_299) );
AND2x2_ASAP7_75t_L g306 ( .A(n_160), .B(n_174), .Y(n_306) );
INVx1_ASAP7_75t_L g337 ( .A(n_160), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_170), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_168), .A2(n_223), .B(n_224), .Y(n_222) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx4_ASAP7_75t_L g483 ( .A(n_169), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g187 ( .A(n_170), .B(n_188), .C(n_191), .Y(n_187) );
INVx2_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_172), .A2(n_206), .B(n_214), .Y(n_205) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_172), .A2(n_216), .B(n_225), .Y(n_215) );
INVx1_ASAP7_75t_L g500 ( .A(n_172), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_172), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_172), .A2(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g313 ( .A(n_173), .Y(n_313) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_185), .Y(n_173) );
INVx2_ASAP7_75t_L g269 ( .A(n_174), .Y(n_269) );
AND2x2_ASAP7_75t_L g291 ( .A(n_174), .B(n_230), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_174), .B(n_337), .Y(n_342) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_175), .B(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g414 ( .A(n_175), .B(n_378), .Y(n_414) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_184), .Y(n_175) );
INVx4_ASAP7_75t_L g191 ( .A(n_176), .Y(n_191) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_176), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_176), .A2(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g228 ( .A(n_185), .Y(n_228) );
INVx3_ASAP7_75t_L g329 ( .A(n_185), .Y(n_329) );
OR2x2_ASAP7_75t_L g359 ( .A(n_185), .B(n_360), .Y(n_359) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_185), .B(n_269), .Y(n_385) );
AND2x4_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
INVx1_ASAP7_75t_L g272 ( .A(n_186), .Y(n_272) );
AO21x1_ASAP7_75t_L g271 ( .A1(n_188), .A2(n_191), .B(n_272), .Y(n_271) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_191), .A2(n_459), .B(n_472), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_191), .B(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g475 ( .A(n_191), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_191), .B(n_516), .Y(n_515) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_191), .A2(n_521), .B(n_528), .Y(n_520) );
AOI33xp33_ASAP7_75t_L g405 ( .A1(n_192), .A2(n_243), .A3(n_257), .B1(n_329), .B2(n_406), .B3(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OR2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
OR2x2_ASAP7_75t_L g258 ( .A(n_194), .B(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_194), .B(n_255), .Y(n_317) );
OR2x2_ASAP7_75t_L g370 ( .A(n_194), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g296 ( .A(n_195), .B(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g321 ( .A(n_195), .B(n_203), .Y(n_321) );
AND2x2_ASAP7_75t_L g388 ( .A(n_195), .B(n_233), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_195), .A2(n_288), .B(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g235 ( .A(n_196), .Y(n_235) );
INVx1_ASAP7_75t_L g248 ( .A(n_196), .Y(n_248) );
AND2x2_ASAP7_75t_L g267 ( .A(n_196), .B(n_237), .Y(n_267) );
AND2x2_ASAP7_75t_L g316 ( .A(n_196), .B(n_236), .Y(n_316) );
INVx2_ASAP7_75t_L g484 ( .A(n_200), .Y(n_484) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_200), .Y(n_514) );
INVx1_ASAP7_75t_L g497 ( .A(n_202), .Y(n_497) );
INVx2_ASAP7_75t_SL g358 ( .A(n_203), .Y(n_358) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_215), .Y(n_203) );
INVx2_ASAP7_75t_L g278 ( .A(n_204), .Y(n_278) );
INVx1_ASAP7_75t_L g409 ( .A(n_204), .Y(n_409) );
AND2x2_ASAP7_75t_L g422 ( .A(n_204), .B(n_303), .Y(n_422) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g249 ( .A(n_205), .Y(n_249) );
OR2x2_ASAP7_75t_L g255 ( .A(n_205), .B(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_205), .Y(n_266) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_215), .Y(n_233) );
AND2x2_ASAP7_75t_L g250 ( .A(n_215), .B(n_236), .Y(n_250) );
INVx1_ASAP7_75t_L g256 ( .A(n_215), .Y(n_256) );
INVx1_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
AND2x2_ASAP7_75t_L g288 ( .A(n_215), .B(n_237), .Y(n_288) );
INVx2_ASAP7_75t_L g304 ( .A(n_215), .Y(n_304) );
AND2x2_ASAP7_75t_L g397 ( .A(n_215), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_215), .B(n_278), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g252 ( .A(n_228), .Y(n_252) );
INVx1_ASAP7_75t_L g281 ( .A(n_228), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_228), .B(n_312), .Y(n_378) );
INVx1_ASAP7_75t_SL g338 ( .A(n_229), .Y(n_338) );
INVx2_ASAP7_75t_L g259 ( .A(n_230), .Y(n_259) );
AND2x2_ASAP7_75t_L g328 ( .A(n_230), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g344 ( .A(n_230), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g406 ( .A(n_232), .Y(n_406) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g261 ( .A(n_234), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g364 ( .A(n_234), .B(n_354), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_234), .A2(n_375), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AND2x2_ASAP7_75t_L g277 ( .A(n_235), .B(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g302 ( .A(n_235), .Y(n_302) );
INVx1_ASAP7_75t_L g326 ( .A(n_235), .Y(n_326) );
OR2x2_ASAP7_75t_L g390 ( .A(n_236), .B(n_249), .Y(n_390) );
NOR2xp67_ASAP7_75t_L g398 ( .A(n_236), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g303 ( .A(n_237), .B(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g310 ( .A(n_237), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_244), .B1(n_251), .B2(n_253), .Y(n_241) );
OR2x2_ASAP7_75t_L g320 ( .A(n_242), .B(n_270), .Y(n_320) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AOI222xp33_ASAP7_75t_L g361 ( .A1(n_243), .A2(n_362), .B1(n_364), .B2(n_365), .C1(n_366), .C2(n_369), .Y(n_361) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_250), .Y(n_245) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g308 ( .A(n_247), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
AND2x2_ASAP7_75t_SL g262 ( .A(n_249), .B(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_249), .Y(n_333) );
AND2x2_ASAP7_75t_L g381 ( .A(n_249), .B(n_250), .Y(n_381) );
INVx1_ASAP7_75t_L g399 ( .A(n_249), .Y(n_399) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g365 ( .A(n_252), .B(n_291), .Y(n_365) );
AND2x2_ASAP7_75t_L g407 ( .A(n_252), .B(n_283), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_254), .B(n_302), .Y(n_389) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_255), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g282 ( .A(n_259), .B(n_283), .Y(n_282) );
INVx3_ASAP7_75t_L g350 ( .A(n_259), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_264), .B(n_268), .C(n_273), .Y(n_260) );
INVxp67_ASAP7_75t_L g274 ( .A(n_261), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_262), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_262), .B(n_309), .Y(n_404) );
BUFx3_ASAP7_75t_L g368 ( .A(n_263), .Y(n_368) );
INVx1_ASAP7_75t_L g275 ( .A(n_264), .Y(n_275) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g294 ( .A(n_266), .B(n_288), .Y(n_294) );
INVx1_ASAP7_75t_SL g334 ( .A(n_267), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx1_ASAP7_75t_L g324 ( .A(n_269), .Y(n_324) );
AND2x2_ASAP7_75t_L g347 ( .A(n_269), .B(n_330), .Y(n_347) );
INVx1_ASAP7_75t_SL g318 ( .A(n_270), .Y(n_318) );
INVx1_ASAP7_75t_L g345 ( .A(n_271), .Y(n_345) );
AOI31xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .A3(n_276), .B(n_279), .Y(n_273) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g366 ( .A(n_277), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g340 ( .A(n_278), .Y(n_340) );
BUFx2_ASAP7_75t_L g354 ( .A(n_278), .Y(n_354) );
AND2x2_ASAP7_75t_L g382 ( .A(n_278), .B(n_303), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_SL g355 ( .A(n_282), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_283), .B(n_350), .Y(n_396) );
AND2x2_ASAP7_75t_L g403 ( .A(n_283), .B(n_329), .Y(n_403) );
AOI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_289), .B(n_292), .C(n_307), .Y(n_284) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_289), .A2(n_316), .B1(n_317), .B2(n_318), .C(n_319), .Y(n_315) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g323 ( .A(n_290), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g360 ( .A(n_291), .Y(n_360) );
OAI32xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_295), .A3(n_298), .B1(n_300), .B2(n_305), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g346 ( .A1(n_294), .A2(n_347), .B(n_348), .C(n_351), .Y(n_346) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
OAI21xp5_ASAP7_75t_SL g410 ( .A1(n_302), .A2(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g371 ( .A(n_303), .Y(n_371) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_309), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g357 ( .A(n_309), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g374 ( .A(n_311), .Y(n_374) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND4xp25_ASAP7_75t_SL g314 ( .A(n_315), .B(n_327), .C(n_346), .D(n_361), .Y(n_314) );
AND2x2_ASAP7_75t_L g353 ( .A(n_316), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g375 ( .A(n_316), .B(n_368), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_318), .B(n_350), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B1(n_322), .B2(n_325), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_320), .A2(n_371), .B1(n_402), .B2(n_404), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_L g408 ( .A1(n_320), .A2(n_409), .B(n_410), .C(n_413), .Y(n_408) );
INVx2_ASAP7_75t_L g379 ( .A(n_321), .Y(n_379) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_323), .A2(n_357), .B1(n_374), .B2(n_375), .C1(n_376), .C2(n_379), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B(n_331), .C(n_335), .Y(n_327) );
INVx1_ASAP7_75t_L g393 ( .A(n_328), .Y(n_393) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g335 ( .A1(n_332), .A2(n_336), .B1(n_339), .B2(n_341), .Y(n_335) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g362 ( .A(n_344), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g420 ( .A(n_347), .Y(n_420) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B1(n_356), .B2(n_359), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_354), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g411 ( .A(n_359), .Y(n_411) );
INVx1_ASAP7_75t_L g392 ( .A(n_363), .Y(n_392) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_365), .Y(n_419) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND5xp2_ASAP7_75t_L g372 ( .A(n_373), .B(n_380), .C(n_394), .D(n_400), .E(n_405), .Y(n_372) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_383), .C(n_386), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI31xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .A3(n_390), .B(n_391), .Y(n_386) );
INVx1_ASAP7_75t_L g412 ( .A(n_388), .Y(n_412) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI222xp33_ASAP7_75t_L g415 ( .A1(n_402), .A2(n_404), .B1(n_416), .B2(n_419), .C1(n_420), .C2(n_421), .Y(n_415) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx2_ASAP7_75t_L g433 ( .A(n_426), .Y(n_433) );
INVx1_ASAP7_75t_SL g442 ( .A(n_426), .Y(n_442) );
NOR2x2_ASAP7_75t_L g738 ( .A(n_427), .B(n_452), .Y(n_738) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g451 ( .A(n_428), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g435 ( .A(n_433), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
NAND2xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_449), .B1(n_450), .B2(n_453), .Y(n_446) );
INVx2_ASAP7_75t_L g740 ( .A(n_447), .Y(n_740) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_449), .A2(n_453), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx2_ASAP7_75t_L g741 ( .A(n_450), .Y(n_741) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR3x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_639), .C(n_688), .Y(n_453) );
NAND5xp2_ASAP7_75t_L g454 ( .A(n_455), .B(n_573), .C(n_602), .D(n_610), .E(n_625), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_501), .B(n_517), .C(n_557), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_486), .Y(n_456) );
AND2x2_ASAP7_75t_L g568 ( .A(n_457), .B(n_565), .Y(n_568) );
AND2x2_ASAP7_75t_L g601 ( .A(n_457), .B(n_487), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_457), .B(n_505), .Y(n_694) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_474), .Y(n_457) );
INVx2_ASAP7_75t_L g504 ( .A(n_458), .Y(n_504) );
BUFx2_ASAP7_75t_L g668 ( .A(n_458), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_469), .Y(n_459) );
INVx5_ASAP7_75t_L g479 ( .A(n_461), .Y(n_479) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_SL g477 ( .A1(n_468), .A2(n_478), .B(n_479), .C(n_480), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_468), .A2(n_479), .B(n_544), .C(n_545), .Y(n_543) );
BUFx2_ASAP7_75t_L g490 ( .A(n_470), .Y(n_490) );
AND2x2_ASAP7_75t_L g486 ( .A(n_474), .B(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g566 ( .A(n_474), .Y(n_566) );
AND2x2_ASAP7_75t_L g652 ( .A(n_474), .B(n_565), .Y(n_652) );
AND2x2_ASAP7_75t_L g707 ( .A(n_474), .B(n_504), .Y(n_707) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_485), .Y(n_474) );
INVx2_ASAP7_75t_L g510 ( .A(n_479), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g624 ( .A(n_486), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_486), .B(n_505), .Y(n_671) );
INVx5_ASAP7_75t_L g565 ( .A(n_487), .Y(n_565) );
AND2x4_ASAP7_75t_L g586 ( .A(n_487), .B(n_566), .Y(n_586) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_487), .Y(n_608) );
AND2x2_ASAP7_75t_L g683 ( .A(n_487), .B(n_668), .Y(n_683) );
AND2x2_ASAP7_75t_L g686 ( .A(n_487), .B(n_506), .Y(n_686) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_498), .Y(n_487) );
AOI21xp5_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_491), .B(n_497), .Y(n_488) );
INVx2_ASAP7_75t_L g496 ( .A(n_494), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_496), .A2(n_512), .B(n_513), .C(n_514), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_496), .A2(n_514), .B(n_535), .C(n_536), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_501), .B(n_566), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_501), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
AND2x2_ASAP7_75t_L g591 ( .A(n_503), .B(n_566), .Y(n_591) );
AND2x2_ASAP7_75t_L g609 ( .A(n_503), .B(n_506), .Y(n_609) );
INVx1_ASAP7_75t_L g629 ( .A(n_503), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_503), .B(n_565), .Y(n_674) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_503), .Y(n_716) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_504), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_505), .B(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_505), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_505), .A2(n_561), .B(n_622), .C(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g628 ( .A(n_505), .B(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g637 ( .A(n_505), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g641 ( .A(n_505), .B(n_565), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_505), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g656 ( .A(n_505), .B(n_566), .Y(n_656) );
AND2x2_ASAP7_75t_L g706 ( .A(n_505), .B(n_707), .Y(n_706) );
INVx5_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g570 ( .A(n_506), .Y(n_570) );
AND2x2_ASAP7_75t_L g611 ( .A(n_506), .B(n_564), .Y(n_611) );
AND2x2_ASAP7_75t_L g623 ( .A(n_506), .B(n_598), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_506), .B(n_652), .Y(n_670) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_515), .Y(n_506) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_538), .Y(n_517) );
INVx1_ASAP7_75t_L g559 ( .A(n_518), .Y(n_559) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
OR2x2_ASAP7_75t_L g561 ( .A(n_519), .B(n_530), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g567 ( .A(n_519), .B(n_568), .C(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_519), .B(n_540), .Y(n_578) );
OR2x2_ASAP7_75t_L g593 ( .A(n_519), .B(n_581), .Y(n_593) );
AND2x2_ASAP7_75t_L g599 ( .A(n_519), .B(n_549), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_519), .B(n_730), .Y(n_729) );
INVx5_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_520), .B(n_540), .Y(n_596) );
AND2x2_ASAP7_75t_L g635 ( .A(n_520), .B(n_550), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_520), .B(n_549), .Y(n_663) );
OR2x2_ASAP7_75t_L g666 ( .A(n_520), .B(n_549), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
INVx5_ASAP7_75t_SL g581 ( .A(n_530), .Y(n_581) );
OR2x2_ASAP7_75t_L g587 ( .A(n_530), .B(n_539), .Y(n_587) );
AND2x2_ASAP7_75t_L g603 ( .A(n_530), .B(n_604), .Y(n_603) );
AOI321xp33_ASAP7_75t_L g610 ( .A1(n_530), .A2(n_611), .A3(n_612), .B1(n_613), .B2(n_619), .C(n_621), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_530), .B(n_538), .Y(n_620) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_530), .Y(n_633) );
OR2x2_ASAP7_75t_L g680 ( .A(n_530), .B(n_578), .Y(n_680) );
AND2x2_ASAP7_75t_L g702 ( .A(n_530), .B(n_599), .Y(n_702) );
AND2x2_ASAP7_75t_L g721 ( .A(n_530), .B(n_540), .Y(n_721) );
OR2x6_ASAP7_75t_L g530 ( .A(n_531), .B(n_537), .Y(n_530) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_549), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_540), .B(n_549), .Y(n_562) );
AND2x2_ASAP7_75t_L g571 ( .A(n_540), .B(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g598 ( .A(n_540), .Y(n_598) );
AND2x2_ASAP7_75t_L g604 ( .A(n_540), .B(n_599), .Y(n_604) );
INVxp67_ASAP7_75t_L g634 ( .A(n_540), .Y(n_634) );
OR2x2_ASAP7_75t_L g676 ( .A(n_540), .B(n_581), .Y(n_676) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_548), .Y(n_540) );
OR2x2_ASAP7_75t_L g558 ( .A(n_549), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_SL g572 ( .A(n_549), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_549), .B(n_561), .Y(n_605) );
AND2x2_ASAP7_75t_L g654 ( .A(n_549), .B(n_598), .Y(n_654) );
AND2x2_ASAP7_75t_L g692 ( .A(n_549), .B(n_581), .Y(n_692) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_550), .B(n_581), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_560), .B(n_563), .C(n_567), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_558), .A2(n_560), .B1(n_685), .B2(n_687), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_560), .A2(n_583), .B1(n_638), .B2(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_SL g712 ( .A(n_561), .Y(n_712) );
INVx1_ASAP7_75t_SL g612 ( .A(n_562), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_564), .B(n_584), .Y(n_614) );
AOI222xp33_ASAP7_75t_L g625 ( .A1(n_564), .A2(n_605), .B1(n_612), .B2(n_626), .C1(n_630), .C2(n_636), .Y(n_625) );
AND2x2_ASAP7_75t_L g715 ( .A(n_564), .B(n_716), .Y(n_715) );
AND2x4_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx2_ASAP7_75t_L g590 ( .A(n_565), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_565), .B(n_585), .Y(n_660) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_565), .Y(n_697) );
AND2x2_ASAP7_75t_L g700 ( .A(n_565), .B(n_609), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_565), .B(n_716), .Y(n_726) );
INVx1_ASAP7_75t_L g617 ( .A(n_566), .Y(n_617) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_566), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_568), .A2(n_709), .B(n_710), .C(n_713), .Y(n_708) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_570), .B(n_632), .C(n_635), .Y(n_631) );
OR2x2_ASAP7_75t_L g659 ( .A(n_570), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_570), .B(n_586), .Y(n_687) );
OR2x2_ASAP7_75t_L g592 ( .A(n_572), .B(n_593), .Y(n_592) );
AOI211xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B(n_582), .C(n_594), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_575), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g681 ( .A(n_576), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_577), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g595 ( .A(n_580), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_581), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g649 ( .A(n_581), .B(n_599), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_581), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_581), .B(n_598), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_587), .B1(n_588), .B2(n_592), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_584), .B(n_656), .Y(n_655) );
BUFx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_586), .B(n_628), .Y(n_627) );
OAI221xp5_ASAP7_75t_SL g650 ( .A1(n_587), .A2(n_651), .B1(n_653), .B2(n_655), .C(n_657), .Y(n_650) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g705 ( .A(n_590), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g718 ( .A(n_590), .B(n_707), .Y(n_718) );
INVx1_ASAP7_75t_L g638 ( .A(n_591), .Y(n_638) );
INVx1_ASAP7_75t_L g709 ( .A(n_592), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_593), .A2(n_676), .B(n_699), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B(n_600), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI21xp5_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_605), .B(n_606), .Y(n_602) );
INVx1_ASAP7_75t_L g642 ( .A(n_603), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_604), .A2(n_690), .B1(n_693), .B2(n_695), .C(n_698), .Y(n_689) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_612), .A2(n_702), .B1(n_703), .B2(n_705), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g678 ( .A(n_614), .Y(n_678) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NOR2xp67_ASAP7_75t_SL g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g682 ( .A(n_618), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g647 ( .A(n_623), .Y(n_647) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_628), .B(n_652), .Y(n_704) );
INVxp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_634), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g720 ( .A(n_635), .B(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g727 ( .A(n_635), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI211xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_642), .B(n_643), .C(n_677), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B(n_650), .C(n_669), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g730 ( .A(n_654), .Y(n_730) );
AND2x2_ASAP7_75t_L g667 ( .A(n_656), .B(n_668), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B1(n_665), .B2(n_667), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
OR2x2_ASAP7_75t_L g675 ( .A(n_663), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g728 ( .A(n_664), .Y(n_728) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI31xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .A3(n_672), .B(n_675), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI211xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B(n_681), .C(n_684), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
CKINVDCx16_ASAP7_75t_R g685 ( .A(n_686), .Y(n_685) );
NAND5xp2_ASAP7_75t_L g688 ( .A(n_689), .B(n_701), .C(n_708), .D(n_722), .E(n_725), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_700), .A2(n_726), .B1(n_727), .B2(n_729), .Y(n_725) );
INVx1_ASAP7_75t_SL g724 ( .A(n_702), .Y(n_724) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI21xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_717), .B(n_719), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
CKINVDCx14_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
endmodule