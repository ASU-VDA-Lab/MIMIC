module real_jpeg_4449_n_32 (n_17, n_8, n_0, n_21, n_2, n_188, n_185, n_29, n_180, n_10, n_31, n_9, n_186, n_12, n_24, n_187, n_6, n_28, n_183, n_179, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_181, n_1, n_26, n_27, n_20, n_19, n_182, n_184, n_30, n_16, n_15, n_13, n_32);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_185;
input n_29;
input n_180;
input n_10;
input n_31;
input n_9;
input n_186;
input n_12;
input n_24;
input n_187;
input n_6;
input n_28;
input n_183;
input n_179;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_181;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_182;
input n_184;
input n_30;
input n_16;
input n_15;
input n_13;

output n_32;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_0),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_1),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_1),
.B(n_68),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_2),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_2),
.B(n_83),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_3),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_4),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_6),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_8),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_9),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_9),
.B(n_133),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_10),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_11),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_11),
.B(n_163),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_12),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_12),
.B(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_14),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_14),
.B(n_64),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_16),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_17),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_18),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_19),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_19),
.B(n_120),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_20),
.B(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_21),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_22),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_22),
.B(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_23),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_23),
.B(n_60),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_24),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_24),
.B(n_143),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_25),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_25),
.B(n_107),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_26),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_27),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_27),
.B(n_160),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_29),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_31),
.B(n_53),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_31),
.A2(n_50),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_174),
.Y(n_32)
);

AO21x1_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_42),
.B(n_172),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_36),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_54),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_38),
.Y(n_145)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B(n_171),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_44),
.B(n_50),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_46),
.B(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_49),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_49),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_50),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B(n_170),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_158),
.B(n_167),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_135),
.B(n_152),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_78),
.B(n_123),
.C(n_132),
.Y(n_57)
);

NOR4xp25_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_67),
.D(n_73),
.Y(n_58)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_89),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_66),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_66),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_67),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_119),
.B(n_122),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_114),
.B(n_118),
.Y(n_79)
);

AO221x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B1(n_111),
.B2(n_112),
.C(n_113),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_121),
.Y(n_120)
);

BUFx8_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_96),
.B(n_110),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_95),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_106),
.B(n_109),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B(n_105),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_104),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_117),
.Y(n_118)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_129),
.C(n_130),
.D(n_131),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.C(n_146),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_146),
.B(n_153),
.C(n_156),
.D(n_157),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_138),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_151),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_179),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_180),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_181),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_182),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_183),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_184),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_185),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_186),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_187),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_188),
.Y(n_121)
);


endmodule