module fake_jpeg_27812_n_290 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp67_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_28),
.Y(n_51)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_58),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_34),
.C(n_33),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_33),
.C(n_32),
.Y(n_99)
);

OR2x2_ASAP7_75t_SL g93 ( 
.A(n_51),
.B(n_17),
.Y(n_93)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

AO22x1_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_19),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_59),
.Y(n_95)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_43),
.Y(n_83)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_23),
.B1(n_20),
.B2(n_34),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_71),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_39),
.B1(n_20),
.B2(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_74),
.B1(n_77),
.B2(n_81),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_23),
.B1(n_20),
.B2(n_36),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_39),
.B1(n_23),
.B2(n_36),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_29),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_93),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_36),
.B1(n_35),
.B2(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_27),
.B1(n_29),
.B2(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_25),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_35),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_100),
.C(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_98),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_37),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_36),
.B1(n_40),
.B2(n_43),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_96),
.B1(n_97),
.B2(n_31),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_21),
.B1(n_33),
.B2(n_32),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_43),
.B1(n_40),
.B2(n_17),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_26),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_37),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_37),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_37),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_112),
.B(n_85),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_24),
.C(n_43),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_110),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_24),
.C(n_30),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_31),
.B(n_28),
.C(n_30),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_78),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_26),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_117),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_15),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_22),
.B(n_31),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_129),
.B(n_124),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_122),
.A2(n_72),
.B1(n_75),
.B2(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_24),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_131),
.A2(n_138),
.B(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_139),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_97),
.B1(n_71),
.B2(n_90),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_137),
.B1(n_114),
.B2(n_122),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_105),
.B1(n_109),
.B2(n_82),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_86),
.B1(n_79),
.B2(n_87),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_142),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_68),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_149),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_107),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_147),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_95),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_22),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_153),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_102),
.B(n_78),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_28),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_155),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_12),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_103),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_108),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_148),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_103),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_131),
.C(n_144),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_169),
.B(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_114),
.B1(n_119),
.B2(n_123),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_174),
.B1(n_180),
.B2(n_183),
.Y(n_205)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_112),
.B(n_121),
.C(n_116),
.D(n_117),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_127),
.B1(n_64),
.B2(n_70),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_105),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_175),
.A2(n_176),
.B(n_184),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_102),
.C(n_78),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_137),
.C(n_147),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_21),
.B1(n_30),
.B2(n_3),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_140),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_1),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_187),
.Y(n_207)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_197),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_167),
.B1(n_179),
.B2(n_188),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_178),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_143),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_202),
.C(n_175),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_141),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_209),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_145),
.B(n_157),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_146),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_150),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_203),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_155),
.C(n_133),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_204),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_156),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_150),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_153),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_177),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_15),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

XNOR2x2_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_1),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_181),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_1),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_205),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_219),
.B1(n_229),
.B2(n_189),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_226),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_222),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_186),
.C(n_184),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_202),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_239),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_213),
.B(n_191),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_234),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_200),
.B(n_213),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_240),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_191),
.B(n_205),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_247),
.B1(n_248),
.B2(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_209),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_222),
.C(n_223),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_189),
.B1(n_181),
.B2(n_196),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_240),
.C(n_247),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_196),
.C(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_254),
.Y(n_262)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_221),
.C(n_218),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_250),
.C(n_257),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_214),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_265),
.B(n_270),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_239),
.Y(n_265)
);

NOR3xp33_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_220),
.C(n_228),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_269),
.Y(n_275)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_274),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_245),
.B(n_260),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_227),
.Y(n_280)
);

OAI321xp33_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_234),
.A3(n_236),
.B1(n_260),
.B2(n_224),
.C(n_256),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_262),
.A2(n_253),
.B(n_233),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_277),
.A2(n_241),
.B(n_261),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_282),
.C(n_272),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_281),
.Y(n_285)
);

NOR2xp67_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_199),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_168),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.C(n_14),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_168),
.C(n_184),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_287),
.B(n_3),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_12),
.C(n_5),
.Y(n_287)
);

OAI21x1_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_5),
.B(n_6),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_5),
.Y(n_290)
);


endmodule