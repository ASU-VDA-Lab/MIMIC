module fake_ibex_299_n_365 (n_85, n_84, n_64, n_3, n_73, n_65, n_95, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_92, n_96, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_365);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_95;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_92;
input n_96;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_365;

wire n_151;
wire n_171;
wire n_103;
wire n_204;
wire n_274;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_124;
wire n_256;
wire n_193;
wire n_108;
wire n_350;
wire n_165;
wire n_255;
wire n_175;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_239;
wire n_134;
wire n_357;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_176;
wire n_216;
wire n_166;
wire n_163;
wire n_114;
wire n_236;
wire n_189;
wire n_280;
wire n_317;
wire n_340;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_170;
wire n_144;
wire n_270;
wire n_346;
wire n_113;
wire n_117;
wire n_265;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_210;
wire n_348;
wire n_220;
wire n_287;
wire n_243;
wire n_228;
wire n_147;
wire n_251;
wire n_244;
wire n_343;
wire n_310;
wire n_323;
wire n_143;
wire n_106;
wire n_224;
wire n_183;
wire n_333;
wire n_110;
wire n_306;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_109;
wire n_127;
wire n_121;
wire n_325;
wire n_301;
wire n_296;
wire n_120;
wire n_168;
wire n_155;
wire n_315;
wire n_122;
wire n_116;
wire n_289;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_215;
wire n_279;
wire n_235;
wire n_136;
wire n_261;
wire n_221;
wire n_355;
wire n_102;
wire n_99;
wire n_269;
wire n_156;
wire n_126;
wire n_356;
wire n_104;
wire n_141;
wire n_222;
wire n_186;
wire n_349;
wire n_295;
wire n_331;
wire n_230;
wire n_185;
wire n_352;
wire n_290;
wire n_174;
wire n_157;
wire n_219;
wire n_246;
wire n_146;
wire n_207;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_139;
wire n_275;
wire n_129;
wire n_98;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_347;
wire n_335;
wire n_263;
wire n_353;
wire n_359;
wire n_262;
wire n_299;
wire n_137;
wire n_338;
wire n_173;
wire n_363;
wire n_180;
wire n_201;
wire n_351;
wire n_257;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_329;
wire n_188;
wire n_200;
wire n_199;
wire n_308;
wire n_135;
wire n_283;
wire n_111;
wire n_322;
wire n_227;
wire n_115;
wire n_248;
wire n_101;
wire n_190;
wire n_138;
wire n_214;
wire n_238;
wire n_332;
wire n_211;
wire n_218;
wire n_314;
wire n_132;
wire n_277;
wire n_337;
wire n_225;
wire n_360;
wire n_272;
wire n_223;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_148;
wire n_342;
wire n_233;
wire n_118;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_178;
wire n_303;
wire n_362;
wire n_162;
wire n_240;
wire n_282;
wire n_266;
wire n_294;
wire n_112;
wire n_284;
wire n_172;
wire n_250;
wire n_313;
wire n_345;
wire n_119;
wire n_361;
wire n_319;
wire n_195;
wire n_212;
wire n_311;
wire n_97;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_302;
wire n_344;
wire n_297;
wire n_252;
wire n_107;
wire n_149;
wire n_254;
wire n_213;
wire n_271;
wire n_241;
wire n_292;
wire n_364;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_160;
wire n_184;
wire n_232;
wire n_281;

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_11),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_33),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_3),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_0),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g107 ( 
.A(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVxp33_ASAP7_75t_SL g112 ( 
.A(n_12),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_16),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_9),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_40),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_13),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_3),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_46),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_38),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_41),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_93),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_94),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_81),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_19),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_67),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_25),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_85),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_7),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_4),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_23),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_31),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_65),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_0),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_14),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_48),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_18),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_49),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_54),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_43),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_6),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_51),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_55),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_57),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_22),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_53),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_15),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_50),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_30),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_20),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_1),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_4),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_80),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_32),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_21),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_70),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_176),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_L g185 ( 
.A(n_100),
.B(n_103),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_134),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_146),
.Y(n_191)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_101),
.B(n_45),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_129),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_172),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_99),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_143),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_112),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_119),
.B(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_98),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_128),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_105),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_140),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_157),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_128),
.B(n_2),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_108),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_169),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_150),
.B(n_2),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_181),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_R g220 ( 
.A(n_110),
.B(n_56),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_170),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_5),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_111),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_139),
.A2(n_158),
.B1(n_154),
.B2(n_164),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_113),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_164),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_139),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_L g229 ( 
.A(n_116),
.B(n_5),
.Y(n_229)
);

NAND2xp33_ASAP7_75t_R g230 ( 
.A(n_117),
.B(n_17),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_118),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_120),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_97),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_121),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_122),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_123),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_124),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_125),
.B(n_29),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_126),
.B(n_35),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_183),
.B(n_144),
.Y(n_243)
);

AO22x2_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_224),
.B1(n_222),
.B2(n_216),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_142),
.B1(n_177),
.B2(n_175),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

AO22x2_ASAP7_75t_L g248 ( 
.A1(n_186),
.A2(n_141),
.B1(n_174),
.B2(n_173),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_136),
.B1(n_107),
.B2(n_180),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_137),
.C(n_166),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_133),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_156),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

AO22x2_ASAP7_75t_L g256 ( 
.A1(n_190),
.A2(n_212),
.B1(n_238),
.B2(n_213),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_194),
.A2(n_167),
.B1(n_165),
.B2(n_163),
.Y(n_258)
);

AO22x2_ASAP7_75t_L g259 ( 
.A1(n_200),
.A2(n_130),
.B1(n_161),
.B2(n_160),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_162),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_204),
.Y(n_261)
);

NAND2x1p5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_153),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_149),
.B1(n_147),
.B2(n_145),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_195),
.B(n_223),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_184),
.A2(n_131),
.B1(n_132),
.B2(n_127),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_201),
.A2(n_132),
.B(n_127),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_223),
.B(n_132),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_206),
.B(n_127),
.Y(n_270)
);

BUFx8_ASAP7_75t_L g271 ( 
.A(n_225),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_36),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_185),
.B(n_39),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_59),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_237),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_77),
.C(n_79),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_198),
.B(n_82),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_196),
.B(n_84),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_192),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_192),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_192),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

AO22x2_ASAP7_75t_L g290 ( 
.A1(n_191),
.A2(n_87),
.B1(n_189),
.B2(n_193),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_255),
.B(n_208),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_279),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_197),
.B(n_209),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_211),
.B(n_215),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_218),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_220),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_274),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_257),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_267),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_243),
.B(n_252),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_247),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_248),
.A2(n_259),
.B1(n_256),
.B2(n_252),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_289),
.B(n_273),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_241),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_274),
.A2(n_270),
.B(n_277),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_260),
.A2(n_280),
.B1(n_249),
.B2(n_259),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_250),
.A2(n_251),
.B(n_276),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_272),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_265),
.B(n_263),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_242),
.B(n_262),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_301),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_304),
.A2(n_248),
.B1(n_244),
.B2(n_290),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_264),
.B(n_281),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_304),
.A2(n_303),
.B1(n_307),
.B2(n_298),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_285),
.B(n_268),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_295),
.A2(n_254),
.B(n_283),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_313),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_295),
.A2(n_246),
.B(n_258),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_278),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_282),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_294),
.A2(n_266),
.B(n_244),
.Y(n_328)
);

BUFx2_ASAP7_75t_R g329 ( 
.A(n_296),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_302),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_326),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_SL g334 ( 
.A1(n_316),
.A2(n_297),
.B(n_294),
.C(n_309),
.Y(n_334)
);

BUFx4f_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_314),
.A2(n_298),
.B(n_308),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_329),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_330),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_331),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_321),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_335),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_315),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_334),
.A2(n_317),
.B(n_318),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_261),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_339),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_315),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_342),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_347),
.B(n_333),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_346),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_349),
.B(n_338),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_350),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_348),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_352),
.A2(n_290),
.B1(n_349),
.B2(n_351),
.Y(n_355)
);

OA21x2_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_345),
.B(n_320),
.Y(n_356)
);

AOI221xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_354),
.B1(n_336),
.B2(n_337),
.C(n_317),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_343),
.B1(n_345),
.B2(n_335),
.Y(n_358)
);

HB1xp67_ASAP7_75t_SL g359 ( 
.A(n_358),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_359),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_360),
.A2(n_336),
.B1(n_319),
.B2(n_324),
.Y(n_361)
);

O2A1O1Ixp33_ASAP7_75t_SL g362 ( 
.A1(n_360),
.A2(n_271),
.B(n_319),
.C(n_292),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_362),
.A2(n_327),
.B1(n_328),
.B2(n_325),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_363),
.A2(n_361),
.B1(n_323),
.B2(n_325),
.Y(n_364)
);

AOI21xp33_ASAP7_75t_L g365 ( 
.A1(n_364),
.A2(n_325),
.B(n_299),
.Y(n_365)
);


endmodule