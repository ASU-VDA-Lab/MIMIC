module fake_jpeg_9665_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_52),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_17),
.B1(n_21),
.B2(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_56),
.B1(n_20),
.B2(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_57),
.Y(n_77)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_37),
.B1(n_35),
.B2(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_41),
.B1(n_57),
.B2(n_59),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_39),
.B(n_38),
.C(n_36),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_82),
.A3(n_83),
.B1(n_79),
.B2(n_72),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_74),
.B1(n_78),
.B2(n_28),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_71),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_81),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_29),
.B1(n_27),
.B2(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_37),
.B1(n_41),
.B2(n_36),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_84),
.B1(n_41),
.B2(n_22),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_27),
.B1(n_31),
.B2(n_30),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_36),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_40),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

OR2x4_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_38),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_38),
.B(n_28),
.C(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_41),
.B1(n_36),
.B2(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_34),
.B1(n_41),
.B2(n_40),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_34),
.B1(n_32),
.B2(n_24),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_88),
.Y(n_103)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_34),
.B1(n_32),
.B2(n_24),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_46),
.Y(n_97)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_94),
.A2(n_77),
.B1(n_75),
.B2(n_63),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_109),
.B1(n_116),
.B2(n_77),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_99),
.B(n_18),
.Y(n_141)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_65),
.B(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_58),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_107),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_32),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_114),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_76),
.B1(n_66),
.B2(n_67),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_84),
.B1(n_63),
.B2(n_75),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_70),
.B1(n_80),
.B2(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_19),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_117),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_19),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_19),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_88),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_34),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_87),
.B(n_90),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_102),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_124),
.C(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_122),
.B(n_123),
.Y(n_178)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_69),
.C(n_81),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_128),
.B(n_132),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_87),
.B(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_131),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_137),
.B1(n_98),
.B2(n_114),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_100),
.B(n_14),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_93),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_14),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_140),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_146),
.B1(n_145),
.B2(n_106),
.Y(n_157)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_147),
.B1(n_103),
.B2(n_115),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_87),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_24),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_63),
.C(n_77),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_34),
.C(n_73),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_75),
.B1(n_70),
.B2(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_115),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_95),
.A2(n_80),
.B1(n_71),
.B2(n_32),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_148),
.A2(n_149),
.B1(n_113),
.B2(n_135),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_24),
.B1(n_16),
.B2(n_26),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_160),
.B1(n_169),
.B2(n_170),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_152),
.A2(n_162),
.B(n_163),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_153),
.B(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_168),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_105),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_172),
.C(n_179),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_158),
.B1(n_182),
.B2(n_171),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_105),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_159),
.B(n_164),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_110),
.B1(n_101),
.B2(n_119),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_161),
.A2(n_167),
.B1(n_181),
.B2(n_34),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_98),
.B(n_112),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_126),
.B(n_104),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_130),
.B1(n_125),
.B2(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_125),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_127),
.A2(n_119),
.B1(n_116),
.B2(n_96),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_176),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_116),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_133),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_116),
.B(n_96),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_34),
.B(n_16),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_115),
.B1(n_16),
.B2(n_26),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_132),
.A2(n_26),
.B1(n_103),
.B2(n_18),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_194),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_141),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_197),
.C(n_207),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_129),
.B(n_136),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_200),
.B(n_204),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_123),
.C(n_122),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_199),
.B(n_205),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_138),
.B1(n_103),
.B2(n_26),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_202),
.B1(n_181),
.B2(n_161),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_18),
.B1(n_34),
.B2(n_88),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_73),
.B(n_34),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_151),
.A2(n_174),
.B(n_164),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_34),
.Y(n_207)
);

OAI22x1_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_0),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_1),
.B(n_2),
.Y(n_236)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_162),
.B1(n_169),
.B2(n_152),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_213),
.A2(n_214),
.B1(n_235),
.B2(n_3),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_159),
.B1(n_173),
.B2(n_155),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_157),
.B1(n_168),
.B2(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_225),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_179),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_230),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_212),
.B1(n_210),
.B2(n_187),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_172),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_232),
.C(n_233),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_188),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_73),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_13),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_207),
.C(n_197),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_205),
.B(n_12),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_209),
.Y(n_249)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_1),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_185),
.C(n_192),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_195),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_256),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_191),
.B(n_193),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_254),
.B1(n_217),
.B2(n_218),
.Y(n_268)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_241),
.A2(n_250),
.B1(n_4),
.B2(n_5),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

OAI221xp5_ASAP7_75t_SL g247 ( 
.A1(n_222),
.A2(n_226),
.B1(n_204),
.B2(n_199),
.C(n_229),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_249),
.C(n_235),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_187),
.B1(n_200),
.B2(n_201),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_237),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_202),
.C(n_2),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_253),
.C(n_234),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_1),
.C(n_2),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_3),
.B(n_4),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_4),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_220),
.B1(n_248),
.B2(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_258),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_267),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_262),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_213),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_265),
.C(n_272),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_229),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_239),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_250),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_230),
.B1(n_219),
.B2(n_221),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_273),
.B1(n_256),
.B2(n_249),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_232),
.C(n_5),
.Y(n_272)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_11),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_251),
.B(n_252),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_280),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_264),
.B(n_267),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_286),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_254),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_6),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_243),
.C(n_253),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_285),
.C(n_272),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_4),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_6),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_294),
.C(n_283),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_259),
.B1(n_265),
.B2(n_8),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_281),
.B1(n_276),
.B2(n_279),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_6),
.C(n_7),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_7),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_6),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_296),
.B(n_298),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_282),
.B(n_284),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_7),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_8),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_304),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_303),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_294),
.B(n_288),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_8),
.B(n_9),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_290),
.B(n_289),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_308),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_291),
.B(n_300),
.Y(n_314)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_307),
.B(n_299),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_313),
.B(n_312),
.C(n_308),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_9),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_11),
.Y(n_319)
);


endmodule