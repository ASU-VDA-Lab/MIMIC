module real_jpeg_14776_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_0),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_61),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_0),
.A2(n_42),
.B1(n_46),
.B2(n_61),
.Y(n_198)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_3),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_4),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_186),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_186),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_4),
.A2(n_42),
.B1(n_46),
.B2(n_186),
.Y(n_273)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_6),
.A2(n_57),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_6),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_6),
.B(n_81),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_6),
.B(n_28),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g251 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_184),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_6),
.A2(n_34),
.B(n_45),
.C(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_6),
.B(n_72),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_6),
.B(n_98),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_6),
.B(n_40),
.Y(n_278)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_6),
.A2(n_28),
.B(n_237),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_7),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_66),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_7),
.A2(n_42),
.B1(n_46),
.B2(n_66),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_9),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_106),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_106),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_9),
.A2(n_42),
.B1(n_46),
.B2(n_106),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_38),
.B1(n_42),
.B2(n_46),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_63),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_12),
.A2(n_42),
.B1(n_46),
.B2(n_63),
.Y(n_162)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_14),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_143),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_143),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_14),
.A2(n_42),
.B1(n_46),
.B2(n_143),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_15),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_171),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_171),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_15),
.A2(n_42),
.B1(n_46),
.B2(n_171),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_16),
.A2(n_36),
.B1(n_57),
.B2(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_16),
.A2(n_36),
.B1(n_42),
.B2(n_46),
.Y(n_134)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_85),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_73),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_73),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_64),
.C(n_67),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_22),
.A2(n_64),
.B1(n_114),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_22),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_50),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_39),
.C(n_51),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_25)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_26),
.A2(n_32),
.B1(n_111),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_26),
.A2(n_32),
.B1(n_140),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_26),
.A2(n_32),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_26),
.A2(n_32),
.B1(n_205),
.B2(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_28),
.A2(n_29),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_28),
.B(n_54),
.Y(n_201)
);

OAI32xp33_ASAP7_75t_L g235 ( 
.A1(n_28),
.A2(n_30),
.A3(n_33),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g200 ( 
.A1(n_29),
.A2(n_55),
.A3(n_57),
.B1(n_183),
.B2(n_201),
.Y(n_200)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_31),
.B(n_34),
.Y(n_238)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_64),
.C(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_39),
.A2(n_50),
.B1(n_68),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_47),
.B(n_49),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_40),
.A2(n_47),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_40),
.A2(n_47),
.B1(n_49),
.B2(n_103),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_40),
.A2(n_47),
.B1(n_102),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_40),
.A2(n_47),
.B1(n_165),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_40),
.A2(n_47),
.B1(n_192),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_40),
.A2(n_47),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_40),
.A2(n_47),
.B1(n_252),
.B2(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_41),
.A2(n_138),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_41),
.A2(n_166),
.B1(n_231),
.B2(n_289),
.Y(n_288)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_42),
.B(n_275),
.Y(n_274)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_44),
.A2(n_46),
.B(n_184),
.Y(n_254)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_47),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_60),
.B2(n_62),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_53),
.B1(n_60),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_52),
.A2(n_53),
.B1(n_65),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_52),
.A2(n_53),
.B1(n_105),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_52),
.A2(n_53),
.B1(n_142),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_52),
.A2(n_53),
.B1(n_181),
.B2(n_185),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_58),
.B(n_184),
.Y(n_183)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_67),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_72),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_70),
.A2(n_72),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_70),
.A2(n_72),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_84),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_79),
.A2(n_81),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_149),
.B(n_319),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_144),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_120),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_90),
.B(n_120),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_107),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_113),
.C(n_118),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B(n_104),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_93),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_95),
.B1(n_104),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_101),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_98),
.B(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_96),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_96),
.A2(n_98),
.B1(n_162),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_96),
.A2(n_98),
.B1(n_198),
.B2(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_96),
.A2(n_98),
.B1(n_209),
.B2(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_96),
.A2(n_98),
.B1(n_240),
.B2(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_96),
.A2(n_98),
.B1(n_184),
.B2(n_273),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_96),
.A2(n_98),
.B1(n_266),
.B2(n_273),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_97),
.A2(n_134),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_97),
.A2(n_160),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_113),
.B1(n_118),
.B2(n_119),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_109),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.C(n_128),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.C(n_141),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_130),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_141),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_144),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_145),
.B(n_146),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_174),
.B(n_318),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_172),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_151),
.B(n_172),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_152),
.B(n_155),
.Y(n_316)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_156),
.B(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_167),
.C(n_169),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_157),
.A2(n_158),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_163),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_167),
.B(n_169),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_313),
.B(n_317),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_223),
.B(n_301),
.C(n_312),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_210),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_177),
.B(n_210),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_195),
.C(n_202),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_178),
.A2(n_179),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_188),
.C(n_194),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_187)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_195),
.B(n_202),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_196),
.B(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.C(n_208),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_203),
.B(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_208),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_212),
.B(n_213),
.C(n_214),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_216),
.B(n_219),
.C(n_222),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_300),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_244),
.B(n_299),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_241),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_226),
.B(n_241),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_227),
.B(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_229),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_234),
.A2(n_235),
.B1(n_239),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_293),
.B(n_298),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_282),
.B(n_292),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_262),
.B(n_281),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_248),
.B(n_255),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_258),
.C(n_260),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_261),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_270),
.B(n_280),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_268),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_276),
.B(n_279),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_284),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_288),
.C(n_290),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_303),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_311),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_309),
.B2(n_310),
.Y(n_304)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_305),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_310),
.C(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);


endmodule