module fake_netlist_1_2710_n_684 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_684);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_684;
wire n_117;
wire n_663;
wire n_513;
wire n_361;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_21), .Y(n_77) );
BUFx8_ASAP7_75t_SL g78 ( .A(n_46), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_67), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_65), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_16), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_75), .Y(n_82) );
BUFx6f_ASAP7_75t_L g83 ( .A(n_36), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_6), .Y(n_84) );
NAND2xp5_ASAP7_75t_L g85 ( .A(n_12), .B(n_49), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_44), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_69), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_13), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_30), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_61), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_43), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_19), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_41), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_23), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_17), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_45), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_71), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_54), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_4), .Y(n_99) );
OR2x2_ASAP7_75t_L g100 ( .A(n_39), .B(n_55), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_6), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_33), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_52), .Y(n_103) );
NOR2xp67_ASAP7_75t_L g104 ( .A(n_10), .B(n_38), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_7), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_18), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_74), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_53), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_66), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_37), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_15), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_28), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_63), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_22), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_8), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_50), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_64), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_42), .Y(n_121) );
INVxp33_ASAP7_75t_L g122 ( .A(n_31), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_11), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_83), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_78), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_109), .B(n_0), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_109), .B(n_0), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_111), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_103), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVxp67_ASAP7_75t_SL g132 ( .A(n_84), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_105), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_106), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_77), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_89), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_89), .A2(n_26), .B(n_73), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_105), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_91), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_83), .B(n_1), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_91), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_108), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_79), .B(n_1), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_95), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_101), .B(n_2), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_95), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_97), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_82), .B(n_3), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_92), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_122), .B(n_3), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_111), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_113), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_101), .B(n_4), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_81), .B(n_5), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_94), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_86), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_94), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_119), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_119), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
AND2x6_ASAP7_75t_L g167 ( .A(n_152), .B(n_120), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_139), .B(n_130), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_128), .B(n_123), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_132), .B(n_118), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
INVx1_ASAP7_75t_SL g172 ( .A(n_156), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_132), .B(n_99), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_157), .Y(n_174) );
XNOR2xp5_ASAP7_75t_L g175 ( .A(n_129), .B(n_123), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_139), .B(n_102), .Y(n_176) );
INVx4_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_130), .B(n_80), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_128), .A2(n_116), .B1(n_88), .B2(n_115), .Y(n_179) );
OAI21xp33_ASAP7_75t_L g180 ( .A1(n_135), .A2(n_93), .B(n_121), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_135), .A2(n_121), .B1(n_120), .B2(n_96), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_152), .B(n_100), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_155), .B(n_86), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_165), .B(n_98), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_157), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_157), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_163), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_165), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_150), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_164), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_138), .B(n_110), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_164), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_138), .B(n_110), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_126), .B(n_117), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_142), .B(n_114), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_155), .B(n_100), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_142), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_134), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_161), .B(n_153), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_153), .B(n_117), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_154), .B(n_107), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_154), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_161), .B(n_112), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_133), .B(n_107), .Y(n_214) );
AND2x6_ASAP7_75t_L g215 ( .A(n_126), .B(n_85), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_145), .B(n_90), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_127), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_127), .B(n_104), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_147), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_133), .B(n_90), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_147), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_125), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_147), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_157), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_146), .A2(n_87), .B1(n_7), .B2(n_8), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_209), .B(n_217), .Y(n_226) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_222), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_209), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_221), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_175), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_209), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_177), .Y(n_233) );
INVx5_ASAP7_75t_L g234 ( .A(n_177), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_177), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_202), .Y(n_236) );
BUFx5_ASAP7_75t_L g237 ( .A(n_184), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_190), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_207), .B(n_158), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_166), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_223), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_187), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_172), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_168), .A2(n_149), .B1(n_159), .B2(n_148), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_168), .B(n_159), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_171), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_218), .B(n_160), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_219), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_183), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_186), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_188), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_219), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_208), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_205), .A2(n_160), .B1(n_148), .B2(n_143), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_186), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_205), .A2(n_149), .B1(n_141), .B2(n_133), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_170), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_190), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_197), .B(n_141), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_167), .A2(n_149), .B1(n_141), .B2(n_133), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_170), .B(n_141), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_193), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_180), .B(n_151), .Y(n_264) );
AOI21xp33_ASAP7_75t_L g265 ( .A1(n_179), .A2(n_140), .B(n_150), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_170), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_218), .B(n_151), .Y(n_267) );
NOR3xp33_ASAP7_75t_SL g268 ( .A(n_176), .B(n_5), .C(n_9), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_173), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_167), .A2(n_151), .B1(n_150), .B2(n_158), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_196), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_173), .B(n_158), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_216), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_215), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_212), .B(n_158), .Y(n_275) );
BUFx3_ASAP7_75t_L g276 ( .A(n_198), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_173), .B(n_158), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_218), .B(n_158), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_199), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_190), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_200), .B(n_151), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_210), .B(n_151), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_201), .B(n_158), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_167), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_194), .B(n_157), .Y(n_285) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_167), .B(n_151), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_214), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_211), .B(n_151), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_190), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_237), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_236), .B(n_176), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_253), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g293 ( .A1(n_227), .A2(n_178), .B1(n_181), .B2(n_225), .C(n_214), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_243), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_234), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_237), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_234), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_228), .Y(n_298) );
INVxp33_ASAP7_75t_SL g299 ( .A(n_242), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_245), .B(n_215), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_257), .A2(n_181), .B1(n_194), .B2(n_220), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_250), .B(n_269), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_229), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_232), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_226), .A2(n_189), .B(n_213), .Y(n_305) );
AND2x4_ASAP7_75t_SL g306 ( .A(n_255), .B(n_178), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_254), .B(n_215), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_265), .A2(n_213), .B(n_203), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_266), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_237), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_261), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_266), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_227), .A2(n_203), .B(n_189), .C(n_136), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_234), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_278), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_278), .Y(n_316) );
BUFx8_ASAP7_75t_SL g317 ( .A(n_231), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_255), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_234), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_237), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_230), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_247), .A2(n_140), .B(n_195), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g323 ( .A1(n_287), .A2(n_124), .B(n_131), .C(n_136), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_241), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_273), .A2(n_167), .B1(n_215), .B2(n_140), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_241), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_276), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_237), .B(n_182), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_261), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_251), .A2(n_150), .B1(n_215), .B2(n_206), .C(n_182), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_281), .A2(n_140), .B(n_206), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_244), .B(n_150), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_261), .A2(n_140), .B1(n_195), .B2(n_204), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_256), .A2(n_124), .B1(n_131), .B2(n_136), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_284), .B(n_9), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_240), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_246), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_237), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_249), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_293), .B(n_244), .Y(n_340) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_325), .A2(n_268), .B(n_288), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_336), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_331), .A2(n_270), .B(n_285), .Y(n_343) );
OAI21xp5_ASAP7_75t_L g344 ( .A1(n_300), .A2(n_260), .B(n_282), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_320), .B(n_233), .Y(n_345) );
INVx8_ASAP7_75t_L g346 ( .A(n_335), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_295), .Y(n_347) );
INVx6_ASAP7_75t_L g348 ( .A(n_295), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_299), .A2(n_272), .B1(n_277), .B2(n_274), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_333), .A2(n_239), .B(n_275), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_322), .A2(n_282), .B(n_268), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_332), .A2(n_239), .B(n_275), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_295), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_337), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_290), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_294), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_290), .Y(n_357) );
OR2x6_ASAP7_75t_L g358 ( .A(n_335), .B(n_277), .Y(n_358) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_320), .B(n_233), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_307), .A2(n_259), .B(n_267), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_323), .A2(n_285), .B(n_283), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_339), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_305), .A2(n_264), .B(n_272), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_334), .A2(n_283), .B(n_174), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_298), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_303), .Y(n_366) );
OAI21x1_ASAP7_75t_L g367 ( .A1(n_328), .A2(n_204), .B(n_174), .Y(n_367) );
OAI21x1_ASAP7_75t_L g368 ( .A1(n_328), .A2(n_192), .B(n_191), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_304), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_296), .Y(n_370) );
OA21x2_ASAP7_75t_L g371 ( .A1(n_343), .A2(n_330), .B(n_264), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_358), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_340), .B(n_291), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g374 ( .A1(n_340), .A2(n_299), .B(n_311), .C(n_301), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_360), .A2(n_338), .B(n_286), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_358), .A2(n_335), .B1(n_311), .B2(n_306), .Y(n_376) );
INVx8_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_342), .B(n_306), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_355), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_356), .Y(n_380) );
OAI211xp5_ASAP7_75t_L g381 ( .A1(n_349), .A2(n_298), .B(n_292), .C(n_329), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_358), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_355), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g384 ( .A1(n_346), .A2(n_313), .B(n_326), .C(n_324), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_346), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_342), .A2(n_292), .B1(n_309), .B2(n_312), .C(n_318), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_354), .B(n_302), .Y(n_387) );
AOI222xp33_ASAP7_75t_L g388 ( .A1(n_354), .A2(n_302), .B1(n_315), .B2(n_316), .C1(n_327), .C2(n_321), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_346), .B(n_302), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g390 ( .A1(n_358), .A2(n_279), .B(n_271), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_362), .A2(n_262), .B1(n_263), .B2(n_248), .C(n_314), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_360), .A2(n_252), .B(n_296), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_346), .A2(n_297), .B1(n_314), .B2(n_317), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_362), .B(n_319), .Y(n_394) );
CKINVDCx6p67_ASAP7_75t_R g395 ( .A(n_358), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_367), .A2(n_310), .B(n_297), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_366), .A2(n_338), .B1(n_310), .B2(n_319), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_379), .B(n_366), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_372), .A2(n_341), .B1(n_351), .B2(n_365), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_380), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_372), .B(n_369), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_382), .B(n_369), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_396), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_379), .B(n_347), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_383), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_383), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_394), .B(n_347), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_387), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_373), .A2(n_341), .B1(n_351), .B2(n_344), .Y(n_410) );
AOI221x1_ASAP7_75t_SL g411 ( .A1(n_378), .A2(n_10), .B1(n_11), .B2(n_12), .C(n_13), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_395), .B(n_341), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_385), .B(n_353), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_396), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_371), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_389), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_386), .B(n_341), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_371), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_395), .B(n_353), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_385), .B(n_347), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_371), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_392), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_385), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_376), .B(n_353), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_385), .B(n_347), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_384), .B(n_370), .Y(n_426) );
AOI211xp5_ASAP7_75t_L g427 ( .A1(n_381), .A2(n_363), .B(n_344), .C(n_319), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
NOR2x1p5_ASAP7_75t_L g429 ( .A(n_389), .B(n_319), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_377), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_390), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_388), .B(n_351), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_405), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_412), .B(n_384), .Y(n_434) );
INVx3_ASAP7_75t_L g435 ( .A(n_403), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_409), .B(n_351), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_429), .A2(n_377), .B1(n_393), .B2(n_374), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_409), .B(n_377), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_398), .B(n_355), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_398), .B(n_357), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_405), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_408), .B(n_377), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_408), .B(n_391), .Y(n_443) );
BUFx3_ASAP7_75t_L g444 ( .A(n_413), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_400), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_430), .B(n_317), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_406), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_414), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_429), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_401), .B(n_357), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_406), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_406), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_418), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_418), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_404), .B(n_357), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_417), .A2(n_308), .B1(n_363), .B2(n_348), .Y(n_459) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_414), .A2(n_375), .B(n_368), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_401), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_418), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_421), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_404), .B(n_370), .Y(n_465) );
OAI321xp33_ASAP7_75t_L g466 ( .A1(n_432), .A2(n_131), .A3(n_137), .B1(n_124), .B2(n_359), .C(n_345), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_430), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_410), .B(n_370), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_427), .B(n_137), .C(n_191), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_421), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_421), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_403), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_411), .A2(n_137), .B1(n_308), .B2(n_192), .C(n_224), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_403), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_402), .B(n_14), .Y(n_475) );
AOI222xp33_ASAP7_75t_L g476 ( .A1(n_416), .A2(n_295), .B1(n_348), .B2(n_16), .C1(n_14), .C2(n_15), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_430), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_403), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_431), .A2(n_224), .B1(n_248), .B2(n_235), .C(n_359), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_402), .Y(n_480) );
AOI32xp33_ASAP7_75t_L g481 ( .A1(n_431), .A2(n_350), .A3(n_364), .B1(n_343), .B2(n_352), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_433), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_433), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_458), .B(n_399), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_467), .Y(n_485) );
AND3x1_ASAP7_75t_L g486 ( .A(n_446), .B(n_423), .C(n_425), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_449), .B(n_423), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_468), .B(n_426), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_468), .B(n_426), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_448), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_434), .B(n_426), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_441), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_453), .B(n_426), .Y(n_494) );
NAND2xp33_ASAP7_75t_L g495 ( .A(n_437), .B(n_419), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_458), .B(n_422), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_461), .B(n_422), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_464), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_480), .B(n_407), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_434), .B(n_403), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_453), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_434), .B(n_403), .Y(n_502) );
AOI22x1_ASAP7_75t_L g503 ( .A1(n_476), .A2(n_419), .B1(n_413), .B2(n_420), .Y(n_503) );
AND3x1_ASAP7_75t_L g504 ( .A(n_445), .B(n_425), .C(n_420), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_434), .B(n_456), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_464), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_435), .Y(n_507) );
NAND3xp33_ASAP7_75t_SL g508 ( .A(n_475), .B(n_424), .C(n_407), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_444), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_456), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_447), .B(n_428), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_447), .B(n_428), .Y(n_512) );
NOR2x1_ASAP7_75t_L g513 ( .A(n_475), .B(n_424), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_477), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_451), .B(n_436), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_451), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_450), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_448), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_439), .B(n_413), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_470), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_452), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_452), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_436), .B(n_428), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_450), .Y(n_525) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_439), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_462), .B(n_413), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_462), .B(n_364), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_462), .B(n_364), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_444), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_440), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_440), .B(n_348), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_463), .B(n_350), .Y(n_533) );
INVx4_ASAP7_75t_L g534 ( .A(n_438), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_448), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_463), .B(n_350), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_444), .Y(n_537) );
INVxp67_ASAP7_75t_SL g538 ( .A(n_463), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_517), .B(n_457), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_485), .Y(n_540) );
AOI21xp33_ASAP7_75t_SL g541 ( .A1(n_503), .A2(n_438), .B(n_442), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_531), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_538), .A2(n_466), .B(n_479), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_526), .B(n_454), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_525), .B(n_457), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_501), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_505), .B(n_465), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_505), .B(n_465), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_514), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_534), .B(n_459), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_501), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_534), .B(n_459), .Y(n_552) );
NAND2x1p5_ASAP7_75t_L g553 ( .A(n_485), .B(n_435), .Y(n_553) );
NOR2x2_ASAP7_75t_L g554 ( .A(n_504), .B(n_455), .Y(n_554) );
NAND2x1_ASAP7_75t_L g555 ( .A(n_534), .B(n_435), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_499), .B(n_455), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_534), .B(n_443), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_504), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_503), .A2(n_473), .B1(n_469), .B2(n_471), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_485), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_497), .B(n_471), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_515), .B(n_454), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_492), .B(n_435), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_510), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_510), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_482), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_482), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_492), .B(n_474), .Y(n_568) );
NOR3xp33_ASAP7_75t_L g569 ( .A(n_495), .B(n_481), .C(n_474), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_497), .B(n_474), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_506), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_515), .B(n_481), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_486), .B(n_472), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_520), .B(n_472), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_496), .B(n_472), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_506), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_483), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_508), .B(n_478), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_527), .B(n_478), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_537), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_527), .B(n_460), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_518), .Y(n_582) );
NAND4xp75_ASAP7_75t_L g583 ( .A(n_486), .B(n_348), .C(n_460), .D(n_25), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_496), .B(n_460), .Y(n_584) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_498), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_483), .B(n_348), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_491), .B(n_368), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_491), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_494), .B(n_368), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g590 ( .A1(n_541), .A2(n_513), .B(n_489), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_549), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_549), .B(n_513), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_572), .B(n_494), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_569), .B(n_487), .C(n_484), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_557), .A2(n_500), .B1(n_502), .B2(n_489), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_557), .A2(n_493), .B1(n_488), .B2(n_521), .C(n_518), .Y(n_596) );
NOR2xp67_ASAP7_75t_L g597 ( .A(n_558), .B(n_507), .Y(n_597) );
NAND2xp33_ASAP7_75t_L g598 ( .A(n_560), .B(n_530), .Y(n_598) );
NAND3xp33_ASAP7_75t_L g599 ( .A(n_569), .B(n_484), .C(n_521), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_542), .B(n_493), .Y(n_600) );
OAI221xp5_ASAP7_75t_SL g601 ( .A1(n_558), .A2(n_488), .B1(n_530), .B2(n_509), .C(n_502), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_546), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_571), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_551), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_539), .B(n_516), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_547), .B(n_516), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_550), .A2(n_500), .B1(n_509), .B2(n_537), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_559), .A2(n_498), .B1(n_537), .B2(n_532), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_544), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_555), .A2(n_522), .B(n_523), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_564), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_565), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_563), .B(n_507), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_552), .A2(n_559), .B1(n_578), .B2(n_540), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_548), .B(n_512), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_576), .A2(n_507), .B1(n_524), .B2(n_522), .C(n_523), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_573), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_554), .Y(n_618) );
OAI22xp33_ASAP7_75t_SL g619 ( .A1(n_553), .A2(n_524), .B1(n_507), .B2(n_490), .Y(n_619) );
NAND4xp75_ASAP7_75t_L g620 ( .A(n_580), .B(n_511), .C(n_512), .D(n_528), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_576), .A2(n_535), .B1(n_490), .B2(n_519), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_562), .B(n_519), .Y(n_622) );
AOI322xp5_ASAP7_75t_L g623 ( .A1(n_571), .A2(n_511), .A3(n_528), .B1(n_529), .B2(n_533), .C1(n_536), .C2(n_519), .Y(n_623) );
OAI211xp5_ASAP7_75t_L g624 ( .A1(n_578), .A2(n_536), .B(n_533), .C(n_529), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_586), .A2(n_535), .B(n_490), .Y(n_625) );
AOI32xp33_ASAP7_75t_L g626 ( .A1(n_618), .A2(n_554), .A3(n_573), .B1(n_585), .B2(n_581), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_617), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_596), .B(n_585), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_613), .B(n_568), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_591), .B(n_556), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_601), .A2(n_583), .B1(n_553), .B2(n_545), .Y(n_631) );
OAI221xp5_ASAP7_75t_SL g632 ( .A1(n_614), .A2(n_584), .B1(n_574), .B2(n_561), .C(n_575), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_598), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_600), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_609), .B(n_579), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_599), .B(n_570), .C(n_588), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_602), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_590), .A2(n_543), .B(n_582), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_608), .A2(n_577), .B1(n_567), .B2(n_566), .C1(n_587), .C2(n_535), .Y(n_639) );
AOI222xp33_ASAP7_75t_L g640 ( .A1(n_594), .A2(n_224), .B1(n_589), .B2(n_543), .C1(n_367), .C2(n_352), .Y(n_640) );
OA22x2_ASAP7_75t_L g641 ( .A1(n_617), .A2(n_367), .B1(n_361), .B2(n_352), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_604), .Y(n_642) );
OAI31xp33_ASAP7_75t_L g643 ( .A1(n_624), .A2(n_359), .A3(n_345), .B(n_27), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_593), .B(n_224), .Y(n_644) );
AO21x1_ASAP7_75t_SL g645 ( .A1(n_607), .A2(n_20), .B(n_24), .Y(n_645) );
XNOR2x1_ASAP7_75t_L g646 ( .A(n_620), .B(n_29), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g647 ( .A1(n_608), .A2(n_345), .B1(n_34), .B2(n_35), .Y(n_647) );
OAI222xp33_ASAP7_75t_L g648 ( .A1(n_595), .A2(n_32), .B1(n_40), .B2(n_47), .C1(n_48), .C2(n_51), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_632), .A2(n_616), .B1(n_592), .B2(n_619), .C(n_603), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_633), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_639), .B(n_623), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_SL g652 ( .A1(n_633), .A2(n_621), .B(n_606), .C(n_605), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_631), .A2(n_597), .B(n_621), .C(n_625), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_639), .B(n_615), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_637), .Y(n_655) );
AOI221x1_ASAP7_75t_SL g656 ( .A1(n_628), .A2(n_625), .B1(n_612), .B2(n_611), .C(n_610), .Y(n_656) );
AOI211x1_ASAP7_75t_L g657 ( .A1(n_638), .A2(n_622), .B(n_57), .C(n_58), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_634), .B(n_361), .Y(n_658) );
OAI21xp33_ASAP7_75t_SL g659 ( .A1(n_626), .A2(n_56), .B(n_60), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_642), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_643), .A2(n_62), .B(n_68), .C(n_70), .Y(n_661) );
XNOR2x1_ASAP7_75t_L g662 ( .A(n_646), .B(n_76), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_655), .Y(n_663) );
NAND2x1_ASAP7_75t_L g664 ( .A(n_660), .B(n_627), .Y(n_664) );
AOI211x1_ASAP7_75t_L g665 ( .A1(n_656), .A2(n_636), .B(n_647), .C(n_648), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_656), .A2(n_630), .B1(n_627), .B2(n_644), .C(n_635), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_651), .A2(n_629), .B1(n_640), .B2(n_641), .C(n_645), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_650), .Y(n_668) );
AOI322xp5_ASAP7_75t_L g669 ( .A1(n_654), .A2(n_238), .A3(n_258), .B1(n_280), .B2(n_289), .C1(n_641), .C2(n_649), .Y(n_669) );
NOR4xp25_ASAP7_75t_L g670 ( .A(n_652), .B(n_238), .C(n_258), .D(n_280), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_668), .B(n_659), .C(n_653), .Y(n_671) );
NAND3xp33_ASAP7_75t_SL g672 ( .A(n_670), .B(n_661), .C(n_657), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_663), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_664), .Y(n_674) );
OR4x1_ASAP7_75t_L g675 ( .A(n_673), .B(n_665), .C(n_669), .D(n_662), .Y(n_675) );
NAND3xp33_ASAP7_75t_SL g676 ( .A(n_671), .B(n_667), .C(n_666), .Y(n_676) );
OAI221xp5_ASAP7_75t_L g677 ( .A1(n_674), .A2(n_658), .B1(n_258), .B2(n_280), .C(n_289), .Y(n_677) );
INVxp67_ASAP7_75t_L g678 ( .A(n_676), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_677), .Y(n_679) );
XNOR2xp5_ASAP7_75t_L g680 ( .A(n_678), .B(n_672), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_680), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_679), .B(n_675), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_682), .A2(n_238), .B1(n_258), .B2(n_280), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_238), .B1(n_289), .B2(n_676), .Y(n_684) );
endmodule