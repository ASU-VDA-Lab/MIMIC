module fake_ibex_1670_n_1510 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_267, n_268, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_266, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_269, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1510);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_267;
input n_268;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_266;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_269;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1510;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1504;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1471;
wire n_1115;
wire n_998;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_291;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1495;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_270;
wire n_1340;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1397;
wire n_1211;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_40),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_110),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_181),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_152),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_183),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_209),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_116),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_167),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_188),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_128),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_224),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_260),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_147),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_238),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_138),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_102),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_132),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_202),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_144),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_36),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_195),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_118),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_166),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_51),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_93),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_149),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_215),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_236),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_134),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_145),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_14),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_43),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_262),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_191),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_7),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_46),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_137),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_124),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_8),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_34),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_66),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_0),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_218),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_139),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_71),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_136),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_204),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_219),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_66),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_81),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_18),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_165),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_17),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_71),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_206),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_229),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_210),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_212),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_190),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_160),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_1),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_196),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_221),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_251),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_95),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_208),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_15),
.B(n_64),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_163),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_177),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_225),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_65),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_75),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_68),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_245),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_41),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_52),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_104),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_100),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_150),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_57),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_243),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_159),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_36),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_200),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_34),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_96),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_194),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_4),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_223),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_228),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_178),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_173),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_222),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_205),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_80),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_84),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_61),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_91),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_161),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_9),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_248),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_89),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_253),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_148),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_211),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_156),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_56),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_131),
.B(n_114),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_92),
.Y(n_387)
);

BUFx5_ASAP7_75t_L g388 ( 
.A(n_143),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_237),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_169),
.Y(n_390)
);

BUFx2_ASAP7_75t_SL g391 ( 
.A(n_35),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_259),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_197),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_151),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_61),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_112),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_220),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_99),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_227),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_23),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_268),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_73),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_43),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_207),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_98),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_6),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_264),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_146),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_256),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_10),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_176),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_98),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_192),
.Y(n_413)
);

BUFx5_ASAP7_75t_L g414 ( 
.A(n_48),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_97),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_257),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_175),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_2),
.Y(n_418)
);

BUFx10_ASAP7_75t_L g419 ( 
.A(n_141),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_91),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_81),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_25),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_20),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_31),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_3),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_55),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_135),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_11),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_7),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_89),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_96),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_203),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_162),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_187),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_154),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_94),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_110),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_254),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_87),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_265),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_129),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_199),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_85),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_29),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_38),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_90),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_249),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_17),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_47),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_95),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_76),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_180),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_115),
.B(n_113),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_69),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_351),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_414),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_355),
.B(n_0),
.Y(n_457)
);

BUFx12f_ASAP7_75t_L g458 ( 
.A(n_274),
.Y(n_458)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_271),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_369),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_274),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_369),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_330),
.B(n_1),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_351),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_358),
.B(n_2),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_358),
.B(n_3),
.Y(n_467)
);

CKINVDCx6p67_ASAP7_75t_R g468 ( 
.A(n_323),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_271),
.Y(n_469)
);

AND2x2_ASAP7_75t_SL g470 ( 
.A(n_409),
.B(n_117),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_388),
.B(n_4),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_363),
.B(n_5),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_293),
.Y(n_473)
);

CKINVDCx11_ASAP7_75t_R g474 ( 
.A(n_316),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

OAI21x1_ASAP7_75t_L g476 ( 
.A1(n_300),
.A2(n_120),
.B(n_119),
.Y(n_476)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_274),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_335),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_429),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_414),
.Y(n_480)
);

BUFx12f_ASAP7_75t_L g481 ( 
.A(n_279),
.Y(n_481)
);

BUFx12f_ASAP7_75t_L g482 ( 
.A(n_279),
.Y(n_482)
);

OA21x2_ASAP7_75t_L g483 ( 
.A1(n_300),
.A2(n_122),
.B(n_121),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_414),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

BUFx8_ASAP7_75t_L g486 ( 
.A(n_414),
.Y(n_486)
);

OAI22x1_ASAP7_75t_SL g487 ( 
.A1(n_316),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_487)
);

CKINVDCx11_ASAP7_75t_R g488 ( 
.A(n_326),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_370),
.B(n_12),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_370),
.B(n_13),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_276),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_361),
.Y(n_492)
);

OAI22x1_ASAP7_75t_SL g493 ( 
.A1(n_326),
.A2(n_18),
.B1(n_14),
.B2(n_16),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_414),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_414),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_361),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_352),
.B(n_16),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_276),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_398),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

INVx6_ASAP7_75t_L g501 ( 
.A(n_279),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_427),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_422),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_388),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_324),
.A2(n_125),
.B(n_123),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_427),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_308),
.B(n_19),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_324),
.A2(n_127),
.B(n_126),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_350),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_416),
.B(n_19),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_388),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_308),
.B(n_20),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_420),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

OAI22x1_ASAP7_75t_L g517 ( 
.A1(n_446),
.A2(n_24),
.B1(n_21),
.B2(n_22),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_420),
.A2(n_27),
.B1(n_24),
.B2(n_26),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_428),
.B(n_26),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_388),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_446),
.Y(n_521)
);

BUFx8_ASAP7_75t_L g522 ( 
.A(n_388),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_331),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_357),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_431),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_525)
);

BUFx8_ASAP7_75t_SL g526 ( 
.A(n_443),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_331),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_359),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_272),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_357),
.B(n_30),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_312),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_359),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_357),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_321),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_273),
.B(n_32),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_294),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_328),
.B(n_130),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_328),
.B(n_33),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_367),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_298),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_367),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_372),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_419),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_372),
.Y(n_544)
);

INVx6_ASAP7_75t_L g545 ( 
.A(n_419),
.Y(n_545)
);

INVxp33_ASAP7_75t_SL g546 ( 
.A(n_338),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_299),
.B(n_33),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_306),
.B(n_37),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_382),
.Y(n_549)
);

BUFx8_ASAP7_75t_L g550 ( 
.A(n_382),
.Y(n_550)
);

NOR2x1_ASAP7_75t_L g551 ( 
.A(n_454),
.B(n_133),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_315),
.B(n_39),
.Y(n_552)
);

OA22x2_ASAP7_75t_SL g553 ( 
.A1(n_283),
.A2(n_319),
.B1(n_320),
.B2(n_310),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_460),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_466),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_486),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_456),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_466),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_456),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_466),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_462),
.B(n_317),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_480),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_480),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_484),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_484),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_494),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_494),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_495),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_495),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_535),
.B(n_270),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_469),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_524),
.B(n_275),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_467),
.Y(n_575)
);

AO21x2_ASAP7_75t_L g576 ( 
.A1(n_471),
.A2(n_278),
.B(n_277),
.Y(n_576)
);

BUFx6f_ASAP7_75t_SL g577 ( 
.A(n_470),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_524),
.B(n_354),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_524),
.B(n_356),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_502),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_502),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_543),
.B(n_281),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_505),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_513),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_513),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_520),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_520),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_543),
.B(n_318),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_477),
.B(n_280),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_503),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_523),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_503),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_523),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_479),
.B(n_468),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_461),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_537),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_537),
.Y(n_598)
);

INVxp33_ASAP7_75t_SL g599 ( 
.A(n_489),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_472),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_533),
.B(n_477),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_486),
.B(n_375),
.C(n_366),
.Y(n_602)
);

AOI21x1_ASAP7_75t_L g603 ( 
.A1(n_471),
.A2(n_452),
.B(n_440),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_533),
.B(n_376),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_533),
.B(n_378),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_477),
.B(n_380),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_531),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_501),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_455),
.Y(n_609)
);

BUFx4f_ASAP7_75t_L g610 ( 
.A(n_535),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_455),
.Y(n_611)
);

NOR2x1p5_ASAP7_75t_L g612 ( 
.A(n_458),
.B(n_325),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_465),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_463),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_537),
.B(n_489),
.Y(n_615)
);

AO21x2_ASAP7_75t_L g616 ( 
.A1(n_476),
.A2(n_284),
.B(n_282),
.Y(n_616)
);

INVxp33_ASAP7_75t_L g617 ( 
.A(n_534),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_527),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_501),
.B(n_285),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_546),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_511),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_507),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_550),
.B(n_286),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_516),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_473),
.B(n_288),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_516),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_516),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_459),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_459),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_459),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_459),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_475),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_522),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_537),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_522),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_474),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_550),
.B(n_287),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_538),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_538),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_538),
.Y(n_641)
);

AOI21x1_ASAP7_75t_L g642 ( 
.A1(n_476),
.A2(n_452),
.B(n_440),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_475),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_522),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_506),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_475),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_475),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_478),
.B(n_291),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_552),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_528),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_532),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_532),
.Y(n_653)
);

INVxp67_ASAP7_75t_R g654 ( 
.A(n_490),
.Y(n_654)
);

BUFx6f_ASAP7_75t_SL g655 ( 
.A(n_537),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_539),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_541),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_541),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_542),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_545),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_506),
.Y(n_661)
);

AND3x2_ASAP7_75t_L g662 ( 
.A(n_508),
.B(n_345),
.C(n_329),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_542),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_544),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_490),
.Y(n_665)
);

CKINVDCx6p67_ASAP7_75t_R g666 ( 
.A(n_458),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_544),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_481),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_549),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_457),
.B(n_327),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_483),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_481),
.B(n_296),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_483),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_483),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_509),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_492),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_482),
.B(n_515),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_485),
.B(n_302),
.Y(n_678)
);

AO21x2_ASAP7_75t_L g679 ( 
.A1(n_547),
.A2(n_548),
.B(n_512),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_508),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_497),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_509),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_457),
.B(n_464),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_509),
.Y(n_684)
);

AO21x2_ASAP7_75t_L g685 ( 
.A1(n_519),
.A2(n_290),
.B(n_289),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_496),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_492),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_514),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_514),
.Y(n_689)
);

INVxp33_ASAP7_75t_SL g690 ( 
.A(n_530),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_530),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_499),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_504),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_688),
.B(n_689),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_679),
.B(n_536),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_597),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_666),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_620),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_572),
.B(n_551),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_679),
.B(n_540),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_679),
.B(n_292),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_595),
.B(n_517),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_554),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_688),
.B(n_491),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_685),
.B(n_295),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_572),
.B(n_303),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_573),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_578),
.B(n_491),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_685),
.B(n_297),
.Y(n_709)
);

OAI221xp5_ASAP7_75t_L g710 ( 
.A1(n_683),
.A2(n_529),
.B1(n_311),
.B2(n_425),
.C(n_374),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_579),
.B(n_498),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_599),
.A2(n_320),
.B1(n_344),
.B2(n_319),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_685),
.B(n_309),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_691),
.B(n_314),
.Y(n_714)
);

INVxp67_ASAP7_75t_SL g715 ( 
.A(n_599),
.Y(n_715)
);

AO221x1_ASAP7_75t_L g716 ( 
.A1(n_621),
.A2(n_553),
.B1(n_518),
.B2(n_517),
.C(n_525),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_554),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_604),
.B(n_510),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_561),
.B(n_499),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_605),
.B(n_607),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_561),
.B(n_500),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_588),
.B(n_500),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_588),
.B(n_500),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_607),
.B(n_521),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_680),
.B(n_304),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_556),
.B(n_634),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_680),
.B(n_305),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_617),
.B(n_301),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_574),
.B(n_313),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_665),
.B(n_322),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_609),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_617),
.B(n_400),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_611),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_570),
.B(n_332),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_595),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_649),
.B(n_606),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_613),
.Y(n_737)
);

BUFx6f_ASAP7_75t_SL g738 ( 
.A(n_677),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_601),
.B(n_333),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_556),
.B(n_337),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_634),
.B(n_636),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_571),
.B(n_334),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_690),
.B(n_347),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_670),
.B(n_589),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_626),
.B(n_343),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_619),
.B(n_348),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_676),
.Y(n_747)
);

INVx8_ASAP7_75t_L g748 ( 
.A(n_572),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_600),
.B(n_336),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_639),
.B(n_339),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_597),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_640),
.B(n_641),
.Y(n_752)
);

AO221x1_ASAP7_75t_L g753 ( 
.A1(n_577),
.A2(n_488),
.B1(n_526),
.B2(n_493),
.C(n_487),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_650),
.B(n_360),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_677),
.B(n_612),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_677),
.B(n_391),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_668),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_577),
.A2(n_346),
.B1(n_371),
.B2(n_344),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_598),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_645),
.B(n_346),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_626),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_687),
.Y(n_762)
);

NOR2xp67_ASAP7_75t_L g763 ( 
.A(n_602),
.B(n_40),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_686),
.Y(n_764)
);

BUFx6f_ASAP7_75t_SL g765 ( 
.A(n_677),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_555),
.B(n_340),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_555),
.B(n_341),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_654),
.A2(n_383),
.B1(n_401),
.B2(n_371),
.Y(n_768)
);

INVx8_ASAP7_75t_L g769 ( 
.A(n_572),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_558),
.B(n_342),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_582),
.B(n_362),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_598),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_678),
.B(n_365),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_681),
.B(n_368),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_610),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_572),
.B(n_558),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_686),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_654),
.B(n_412),
.Y(n_778)
);

INVxp67_ASAP7_75t_SL g779 ( 
.A(n_610),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_693),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_672),
.B(n_438),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_693),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_692),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_598),
.B(n_384),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_560),
.B(n_575),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_560),
.B(n_389),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_575),
.B(n_392),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_598),
.B(n_393),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_608),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_575),
.B(n_399),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_591),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_635),
.B(n_417),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_651),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_635),
.B(n_433),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_635),
.B(n_434),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_635),
.B(n_435),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_644),
.B(n_441),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_644),
.B(n_442),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_662),
.B(n_418),
.C(n_415),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_594),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_644),
.B(n_447),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_652),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_652),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_653),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_586),
.B(n_377),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_653),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_656),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_618),
.B(n_436),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_576),
.B(n_379),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_658),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_644),
.B(n_681),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_576),
.B(n_381),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_660),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_637),
.Y(n_814)
);

BUFx6f_ASAP7_75t_SL g815 ( 
.A(n_660),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_618),
.B(n_439),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_624),
.B(n_390),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_657),
.B(n_445),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_638),
.B(n_394),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_646),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_658),
.Y(n_821)
);

AND2x6_ASAP7_75t_L g822 ( 
.A(n_655),
.B(n_396),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_669),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_616),
.B(n_349),
.Y(n_825)
);

AO221x1_ASAP7_75t_L g826 ( 
.A1(n_646),
.A2(n_661),
.B1(n_637),
.B2(n_449),
.C(n_395),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_663),
.B(n_451),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_564),
.A2(n_567),
.B1(n_581),
.B2(n_580),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_671),
.B(n_397),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_646),
.B(n_404),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_663),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_664),
.B(n_42),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_667),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_564),
.B(n_407),
.Y(n_834)
);

AO221x1_ASAP7_75t_L g835 ( 
.A1(n_646),
.A2(n_307),
.B1(n_449),
.B2(n_395),
.C(n_432),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_581),
.B(n_408),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_671),
.B(n_411),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_673),
.B(n_413),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_655),
.A2(n_345),
.B1(n_364),
.B2(n_353),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_661),
.B(n_673),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_SL g841 ( 
.A(n_655),
.B(n_373),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_761),
.A2(n_385),
.B(n_402),
.C(n_387),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_720),
.B(n_583),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_830),
.A2(n_642),
.B(n_603),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_698),
.B(n_735),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_827),
.B(n_583),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_703),
.B(n_684),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_816),
.B(n_584),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_716),
.A2(n_702),
.B1(n_695),
.B2(n_700),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_707),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_748),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_694),
.B(n_403),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_840),
.A2(n_675),
.B(n_674),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_717),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_710),
.A2(n_406),
.B(n_410),
.C(n_405),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_757),
.Y(n_856)
);

CKINVDCx6p67_ASAP7_75t_R g857 ( 
.A(n_697),
.Y(n_857)
);

CKINVDCx10_ASAP7_75t_R g858 ( 
.A(n_738),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_708),
.B(n_675),
.Y(n_859)
);

AOI21x1_ASAP7_75t_L g860 ( 
.A1(n_695),
.A2(n_642),
.B(n_603),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_825),
.A2(n_684),
.B(n_682),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_701),
.A2(n_837),
.B(n_838),
.C(n_829),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_701),
.A2(n_682),
.B(n_585),
.C(n_587),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_768),
.B(n_423),
.C(n_421),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_715),
.B(n_745),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_785),
.Y(n_866)
);

OAI321xp33_ASAP7_75t_L g867 ( 
.A1(n_705),
.A2(n_437),
.A3(n_448),
.B1(n_424),
.B2(n_426),
.C(n_430),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_704),
.B(n_444),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_764),
.A2(n_587),
.B(n_559),
.C(n_562),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_809),
.A2(n_559),
.B(n_557),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_769),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_812),
.A2(n_562),
.B(n_557),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_776),
.A2(n_661),
.B(n_616),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_818),
.B(n_616),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_752),
.A2(n_565),
.B(n_563),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_777),
.A2(n_568),
.B(n_569),
.C(n_566),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_758),
.B(n_42),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_732),
.Y(n_878)
);

CKINVDCx10_ASAP7_75t_R g879 ( 
.A(n_738),
.Y(n_879)
);

AOI21xp33_ASAP7_75t_L g880 ( 
.A1(n_711),
.A2(n_743),
.B(n_728),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_760),
.B(n_307),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_724),
.B(n_395),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_778),
.A2(n_449),
.B1(n_453),
.B2(n_386),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_760),
.B(n_44),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_744),
.B(n_629),
.Y(n_885)
);

BUFx4f_ASAP7_75t_L g886 ( 
.A(n_756),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_766),
.A2(n_631),
.B(n_630),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_766),
.A2(n_632),
.B(n_631),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_705),
.A2(n_633),
.B(n_632),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_767),
.A2(n_643),
.B(n_633),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_780),
.A2(n_782),
.B(n_718),
.C(n_713),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_824),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_770),
.A2(n_648),
.B(n_647),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_719),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_709),
.A2(n_590),
.B(n_593),
.C(n_592),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_808),
.B(n_45),
.Y(n_896)
);

BUFx12f_ASAP7_75t_L g897 ( 
.A(n_814),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_781),
.B(n_45),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_758),
.B(n_714),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_714),
.B(n_46),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_721),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_722),
.Y(n_902)
);

OR2x6_ASAP7_75t_L g903 ( 
.A(n_756),
.B(n_47),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_820),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_736),
.B(n_48),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_799),
.B(n_49),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_723),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_756),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_775),
.B(n_49),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_779),
.B(n_50),
.Y(n_910)
);

BUFx4f_ASAP7_75t_L g911 ( 
.A(n_755),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_774),
.B(n_50),
.Y(n_912)
);

OAI321xp33_ASAP7_75t_L g913 ( 
.A1(n_713),
.A2(n_628),
.A3(n_627),
.B1(n_625),
.B2(n_623),
.C(n_622),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_731),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_811),
.A2(n_614),
.B(n_596),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_817),
.B(n_51),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_725),
.B(n_53),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_699),
.A2(n_53),
.B(n_54),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_819),
.B(n_54),
.Y(n_919)
);

NAND2x1p5_ASAP7_75t_L g920 ( 
.A(n_789),
.B(n_55),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_727),
.B(n_57),
.Y(n_921)
);

NOR2x1_ASAP7_75t_L g922 ( 
.A(n_755),
.B(n_596),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_733),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_822),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_755),
.B(n_58),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_791),
.A2(n_622),
.B(n_614),
.C(n_60),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_734),
.B(n_58),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_734),
.B(n_59),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_742),
.B(n_59),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_749),
.B(n_62),
.Y(n_930)
);

BUFx8_ASAP7_75t_L g931 ( 
.A(n_765),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_749),
.B(n_62),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_786),
.A2(n_790),
.B(n_787),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_737),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_730),
.Y(n_935)
);

NAND3xp33_ASAP7_75t_SL g936 ( 
.A(n_839),
.B(n_63),
.C(n_64),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_750),
.A2(n_805),
.B(n_834),
.C(n_800),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_828),
.A2(n_142),
.B(n_140),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_754),
.B(n_67),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_831),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_696),
.B(n_72),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_696),
.B(n_74),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_834),
.B(n_76),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_822),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_822),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_805),
.B(n_77),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_726),
.Y(n_947)
);

NOR2x1_ASAP7_75t_L g948 ( 
.A(n_763),
.B(n_78),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_793),
.A2(n_182),
.B(n_263),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_741),
.B(n_79),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_802),
.A2(n_179),
.B(n_255),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_739),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_706),
.A2(n_184),
.B(n_250),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_803),
.A2(n_806),
.B(n_804),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_L g955 ( 
.A(n_740),
.B(n_82),
.C(n_83),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_807),
.A2(n_185),
.B(n_246),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_784),
.A2(n_174),
.B(n_242),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_810),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_813),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_696),
.B(n_84),
.Y(n_960)
);

BUFx4f_ASAP7_75t_L g961 ( 
.A(n_822),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_836),
.Y(n_962)
);

AND2x2_ASAP7_75t_SL g963 ( 
.A(n_765),
.B(n_86),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_788),
.A2(n_186),
.B(n_241),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_792),
.A2(n_172),
.B(n_239),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_821),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_794),
.A2(n_189),
.B(n_235),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_823),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_773),
.B(n_88),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_795),
.A2(n_171),
.B(n_234),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_796),
.A2(n_170),
.B(n_233),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_797),
.A2(n_198),
.B(n_232),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_798),
.A2(n_193),
.B(n_231),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_833),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_801),
.A2(n_168),
.B(n_230),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_826),
.Y(n_976)
);

BUFx4f_ASAP7_75t_L g977 ( 
.A(n_747),
.Y(n_977)
);

INVx5_ASAP7_75t_L g978 ( 
.A(n_903),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_L g979 ( 
.A(n_904),
.B(n_751),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_914),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_860),
.A2(n_832),
.B(n_835),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_861),
.A2(n_841),
.B(n_729),
.Y(n_982)
);

AOI21x1_ASAP7_75t_L g983 ( 
.A1(n_915),
.A2(n_762),
.B(n_783),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_923),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_934),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_861),
.A2(n_746),
.B(n_771),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_874),
.A2(n_772),
.B(n_759),
.Y(n_987)
);

AO31x2_ASAP7_75t_L g988 ( 
.A1(n_862),
.A2(n_895),
.A3(n_863),
.B(n_918),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_865),
.B(n_850),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_962),
.A2(n_815),
.B1(n_772),
.B2(n_759),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_937),
.A2(n_772),
.B(n_815),
.C(n_753),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_L g992 ( 
.A(n_880),
.B(n_936),
.C(n_845),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_844),
.A2(n_201),
.B(n_269),
.Y(n_993)
);

AO21x1_ASAP7_75t_L g994 ( 
.A1(n_938),
.A2(n_164),
.B(n_226),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_851),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_854),
.Y(n_996)
);

INVx1_ASAP7_75t_SL g997 ( 
.A(n_968),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_894),
.B(n_101),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_856),
.B(n_101),
.Y(n_999)
);

OAI21x1_ASAP7_75t_SL g1000 ( 
.A1(n_924),
.A2(n_103),
.B(n_104),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_943),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_881),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_859),
.A2(n_105),
.B(n_107),
.C(n_108),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_903),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_899),
.B(n_878),
.Y(n_1005)
);

AND3x4_ASAP7_75t_L g1006 ( 
.A(n_864),
.B(n_153),
.C(n_155),
.Y(n_1006)
);

AOI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_976),
.A2(n_157),
.B(n_158),
.Y(n_1007)
);

AO31x2_ASAP7_75t_L g1008 ( 
.A1(n_926),
.A2(n_213),
.A3(n_216),
.B(n_217),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_897),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_901),
.B(n_902),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_858),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_886),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_907),
.B(n_868),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_946),
.A2(n_927),
.B1(n_929),
.B2(n_928),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_935),
.B(n_852),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_968),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_843),
.B(n_952),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_939),
.A2(n_917),
.B(n_921),
.C(n_969),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_SL g1019 ( 
.A(n_944),
.B(n_945),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_889),
.A2(n_872),
.B(n_870),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_866),
.B(n_884),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_847),
.A2(n_905),
.B(n_932),
.C(n_930),
.Y(n_1022)
);

OA21x2_ASAP7_75t_L g1023 ( 
.A1(n_913),
.A2(n_951),
.B(n_949),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_886),
.B(n_963),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_848),
.B(n_842),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_871),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_898),
.B(n_900),
.Y(n_1027)
);

AND3x1_ASAP7_75t_SL g1028 ( 
.A(n_879),
.B(n_911),
.C(n_931),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_846),
.B(n_958),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_857),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_877),
.B(n_911),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_871),
.B(n_922),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_949),
.A2(n_956),
.B(n_951),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_954),
.A2(n_875),
.B(n_887),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_892),
.B(n_974),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_869),
.A2(n_876),
.B(n_888),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_890),
.A2(n_893),
.B(n_913),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_974),
.B(n_885),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_882),
.A2(n_953),
.B(n_912),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_SL g1040 ( 
.A1(n_920),
.A2(n_940),
.B(n_855),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_896),
.B(n_966),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_931),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_957),
.A2(n_971),
.B(n_970),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_925),
.B(n_959),
.Y(n_1044)
);

OAI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_916),
.A2(n_919),
.B(n_883),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_920),
.A2(n_961),
.B1(n_910),
.B2(n_909),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_964),
.A2(n_973),
.B(n_972),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_965),
.A2(n_975),
.B(n_967),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_977),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_867),
.B(n_977),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_950),
.B(n_947),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_867),
.A2(n_906),
.B(n_955),
.C(n_948),
.Y(n_1052)
);

OAI21xp33_ASAP7_75t_SL g1053 ( 
.A1(n_941),
.A2(n_942),
.B(n_960),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_851),
.B(n_871),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_865),
.B(n_761),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_865),
.B(n_761),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_861),
.A2(n_873),
.B(n_874),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_864),
.A2(n_716),
.B1(n_577),
.B2(n_690),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_937),
.A2(n_859),
.B(n_891),
.C(n_933),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_914),
.Y(n_1060)
);

NOR2x1_ASAP7_75t_SL g1061 ( 
.A(n_903),
.B(n_924),
.Y(n_1061)
);

AOI221xp5_ASAP7_75t_SL g1062 ( 
.A1(n_937),
.A2(n_862),
.B1(n_891),
.B2(n_849),
.C(n_874),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_865),
.B(n_761),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_858),
.Y(n_1064)
);

AOI21x1_ASAP7_75t_L g1065 ( 
.A1(n_860),
.A2(n_915),
.B(n_642),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_860),
.A2(n_853),
.B(n_873),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_850),
.B(n_707),
.Y(n_1067)
);

AND3x2_ASAP7_75t_L g1068 ( 
.A(n_850),
.B(n_757),
.C(n_620),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_861),
.A2(n_873),
.B(n_874),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_861),
.A2(n_873),
.B(n_874),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_850),
.B(n_908),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_865),
.B(n_761),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_860),
.A2(n_853),
.B(n_873),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_860),
.A2(n_853),
.B(n_873),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_865),
.B(n_761),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_962),
.B(n_849),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_850),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_851),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_962),
.B(n_849),
.Y(n_1079)
);

NAND2x1p5_ASAP7_75t_L g1080 ( 
.A(n_851),
.B(n_871),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_850),
.B(n_908),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_899),
.B(n_735),
.Y(n_1082)
);

OA22x2_ASAP7_75t_L g1083 ( 
.A1(n_903),
.A2(n_712),
.B1(n_758),
.B2(n_716),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_850),
.B(n_908),
.Y(n_1084)
);

NOR2x1p5_ASAP7_75t_L g1085 ( 
.A(n_857),
.B(n_666),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_861),
.A2(n_840),
.B(n_615),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_891),
.A2(n_862),
.A3(n_873),
.B(n_874),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_SL g1088 ( 
.A(n_924),
.B(n_944),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_850),
.Y(n_1089)
);

AOI21x1_ASAP7_75t_L g1090 ( 
.A1(n_860),
.A2(n_915),
.B(n_642),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_865),
.B(n_761),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_861),
.A2(n_873),
.B(n_874),
.Y(n_1092)
);

BUFx8_ASAP7_75t_SL g1093 ( 
.A(n_897),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_850),
.B(n_908),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_865),
.B(n_761),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_891),
.A2(n_962),
.B1(n_862),
.B2(n_700),
.Y(n_1096)
);

AO31x2_ASAP7_75t_L g1097 ( 
.A1(n_891),
.A2(n_862),
.A3(n_873),
.B(n_874),
.Y(n_1097)
);

OR2x6_ASAP7_75t_L g1098 ( 
.A(n_903),
.B(n_748),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_865),
.B(n_761),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_851),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_914),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_861),
.A2(n_840),
.B(n_615),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_899),
.B(n_735),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_850),
.B(n_707),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_850),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_861),
.A2(n_840),
.B(n_615),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_850),
.Y(n_1107)
);

CKINVDCx11_ASAP7_75t_R g1108 ( 
.A(n_897),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_891),
.A2(n_962),
.B1(n_862),
.B2(n_700),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_865),
.B(n_761),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_937),
.A2(n_859),
.B(n_891),
.C(n_933),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_861),
.A2(n_840),
.B(n_615),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_850),
.B(n_908),
.Y(n_1113)
);

AND2x2_ASAP7_75t_SL g1114 ( 
.A(n_886),
.B(n_963),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_903),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_850),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_865),
.B(n_761),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_865),
.B(n_761),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_865),
.B(n_761),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_891),
.A2(n_862),
.A3(n_873),
.B(n_874),
.Y(n_1120)
);

XOR2xp5_ASAP7_75t_L g1121 ( 
.A(n_850),
.B(n_637),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_937),
.A2(n_859),
.B(n_891),
.C(n_933),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_865),
.B(n_761),
.Y(n_1123)
);

AOI221xp5_ASAP7_75t_SL g1124 ( 
.A1(n_937),
.A2(n_862),
.B1(n_891),
.B2(n_849),
.C(n_874),
.Y(n_1124)
);

OA22x2_ASAP7_75t_L g1125 ( 
.A1(n_903),
.A2(n_712),
.B1(n_758),
.B2(n_716),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_899),
.B(n_735),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_861),
.A2(n_840),
.B(n_615),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_865),
.B(n_761),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_861),
.A2(n_873),
.B(n_874),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_865),
.B(n_761),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_914),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_850),
.B(n_707),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_850),
.B(n_908),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_899),
.B(n_735),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_865),
.B(n_761),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_861),
.A2(n_840),
.B(n_615),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_962),
.B(n_849),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_897),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_850),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_914),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_861),
.A2(n_840),
.B(n_615),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_1098),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_SL g1143 ( 
.A1(n_1114),
.A2(n_1115),
.B1(n_978),
.B2(n_1061),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_992),
.A2(n_1125),
.B1(n_1083),
.B2(n_1103),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_997),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1082),
.B(n_1126),
.Y(n_1146)
);

AO21x2_ASAP7_75t_L g1147 ( 
.A1(n_1037),
.A2(n_1069),
.B(n_1057),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_SL g1148 ( 
.A1(n_1115),
.A2(n_1046),
.B(n_994),
.Y(n_1148)
);

OR3x4_ASAP7_75t_SL g1149 ( 
.A(n_1028),
.B(n_1108),
.C(n_1093),
.Y(n_1149)
);

INVx6_ASAP7_75t_L g1150 ( 
.A(n_978),
.Y(n_1150)
);

OA21x2_ASAP7_75t_L g1151 ( 
.A1(n_1066),
.A2(n_1074),
.B(n_1073),
.Y(n_1151)
);

INVx6_ASAP7_75t_L g1152 ( 
.A(n_978),
.Y(n_1152)
);

AO21x2_ASAP7_75t_L g1153 ( 
.A1(n_1057),
.A2(n_1070),
.B(n_1069),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_1098),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1005),
.B(n_1096),
.Y(n_1155)
);

INVx8_ASAP7_75t_L g1156 ( 
.A(n_1098),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1059),
.A2(n_1122),
.B(n_1111),
.Y(n_1157)
);

NAND2x1p5_ASAP7_75t_L g1158 ( 
.A(n_997),
.B(n_1016),
.Y(n_1158)
);

CKINVDCx11_ASAP7_75t_R g1159 ( 
.A(n_1009),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1134),
.A2(n_1025),
.B1(n_1031),
.B2(n_1001),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1096),
.A2(n_1109),
.B(n_1020),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1109),
.B(n_1010),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1022),
.A2(n_1034),
.B(n_1014),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_996),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_1070),
.A2(n_1129),
.B(n_1092),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1012),
.B(n_1085),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1012),
.B(n_995),
.Y(n_1167)
);

OAI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1040),
.A2(n_1058),
.B1(n_1017),
.B2(n_1015),
.C(n_1027),
.Y(n_1168)
);

AO21x2_ASAP7_75t_L g1169 ( 
.A1(n_1092),
.A2(n_1129),
.B(n_1033),
.Y(n_1169)
);

BUFx2_ASAP7_75t_R g1170 ( 
.A(n_1011),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1062),
.B(n_1124),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_1030),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_980),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_SL g1174 ( 
.A1(n_1046),
.A2(n_1000),
.B(n_990),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_984),
.Y(n_1175)
);

NAND2x1p5_ASAP7_75t_L g1176 ( 
.A(n_1026),
.B(n_1078),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1038),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_1020),
.A2(n_981),
.B(n_1036),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1060),
.Y(n_1179)
);

INVxp67_ASAP7_75t_SL g1180 ( 
.A(n_1038),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1055),
.B(n_1056),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1026),
.B(n_1078),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_996),
.Y(n_1183)
);

BUFx8_ASAP7_75t_L g1184 ( 
.A(n_1138),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1063),
.B(n_1095),
.Y(n_1185)
);

BUFx4f_ASAP7_75t_L g1186 ( 
.A(n_1006),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1014),
.A2(n_1036),
.B(n_1086),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1132),
.B(n_1118),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1102),
.A2(n_1112),
.B(n_1106),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1141),
.A2(n_1136),
.B(n_1127),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1042),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_1064),
.Y(n_1193)
);

NOR2x1_ASAP7_75t_R g1194 ( 
.A(n_1024),
.B(n_1089),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1105),
.Y(n_1195)
);

INVx3_ASAP7_75t_SL g1196 ( 
.A(n_1071),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1043),
.A2(n_1048),
.B(n_1047),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1039),
.A2(n_993),
.B(n_987),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1101),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1131),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1140),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_989),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1123),
.B(n_1128),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1091),
.B(n_1099),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_1035),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1001),
.A2(n_1079),
.B1(n_1076),
.B2(n_1137),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_998),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1023),
.A2(n_982),
.B(n_1045),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1035),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1110),
.B(n_1117),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1100),
.B(n_1071),
.Y(n_1211)
);

AO21x1_ASAP7_75t_L g1212 ( 
.A1(n_1007),
.A2(n_1050),
.B(n_1040),
.Y(n_1212)
);

NAND3xp33_ASAP7_75t_L g1213 ( 
.A(n_1018),
.B(n_1052),
.C(n_1003),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1023),
.A2(n_1045),
.B(n_986),
.Y(n_1214)
);

OR2x6_ASAP7_75t_L g1215 ( 
.A(n_1054),
.B(n_1080),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1119),
.B(n_1130),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1054),
.Y(n_1217)
);

AO222x2_ASAP7_75t_SL g1218 ( 
.A1(n_1121),
.A2(n_1081),
.B1(n_1084),
.B2(n_1133),
.C1(n_1113),
.C2(n_1094),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1219)
);

BUFx2_ASAP7_75t_R g1220 ( 
.A(n_1013),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_998),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1135),
.B(n_1021),
.Y(n_1222)
);

BUFx8_ASAP7_75t_SL g1223 ( 
.A(n_1113),
.Y(n_1223)
);

CKINVDCx6p67_ASAP7_75t_R g1224 ( 
.A(n_1133),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1080),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1053),
.A2(n_1002),
.B(n_1041),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1116),
.B(n_1139),
.Y(n_1227)
);

OA21x2_ASAP7_75t_L g1228 ( 
.A1(n_1087),
.A2(n_1120),
.B(n_1097),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1077),
.B(n_1107),
.Y(n_1229)
);

AO21x2_ASAP7_75t_L g1230 ( 
.A1(n_979),
.A2(n_1041),
.B(n_1097),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1032),
.B(n_1029),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1068),
.Y(n_1232)
);

BUFx4_ASAP7_75t_SL g1233 ( 
.A(n_1004),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1049),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1004),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1044),
.B(n_1104),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1067),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_1087),
.A2(n_1051),
.B(n_988),
.Y(n_1238)
);

AO21x1_ASAP7_75t_L g1239 ( 
.A1(n_999),
.A2(n_1088),
.B(n_1019),
.Y(n_1239)
);

AO21x2_ASAP7_75t_L g1240 ( 
.A1(n_988),
.A2(n_991),
.B(n_1008),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1082),
.B(n_899),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_985),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1054),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1065),
.A2(n_1090),
.B(n_983),
.Y(n_1244)
);

NAND2x1p5_ASAP7_75t_L g1245 ( 
.A(n_978),
.B(n_1115),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_997),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_997),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1098),
.B(n_1115),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1065),
.A2(n_1090),
.B(n_983),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1065),
.A2(n_1090),
.B(n_983),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1218),
.A2(n_1186),
.B1(n_1156),
.B2(n_1168),
.Y(n_1252)
);

AO21x1_ASAP7_75t_L g1253 ( 
.A1(n_1163),
.A2(n_1187),
.B(n_1171),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1181),
.B(n_1185),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1151),
.Y(n_1255)
);

CKINVDCx16_ASAP7_75t_R g1256 ( 
.A(n_1149),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1160),
.A2(n_1220),
.B1(n_1186),
.B2(n_1168),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1195),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1173),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1160),
.A2(n_1220),
.B1(n_1144),
.B2(n_1206),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1146),
.A2(n_1241),
.B1(n_1185),
.B2(n_1203),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1175),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1179),
.Y(n_1263)
);

CKINVDCx11_ASAP7_75t_R g1264 ( 
.A(n_1149),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1199),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1200),
.Y(n_1266)
);

INVx6_ASAP7_75t_L g1267 ( 
.A(n_1215),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1215),
.A2(n_1217),
.B1(n_1233),
.B2(n_1224),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1145),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1215),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1217),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1201),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1159),
.Y(n_1273)
);

BUFx2_ASAP7_75t_SL g1274 ( 
.A(n_1142),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1177),
.B(n_1209),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1181),
.B(n_1203),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1225),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1142),
.B(n_1225),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1174),
.A2(n_1148),
.B(n_1212),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1144),
.A2(n_1206),
.B1(n_1241),
.B2(n_1146),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1235),
.A2(n_1155),
.B1(n_1210),
.B2(n_1204),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1243),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1180),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1177),
.B(n_1209),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1208),
.A2(n_1197),
.B(n_1214),
.Y(n_1285)
);

AOI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1163),
.A2(n_1208),
.B(n_1190),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1145),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1205),
.B(n_1180),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1196),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1246),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1142),
.B(n_1249),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1158),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1155),
.A2(n_1210),
.B1(n_1248),
.B2(n_1191),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1205),
.B(n_1242),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1142),
.B(n_1249),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1196),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1223),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1246),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1247),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1247),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1222),
.B(n_1202),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1222),
.B(n_1216),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1188),
.B(n_1231),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1159),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1244),
.A2(n_1251),
.B(n_1250),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1223),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1147),
.Y(n_1307)
);

AO21x1_ASAP7_75t_SL g1308 ( 
.A1(n_1162),
.A2(n_1161),
.B(n_1157),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1236),
.B(n_1229),
.Y(n_1309)
);

INVx4_ASAP7_75t_L g1310 ( 
.A(n_1156),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1236),
.A2(n_1221),
.B1(n_1207),
.B2(n_1237),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1187),
.A2(n_1189),
.B(n_1198),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1227),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1164),
.Y(n_1314)
);

OR2x6_ASAP7_75t_L g1315 ( 
.A(n_1279),
.B(n_1156),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1283),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1308),
.B(n_1238),
.Y(n_1317)
);

INVx4_ASAP7_75t_L g1318 ( 
.A(n_1291),
.Y(n_1318)
);

INVxp67_ASAP7_75t_SL g1319 ( 
.A(n_1288),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1271),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1255),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1308),
.B(n_1153),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1260),
.A2(n_1232),
.B1(n_1213),
.B2(n_1183),
.Y(n_1323)
);

BUFx8_ASAP7_75t_L g1324 ( 
.A(n_1297),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1288),
.B(n_1153),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1253),
.B(n_1165),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1253),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1271),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1269),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1287),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1292),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1307),
.B(n_1165),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1275),
.B(n_1238),
.Y(n_1333)
);

INVxp33_ASAP7_75t_L g1334 ( 
.A(n_1273),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1294),
.B(n_1228),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1257),
.A2(n_1226),
.B1(n_1161),
.B2(n_1143),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1275),
.B(n_1169),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1254),
.B(n_1193),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1286),
.A2(n_1157),
.B(n_1189),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1290),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1298),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1284),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_L g1343 ( 
.A(n_1268),
.B(n_1249),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1280),
.A2(n_1226),
.B1(n_1143),
.B2(n_1154),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1252),
.A2(n_1237),
.B1(n_1230),
.B2(n_1233),
.Y(n_1345)
);

NAND2xp33_ASAP7_75t_R g1346 ( 
.A(n_1271),
.B(n_1166),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1312),
.B(n_1240),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1294),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1344),
.A2(n_1261),
.B1(n_1302),
.B2(n_1281),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1316),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1343),
.A2(n_1293),
.B1(n_1276),
.B2(n_1264),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1319),
.B(n_1299),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1316),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1321),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1325),
.B(n_1240),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1331),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1343),
.A2(n_1311),
.B1(n_1267),
.B2(n_1270),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1320),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1330),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1342),
.B(n_1259),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1325),
.B(n_1178),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1334),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1342),
.B(n_1262),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1325),
.B(n_1178),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1336),
.A2(n_1264),
.B1(n_1309),
.B2(n_1297),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1335),
.B(n_1230),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1348),
.B(n_1263),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1319),
.B(n_1300),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1322),
.B(n_1305),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1346),
.A2(n_1256),
.B1(n_1303),
.B2(n_1301),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1348),
.B(n_1265),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1333),
.B(n_1314),
.Y(n_1372)
);

AND2x4_ASAP7_75t_SL g1373 ( 
.A(n_1318),
.B(n_1291),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1330),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1323),
.A2(n_1258),
.B1(n_1267),
.B2(n_1291),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1331),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1335),
.B(n_1285),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1328),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1328),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1345),
.A2(n_1267),
.B1(n_1295),
.B2(n_1313),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1350),
.B(n_1326),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1351),
.A2(n_1338),
.B1(n_1322),
.B2(n_1315),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1358),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1369),
.B(n_1322),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1372),
.B(n_1337),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1369),
.B(n_1317),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1350),
.B(n_1326),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1377),
.B(n_1326),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1377),
.B(n_1317),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1361),
.B(n_1347),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1354),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1372),
.B(n_1359),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1362),
.B(n_1306),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1353),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1364),
.B(n_1366),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1353),
.B(n_1327),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1366),
.B(n_1339),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1369),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1369),
.B(n_1332),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1355),
.B(n_1339),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1355),
.B(n_1339),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1357),
.A2(n_1315),
.B1(n_1324),
.B2(n_1279),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1388),
.B(n_1339),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1395),
.B(n_1374),
.Y(n_1404)
);

AOI32xp33_ASAP7_75t_L g1405 ( 
.A1(n_1402),
.A2(n_1357),
.A3(n_1373),
.B1(n_1356),
.B2(n_1376),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1391),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1382),
.A2(n_1378),
.B(n_1373),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_SL g1408 ( 
.A(n_1398),
.B(n_1304),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1398),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1388),
.B(n_1389),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1385),
.B(n_1352),
.Y(n_1411)
);

AOI221xp5_ASAP7_75t_L g1412 ( 
.A1(n_1381),
.A2(n_1329),
.B1(n_1349),
.B2(n_1387),
.C(n_1397),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1395),
.B(n_1356),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1385),
.B(n_1352),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1392),
.B(n_1368),
.Y(n_1415)
);

NAND4xp25_ASAP7_75t_L g1416 ( 
.A(n_1393),
.B(n_1365),
.C(n_1370),
.D(n_1380),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1392),
.B(n_1368),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1384),
.B(n_1379),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1395),
.B(n_1337),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1394),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1383),
.B(n_1370),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1388),
.B(n_1327),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1411),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1407),
.A2(n_1421),
.B1(n_1416),
.B2(n_1376),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1403),
.B(n_1397),
.Y(n_1425)
);

NOR2x1_ASAP7_75t_L g1426 ( 
.A(n_1421),
.B(n_1304),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1408),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1414),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1415),
.Y(n_1429)
);

NAND2x1p5_ASAP7_75t_L g1430 ( 
.A(n_1418),
.B(n_1289),
.Y(n_1430)
);

OR2x6_ASAP7_75t_L g1431 ( 
.A(n_1418),
.B(n_1315),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1408),
.Y(n_1432)
);

NAND4xp25_ASAP7_75t_L g1433 ( 
.A(n_1405),
.B(n_1375),
.C(n_1193),
.D(n_1296),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1406),
.Y(n_1434)
);

AOI322xp5_ASAP7_75t_L g1435 ( 
.A1(n_1412),
.A2(n_1410),
.A3(n_1403),
.B1(n_1422),
.B2(n_1404),
.C1(n_1413),
.C2(n_1397),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1410),
.A2(n_1329),
.B(n_1340),
.Y(n_1436)
);

OR2x6_ASAP7_75t_SL g1437 ( 
.A(n_1417),
.B(n_1192),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1420),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1422),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1419),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1418),
.A2(n_1384),
.B1(n_1401),
.B2(n_1400),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1409),
.B(n_1389),
.Y(n_1442)
);

OAI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1427),
.A2(n_1398),
.B1(n_1409),
.B2(n_1318),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1438),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1424),
.A2(n_1409),
.B(n_1373),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1432),
.A2(n_1324),
.B1(n_1398),
.B2(n_1289),
.Y(n_1446)
);

NOR3xp33_ASAP7_75t_L g1447 ( 
.A(n_1424),
.B(n_1273),
.C(n_1172),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1434),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1442),
.B(n_1389),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1439),
.Y(n_1450)
);

OAI221xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1435),
.A2(n_1315),
.B1(n_1400),
.B2(n_1401),
.C(n_1387),
.Y(n_1451)
);

AOI321xp33_ASAP7_75t_L g1452 ( 
.A1(n_1426),
.A2(n_1400),
.A3(n_1401),
.B1(n_1399),
.B2(n_1384),
.C(n_1386),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1437),
.A2(n_1386),
.B1(n_1384),
.B2(n_1318),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1446),
.B(n_1447),
.Y(n_1454)
);

AND2x4_ASAP7_75t_SL g1455 ( 
.A(n_1447),
.B(n_1431),
.Y(n_1455)
);

NAND2x2_ASAP7_75t_L g1456 ( 
.A(n_1446),
.B(n_1170),
.Y(n_1456)
);

AOI21xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1453),
.A2(n_1430),
.B(n_1436),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1448),
.Y(n_1458)
);

OAI322xp33_ASAP7_75t_L g1459 ( 
.A1(n_1443),
.A2(n_1429),
.A3(n_1423),
.B1(n_1428),
.B2(n_1425),
.C1(n_1440),
.C2(n_1430),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1444),
.Y(n_1460)
);

AOI211xp5_ASAP7_75t_L g1461 ( 
.A1(n_1451),
.A2(n_1433),
.B(n_1436),
.C(n_1194),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1450),
.Y(n_1462)
);

OAI211xp5_ASAP7_75t_L g1463 ( 
.A1(n_1452),
.A2(n_1441),
.B(n_1296),
.C(n_1425),
.Y(n_1463)
);

AOI211xp5_ASAP7_75t_L g1464 ( 
.A1(n_1445),
.A2(n_1166),
.B(n_1383),
.C(n_1384),
.Y(n_1464)
);

AOI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1449),
.A2(n_1381),
.B1(n_1340),
.B2(n_1341),
.C(n_1399),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_SL g1466 ( 
.A(n_1447),
.B(n_1245),
.C(n_1192),
.Y(n_1466)
);

NAND3x1_ASAP7_75t_L g1467 ( 
.A(n_1447),
.B(n_1324),
.C(n_1170),
.Y(n_1467)
);

NOR3xp33_ASAP7_75t_L g1468 ( 
.A(n_1466),
.B(n_1454),
.C(n_1457),
.Y(n_1468)
);

NOR2x1_ASAP7_75t_SL g1469 ( 
.A(n_1463),
.B(n_1431),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1467),
.A2(n_1431),
.B1(n_1324),
.B2(n_1386),
.Y(n_1470)
);

NAND4xp25_ASAP7_75t_L g1471 ( 
.A(n_1461),
.B(n_1310),
.C(n_1295),
.D(n_1318),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1465),
.B(n_1390),
.Y(n_1472)
);

NAND3xp33_ASAP7_75t_L g1473 ( 
.A(n_1457),
.B(n_1184),
.C(n_1341),
.Y(n_1473)
);

NOR3xp33_ASAP7_75t_L g1474 ( 
.A(n_1459),
.B(n_1310),
.C(n_1282),
.Y(n_1474)
);

NOR2x1_ASAP7_75t_L g1475 ( 
.A(n_1456),
.B(n_1310),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1460),
.B(n_1390),
.Y(n_1476)
);

NOR3x1_ASAP7_75t_L g1477 ( 
.A(n_1455),
.B(n_1184),
.C(n_1379),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1477),
.B(n_1464),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1476),
.Y(n_1479)
);

NOR2x1_ASAP7_75t_L g1480 ( 
.A(n_1473),
.B(n_1462),
.Y(n_1480)
);

OA22x2_ASAP7_75t_L g1481 ( 
.A1(n_1470),
.A2(n_1458),
.B1(n_1461),
.B2(n_1315),
.Y(n_1481)
);

AOI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1468),
.A2(n_1371),
.B1(n_1367),
.B2(n_1363),
.C(n_1360),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1475),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1471),
.A2(n_1386),
.B1(n_1399),
.B2(n_1315),
.Y(n_1484)
);

NOR3xp33_ASAP7_75t_L g1485 ( 
.A(n_1474),
.B(n_1167),
.C(n_1277),
.Y(n_1485)
);

NOR3xp33_ASAP7_75t_L g1486 ( 
.A(n_1472),
.B(n_1167),
.C(n_1277),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1469),
.B(n_1396),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1482),
.B(n_1486),
.Y(n_1488)
);

NAND3xp33_ASAP7_75t_L g1489 ( 
.A(n_1480),
.B(n_1272),
.C(n_1266),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_L g1490 ( 
.A(n_1478),
.B(n_1274),
.Y(n_1490)
);

NOR3xp33_ASAP7_75t_L g1491 ( 
.A(n_1483),
.B(n_1282),
.C(n_1277),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1481),
.Y(n_1492)
);

OAI222xp33_ASAP7_75t_L g1493 ( 
.A1(n_1487),
.A2(n_1245),
.B1(n_1358),
.B2(n_1378),
.C1(n_1270),
.C2(n_1386),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1479),
.B(n_1396),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1485),
.Y(n_1495)
);

NAND4xp75_ASAP7_75t_L g1496 ( 
.A(n_1490),
.B(n_1484),
.C(n_1239),
.D(n_1152),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1494),
.B(n_1406),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1495),
.Y(n_1498)
);

AOI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1492),
.A2(n_1295),
.B(n_1234),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1488),
.B(n_1489),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1499),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1500),
.Y(n_1502)
);

AND3x1_ASAP7_75t_L g1503 ( 
.A(n_1501),
.B(n_1498),
.C(n_1491),
.Y(n_1503)
);

AOI211xp5_ASAP7_75t_L g1504 ( 
.A1(n_1503),
.A2(n_1502),
.B(n_1493),
.C(n_1497),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1504),
.A2(n_1496),
.B(n_1182),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1505),
.A2(n_1278),
.B(n_1176),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1506),
.B(n_1150),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1507),
.A2(n_1211),
.B(n_1219),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1508),
.A2(n_1219),
.B(n_1211),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1509),
.A2(n_1150),
.B1(n_1152),
.B2(n_1267),
.Y(n_1510)
);


endmodule