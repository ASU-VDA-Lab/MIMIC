module fake_jpeg_235_n_227 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_227);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_0),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_76),
.B1(n_56),
.B2(n_65),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_94),
.B1(n_65),
.B2(n_76),
.Y(n_109)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_60),
.B1(n_56),
.B2(n_71),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_68),
.B(n_58),
.Y(n_97)
);

XNOR2x2_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_63),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_77),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_67),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_108),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_55),
.B(n_64),
.C(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_70),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_60),
.C(n_67),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_74),
.B(n_69),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_110),
.A2(n_57),
.B(n_69),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_83),
.B1(n_80),
.B2(n_82),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_115),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_106),
.B1(n_100),
.B2(n_101),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_70),
.B(n_78),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_89),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_131),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_81),
.B1(n_92),
.B2(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_81),
.B1(n_83),
.B2(n_91),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_71),
.B1(n_53),
.B2(n_72),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_75),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_75),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_87),
.B(n_82),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_144),
.B(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_128),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_158),
.C(n_159),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_0),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_149),
.B(n_152),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_78),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_121),
.Y(n_152)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_72),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_157),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_87),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_134),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_61),
.B(n_2),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_1),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_51),
.C(n_50),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_45),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_130),
.B1(n_137),
.B2(n_132),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_169),
.B1(n_7),
.B2(n_10),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_170),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_2),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_167),
.B(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_171),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_140),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_6),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_44),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_175),
.C(n_158),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_43),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_176),
.B(n_156),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_42),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_160),
.C(n_162),
.Y(n_193)
);

AO22x1_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_155),
.B1(n_140),
.B2(n_144),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_143),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_188),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_153),
.B(n_9),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_41),
.C(n_40),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_39),
.C(n_38),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_175),
.C(n_179),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_193),
.B(n_35),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_196),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_202),
.C(n_177),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_184),
.A2(n_190),
.B1(n_182),
.B2(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_166),
.C(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_10),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_203),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_211),
.B1(n_201),
.B2(n_199),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_177),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_209),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_33),
.C(n_32),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_24),
.C(n_14),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_200),
.B(n_11),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_30),
.B(n_29),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_214),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_204),
.B1(n_208),
.B2(n_202),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.C(n_210),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_217),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_217),
.B1(n_206),
.B2(n_216),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_12),
.B(n_14),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_15),
.C(n_16),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_15),
.A3(n_16),
.B1(n_18),
.B2(n_19),
.C1(n_20),
.C2(n_21),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_18),
.B(n_19),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_20),
.Y(n_227)
);


endmodule