module fake_jpeg_27186_n_163 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_5),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_68),
.Y(n_86)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_66),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_81),
.B(n_0),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_61),
.B(n_58),
.C(n_65),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_69),
.B1(n_59),
.B2(n_55),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_85),
.B1(n_88),
.B2(n_83),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_59),
.B1(n_44),
.B2(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_60),
.C(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_61),
.B1(n_48),
.B2(n_52),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_67),
.B1(n_49),
.B2(n_68),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_67),
.B1(n_53),
.B2(n_62),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_54),
.B1(n_50),
.B2(n_64),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_49),
.B1(n_51),
.B2(n_46),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_46),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_94),
.B1(n_95),
.B2(n_92),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_113),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_112),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_4),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_6),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_7),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_124),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_25),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_123),
.Y(n_129)
);

OR2x6_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_97),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_8),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_126),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_109),
.B1(n_110),
.B2(n_10),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_131),
.B1(n_135),
.B2(n_137),
.Y(n_142)
);

AOI32xp33_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_109),
.A3(n_26),
.B1(n_39),
.B2(n_38),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_110),
.B(n_9),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_14),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_8),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_138),
.B1(n_37),
.B2(n_29),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_122),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_24),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_11),
.C(n_13),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_18),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_140),
.Y(n_143)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_16),
.C(n_17),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_154),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_151),
.C(n_145),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_147),
.B(n_144),
.C(n_152),
.D(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_147),
.Y(n_161)
);

OAI211xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_129),
.B(n_149),
.C(n_141),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_146),
.Y(n_163)
);


endmodule