module fake_netlist_1_6792_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
BUFx6f_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_1), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_14), .B(n_0), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_5), .B(n_6), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_15), .B(n_0), .C(n_2), .Y(n_20) );
OR2x6_ASAP7_75t_L g21 ( .A(n_12), .B(n_2), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_16), .A2(n_7), .B(n_3), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_18), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
BUFx3_ASAP7_75t_L g26 ( .A(n_21), .Y(n_26) );
NOR2xp33_ASAP7_75t_L g27 ( .A(n_24), .B(n_13), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_24), .B(n_20), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
NAND2x1p5_ASAP7_75t_L g30 ( .A(n_28), .B(n_26), .Y(n_30) );
AOI211xp5_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_25), .B(n_29), .C(n_27), .Y(n_31) );
A2O1A1Ixp33_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_23), .B(n_19), .C(n_11), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_30), .B(n_17), .Y(n_33) );
CKINVDCx5p33_ASAP7_75t_R g34 ( .A(n_33), .Y(n_34) );
INVxp33_ASAP7_75t_SL g35 ( .A(n_32), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_33), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_23), .B1(n_11), .B2(n_4), .Y(n_37) );
XNOR2xp5_ASAP7_75t_L g38 ( .A(n_36), .B(n_11), .Y(n_38) );
AOI22xp33_ASAP7_75t_L g39 ( .A1(n_37), .A2(n_11), .B1(n_35), .B2(n_38), .Y(n_39) );
endmodule