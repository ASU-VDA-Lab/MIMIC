module fake_jpeg_19043_n_142 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_1),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_6),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_26),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_22),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_48),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_18),
.B1(n_19),
.B2(n_29),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_31),
.B(n_25),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_40),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_63),
.B(n_70),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_39),
.B1(n_23),
.B2(n_29),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_68),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_35),
.B1(n_41),
.B2(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_78),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_22),
.B(n_20),
.C(n_16),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_58),
.A3(n_43),
.B1(n_42),
.B2(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_9),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_49),
.C(n_48),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_85),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_76),
.Y(n_99)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

CKINVDCx11_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_60),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_57),
.C(n_52),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_78),
.Y(n_101)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_104),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_74),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_101),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_96),
.B(n_86),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_75),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_76),
.B1(n_60),
.B2(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_107),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_87),
.B(n_84),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_92),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_71),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_35),
.Y(n_118)
);

AOI331xp33_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_66),
.A3(n_65),
.B1(n_61),
.B2(n_79),
.B3(n_69),
.C1(n_41),
.Y(n_109)
);

OAI321xp33_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_81),
.A3(n_35),
.B1(n_54),
.B2(n_90),
.C(n_28),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_95),
.B(n_84),
.C(n_96),
.D(n_89),
.Y(n_110)
);

NOR4xp25_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_118),
.C(n_109),
.D(n_98),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_89),
.B(n_86),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_125),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_124),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_100),
.C(n_104),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_54),
.C(n_28),
.Y(n_131)
);

NOR2xp67_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_129),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_111),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_131),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_112),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_120),
.B(n_7),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_130),
.B(n_3),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_54),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_137),
.B(n_138),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_132),
.B1(n_128),
.B2(n_4),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_54),
.C(n_3),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_139),
.Y(n_142)
);


endmodule