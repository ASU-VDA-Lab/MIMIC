module fake_jpeg_4869_n_330 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_37),
.B(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_42),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_17),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_14),
.B(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_49),
.B(n_11),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_16),
.B1(n_14),
.B2(n_20),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_55),
.A2(n_65),
.B1(n_91),
.B2(n_92),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_71),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_16),
.B1(n_29),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_57),
.A2(n_101),
.B1(n_102),
.B2(n_71),
.Y(n_118)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_61),
.Y(n_110)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_16),
.B1(n_34),
.B2(n_25),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_63),
.A2(n_79),
.B1(n_96),
.B2(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_15),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_31),
.B1(n_29),
.B2(n_24),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_15),
.Y(n_72)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_17),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_78),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_42),
.A2(n_34),
.B1(n_24),
.B2(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_42),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_81),
.Y(n_112)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_35),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_36),
.B(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_36),
.B(n_35),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_85),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_35),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_40),
.B(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_40),
.B(n_30),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_37),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_37),
.B(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_95),
.Y(n_107)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_44),
.A2(n_32),
.B1(n_22),
.B2(n_33),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_100),
.B1(n_23),
.B2(n_22),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_44),
.A2(n_22),
.B1(n_33),
.B2(n_23),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_44),
.A2(n_23),
.B1(n_22),
.B2(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_22),
.B1(n_23),
.B2(n_33),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_106),
.A2(n_118),
.B1(n_129),
.B2(n_61),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_75),
.C(n_89),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_116),
.C(n_74),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_113),
.A2(n_88),
.B1(n_53),
.B2(n_80),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_21),
.C(n_33),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_60),
.B(n_54),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_126),
.B(n_69),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_58),
.A2(n_21),
.B(n_35),
.Y(n_126)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_136),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_56),
.Y(n_135)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_137),
.B(n_139),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_54),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_138),
.A2(n_156),
.B(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_140),
.A2(n_115),
.B1(n_13),
.B2(n_12),
.Y(n_210)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_141),
.B(n_142),
.Y(n_197)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_124),
.B(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_76),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_144),
.B(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_149),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_163),
.B(n_133),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_62),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_154),
.C(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_52),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_155),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_96),
.B1(n_94),
.B2(n_59),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_167),
.B1(n_130),
.B2(n_108),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_56),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_82),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_18),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_107),
.B(n_70),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_157),
.B(n_161),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_104),
.B(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_53),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_66),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_73),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_119),
.B(n_93),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_93),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_88),
.B1(n_80),
.B2(n_81),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_115),
.B1(n_21),
.B2(n_18),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_105),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_105),
.B(n_81),
.C(n_18),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_128),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_172),
.A2(n_195),
.B(n_203),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_177),
.B1(n_188),
.B2(n_194),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_154),
.B(n_128),
.CI(n_127),
.CON(n_176),
.SN(n_176)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_139),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_149),
.B1(n_162),
.B2(n_166),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_190),
.B(n_201),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_114),
.B1(n_103),
.B2(n_120),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_200),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_114),
.B1(n_103),
.B2(n_120),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_143),
.A2(n_21),
.B(n_18),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_148),
.A2(n_21),
.B(n_125),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_108),
.C(n_121),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_204),
.C(n_134),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_138),
.B(n_121),
.C(n_67),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g208 ( 
.A1(n_156),
.A2(n_67),
.B1(n_21),
.B2(n_115),
.Y(n_208)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_0),
.B(n_1),
.Y(n_230)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_150),
.B1(n_142),
.B2(n_136),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_147),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_215),
.C(n_222),
.Y(n_247)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_156),
.B1(n_171),
.B2(n_169),
.Y(n_212)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_230),
.B(n_208),
.C(n_194),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_144),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_186),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_219),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_0),
.B(n_1),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_224),
.B(n_232),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_141),
.C(n_170),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_226),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_190),
.A2(n_183),
.B(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_137),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

HAxp5_ASAP7_75t_SL g227 ( 
.A(n_177),
.B(n_170),
.CON(n_227),
.SN(n_227)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_227),
.A2(n_234),
.B(n_237),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_196),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_229),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_0),
.C(n_2),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_233),
.C(n_238),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_3),
.B(n_5),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_3),
.C(n_5),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_3),
.B(n_6),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_185),
.A2(n_6),
.B(n_7),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_172),
.A2(n_10),
.A3(n_13),
.B1(n_8),
.B2(n_9),
.C1(n_6),
.C2(n_7),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_181),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_239),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_225),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_252),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_206),
.B1(n_173),
.B2(n_207),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_263),
.B1(n_227),
.B2(n_235),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_253),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_200),
.B1(n_209),
.B2(n_176),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_250),
.B1(n_261),
.B2(n_232),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_176),
.B1(n_202),
.B2(n_204),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_201),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_230),
.B1(n_234),
.B2(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

OA21x2_ASAP7_75t_SL g255 ( 
.A1(n_212),
.A2(n_195),
.B(n_198),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_217),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_188),
.C(n_191),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_260),
.C(n_262),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_191),
.C(n_187),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_216),
.A2(n_186),
.B1(n_182),
.B2(n_187),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_212),
.A2(n_182),
.B1(n_174),
.B2(n_180),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_267),
.B1(n_273),
.B2(n_244),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_263),
.A2(n_217),
.B1(n_219),
.B2(n_228),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_216),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_269),
.C(n_277),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_222),
.C(n_224),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_248),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_175),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_278),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_251),
.B1(n_256),
.B2(n_248),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_213),
.C(n_233),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_231),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_237),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_174),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_251),
.B1(n_246),
.B2(n_245),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_259),
.B1(n_279),
.B2(n_260),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_245),
.Y(n_285)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_287),
.A2(n_289),
.B(n_291),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_249),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_296),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_243),
.B(n_241),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_243),
.B(n_241),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_230),
.B(n_258),
.C(n_264),
.Y(n_304)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_261),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_269),
.C(n_268),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_278),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_246),
.B1(n_270),
.B2(n_254),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_257),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_264),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_277),
.C(n_257),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_295),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_312),
.B(n_307),
.Y(n_321)
);

AOI31xp67_ASAP7_75t_SL g311 ( 
.A1(n_297),
.A2(n_288),
.A3(n_292),
.B(n_289),
.Y(n_311)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_290),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_291),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_299),
.B(n_290),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_298),
.C(n_306),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_302),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_319),
.C(n_314),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_321),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_303),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_308),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_317),
.B(n_320),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_326),
.A2(n_327),
.B(n_304),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_324),
.C(n_319),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_315),
.Y(n_330)
);


endmodule