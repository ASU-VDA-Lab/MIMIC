module real_jpeg_30549_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_679;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_682;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_704;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_650;
wire n_250;
wire n_254;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_707;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_710;
wire n_703;
wire n_110;
wire n_195;
wire n_533;
wire n_592;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_594;
wire n_316;
wire n_161;
wire n_207;
wire n_711;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_708;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_709;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_268;
wire n_597;
wire n_42;
wire n_313;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_361;
wire n_694;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_0),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_0),
.Y(n_219)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_0),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_2),
.A2(n_241),
.B1(n_244),
.B2(n_245),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_2),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_2),
.A2(n_244),
.B1(n_265),
.B2(n_268),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_2),
.A2(n_244),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_2),
.A2(n_244),
.B1(n_413),
.B2(n_415),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_3),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_4),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_4),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_4),
.A2(n_171),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_4),
.A2(n_171),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

AO22x1_ASAP7_75t_L g671 ( 
.A1(n_4),
.A2(n_171),
.B1(n_645),
.B2(n_672),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_5),
.A2(n_233),
.B1(n_234),
.B2(n_237),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_5),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_5),
.A2(n_168),
.B1(n_233),
.B2(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_5),
.A2(n_233),
.B1(n_463),
.B2(n_466),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g538 ( 
.A1(n_5),
.A2(n_233),
.B1(n_539),
.B2(n_543),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_6),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_6),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_6),
.A2(n_228),
.B1(n_310),
.B2(n_315),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_6),
.A2(n_228),
.B1(n_392),
.B2(n_394),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_6),
.A2(n_228),
.B1(n_491),
.B2(n_495),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_7),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_7),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g420 ( 
.A(n_7),
.B(n_72),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_7),
.A2(n_386),
.B1(n_524),
.B2(n_527),
.Y(n_523)
);

OAI21xp33_ASAP7_75t_L g613 ( 
.A1(n_7),
.A2(n_205),
.B(n_548),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_9),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_10),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_10),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_11),
.A2(n_301),
.B1(n_302),
.B2(n_305),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_11),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_11),
.A2(n_301),
.B1(n_399),
.B2(n_403),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_11),
.A2(n_301),
.B1(n_515),
.B2(n_519),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_11),
.A2(n_301),
.B1(n_597),
.B2(n_600),
.Y(n_596)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_12),
.Y(n_110)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_12),
.Y(n_121)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_12),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_20),
.B(n_710),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_13),
.B(n_711),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_14),
.A2(n_57),
.B1(n_97),
.B2(n_101),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_14),
.A2(n_57),
.B1(n_197),
.B2(n_200),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_14),
.A2(n_57),
.B1(n_525),
.B2(n_650),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_15),
.Y(n_129)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_15),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_16),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_16),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_16),
.A2(n_138),
.B1(n_183),
.B2(n_186),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_16),
.A2(n_138),
.B1(n_352),
.B2(n_354),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_16),
.A2(n_138),
.B1(n_639),
.B2(n_645),
.Y(n_638)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_17),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_17),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_17),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_18),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_18),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_18),
.A2(n_75),
.B1(n_126),
.B2(n_130),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g212 ( 
.A1(n_18),
.A2(n_75),
.B1(n_122),
.B2(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_18),
.A2(n_75),
.B1(n_679),
.B2(n_680),
.Y(n_678)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_83),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_81),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_23),
.B(n_703),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_23),
.B(n_703),
.Y(n_709)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_55),
.B1(n_70),
.B2(n_73),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g82 ( 
.A1(n_24),
.A2(n_70),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_24),
.Y(n_637)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2x1_ASAP7_75t_L g231 ( 
.A(n_25),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_25),
.B(n_223),
.Y(n_272)
);

AO22x1_ASAP7_75t_SL g299 ( 
.A1(n_25),
.A2(n_72),
.B1(n_232),
.B2(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_25),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_35),
.B2(n_38),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_27),
.Y(n_237)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_29),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_29),
.Y(n_646)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_34),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_34),
.Y(n_348)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_38),
.Y(n_344)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_41),
.Y(n_644)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_42),
.Y(n_270)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_45),
.Y(n_137)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_45),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_46),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_46),
.Y(n_243)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_54),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_56),
.A2(n_71),
.B1(n_637),
.B2(n_671),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_62),
.Y(n_236)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_62),
.Y(n_304)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_66),
.Y(n_305)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_67),
.Y(n_267)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_67),
.Y(n_674)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_70),
.Y(n_670)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g263 ( 
.A(n_71),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_71),
.A2(n_264),
.B1(n_637),
.B2(n_638),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_72),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_72),
.B(n_300),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_78),
.Y(n_230)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g333 ( 
.A1(n_80),
.A2(n_334),
.A3(n_340),
.B1(n_343),
.B2(n_345),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_84),
.Y(n_83)
);

AO21x2_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_629),
.B(n_704),
.Y(n_85)
);

NAND2x1_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_446),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_378),
.B(n_442),
.Y(n_87)
);

NOR2xp67_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_324),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_89),
.A2(n_443),
.B(n_444),
.Y(n_442)
);

NOR3xp33_ASAP7_75t_L g447 ( 
.A(n_89),
.B(n_324),
.C(n_448),
.Y(n_447)
);

AOI21x1_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_273),
.B(n_276),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_253),
.Y(n_90)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_91),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_91),
.A2(n_253),
.B1(n_274),
.B2(n_275),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_178),
.B1(n_179),
.B2(n_252),
.Y(n_91)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_92),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_92),
.B(n_178),
.C(n_274),
.Y(n_632)
);

NAND2x1_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_177),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_133),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_94),
.B(n_133),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_103),
.B1(n_125),
.B2(n_132),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_96),
.A2(n_104),
.B1(n_188),
.B2(n_189),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_100),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_102),
.Y(n_185)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

AO22x1_ASAP7_75t_L g389 ( 
.A1(n_103),
.A2(n_132),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_103),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_103),
.A2(n_511),
.B1(n_512),
.B2(n_513),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_103),
.B(n_579),
.Y(n_578)
);

OA21x2_ASAP7_75t_L g654 ( 
.A1(n_103),
.A2(n_125),
.B(n_132),
.Y(n_654)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_104),
.A2(n_182),
.B1(n_188),
.B2(n_189),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_104),
.A2(n_182),
.B1(n_188),
.B2(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_104),
.A2(n_514),
.B1(n_553),
.B2(n_554),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_105)
);

BUFx4f_ASAP7_75t_SL g563 ( 
.A(n_106),
.Y(n_563)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_108),
.Y(n_147)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_108),
.Y(n_476)
);

OAI22x1_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_116),
.B1(n_119),
.B2(n_122),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_110),
.Y(n_574)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_115),
.Y(n_188)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_116),
.Y(n_353)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_117),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_118),
.Y(n_288)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_123),
.Y(n_547)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_124),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_124),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_124),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_127),
.Y(n_395)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_128),
.Y(n_520)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_129),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_129),
.Y(n_487)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_131),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_132),
.B(n_391),
.Y(n_470)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_132),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_144),
.B1(n_167),
.B2(n_175),
.Y(n_133)
);

AOI22x1_ASAP7_75t_L g239 ( 
.A1(n_134),
.A2(n_144),
.B1(n_240),
.B2(n_249),
.Y(n_239)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_143),
.Y(n_339)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_143),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_144),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_144),
.A2(n_175),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_144),
.B(n_309),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g648 ( 
.A1(n_144),
.A2(n_167),
.B1(n_175),
.B2(n_649),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_144),
.B(n_649),
.Y(n_682)
);

OA21x2_ASAP7_75t_SL g696 ( 
.A1(n_144),
.A2(n_175),
.B(n_697),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_158),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_145),
.Y(n_249)
);

AOI22x1_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_148),
.B1(n_151),
.B2(n_154),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_159),
.B1(n_162),
.B2(n_165),
.Y(n_158)
);

INVx5_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_150),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_156),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g469 ( 
.A(n_157),
.Y(n_469)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_165),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_170),
.Y(n_402)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_170),
.Y(n_527)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_176),
.A2(n_307),
.B1(n_308),
.B2(n_319),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_176),
.A2(n_409),
.B(n_410),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_R g551 ( 
.A(n_176),
.B(n_386),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_176),
.A2(n_677),
.B(n_682),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_177),
.A2(n_635),
.B1(n_656),
.B2(n_657),
.Y(n_634)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_177),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_220),
.B(n_250),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_180),
.B(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_195),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_181),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_188),
.Y(n_511)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2x2_ASAP7_75t_L g374 ( 
.A(n_195),
.B(n_375),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_205),
.B1(n_211),
.B2(n_215),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_196),
.A2(n_205),
.B1(n_283),
.B2(n_285),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_198),
.Y(n_560)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_199),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_199),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_199),
.Y(n_572)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_205),
.B(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_205),
.A2(n_351),
.B1(n_412),
.B2(n_417),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_205),
.A2(n_538),
.B(n_548),
.Y(n_537)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_206),
.A2(n_286),
.B1(n_350),
.B2(n_357),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_206),
.B(n_490),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_206),
.A2(n_591),
.B1(n_594),
.B2(n_595),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_209),
.Y(n_418)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_SL g550 ( 
.A(n_210),
.Y(n_550)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_213),
.Y(n_414)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx2_ASAP7_75t_R g284 ( 
.A(n_218),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_219),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_238),
.Y(n_220)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_221),
.A2(n_238),
.B1(n_239),
.B2(n_251),
.Y(n_279)
);

NAND2x1_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_231),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_222),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_249),
.B(n_309),
.Y(n_372)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_261),
.Y(n_253)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_254),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_255),
.A2(n_260),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_255),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_259),
.Y(n_593)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_260),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_262),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_271),
.Y(n_262)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_268),
.Y(n_385)
);

INVx11_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_272),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_276),
.B(n_445),
.Y(n_444)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.C(n_320),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_278),
.B(n_321),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_280),
.B(n_377),
.Y(n_376)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_299),
.C(n_306),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_R g326 ( 
.A1(n_281),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_293),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_282),
.B(n_293),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx2_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_291),
.Y(n_497)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_292),
.Y(n_542)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_294),
.Y(n_390)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_296),
.Y(n_465)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_298),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_306),
.Y(n_327)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_313),
.Y(n_485)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_314),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_314),
.Y(n_652)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_319),
.A2(n_367),
.B(n_372),
.Y(n_366)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_319),
.A2(n_372),
.B(n_523),
.Y(n_522)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_322),
.A2(n_659),
.B(n_660),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_376),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_325),
.B(n_376),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.C(n_373),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_327),
.A2(n_328),
.B1(n_374),
.B2(n_441),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_329),
.B(n_331),
.Y(n_439)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_362),
.C(n_365),
.Y(n_331)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_332),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_349),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g405 ( 
.A(n_333),
.B(n_349),
.Y(n_405)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_338),
.Y(n_346)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx2_ASAP7_75t_SL g599 ( 
.A(n_356),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_357),
.B(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_362),
.A2(n_363),
.B1(n_365),
.B2(n_366),
.Y(n_431)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_367),
.Y(n_397)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_368),
.Y(n_679)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_434),
.C(n_437),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_421),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_380),
.B(n_421),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_405),
.C(n_406),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_381),
.B(n_501),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_388),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_382),
.B(n_389),
.C(n_426),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_386),
.B(n_387),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_386),
.B(n_474),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_386),
.B(n_484),
.C(n_486),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_386),
.B(n_576),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_386),
.A2(n_575),
.B(n_580),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g607 ( 
.A(n_386),
.B(n_553),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_386),
.B(n_616),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_396),
.Y(n_388)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_391),
.Y(n_554)
);

INVx3_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_398),
.Y(n_409)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_405),
.A2(n_406),
.B1(n_407),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_411),
.C(n_419),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_408),
.B(n_457),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_411),
.A2(n_419),
.B1(n_420),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_428),
.B(n_432),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_433),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_425),
.B2(n_427),
.Y(n_422)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_425),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_427),
.Y(n_436)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_435),
.C(n_436),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_429),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_434),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_438),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_438),
.A2(n_449),
.B(n_450),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_451),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_503),
.B(n_627),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_500),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_454),
.B(n_628),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_459),
.C(n_471),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_456),
.B(n_529),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_459),
.A2(n_460),
.B1(n_471),
.B2(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_461),
.A2(n_462),
.B(n_470),
.Y(n_460)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_462),
.Y(n_512)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_470),
.B(n_578),
.Y(n_577)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_471),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_488),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_488),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_477),
.B(n_483),
.Y(n_472)
);

INVx4_ASAP7_75t_SL g474 ( 
.A(n_475),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_486),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_498),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_489),
.A2(n_596),
.B(n_609),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_490),
.B(n_549),
.Y(n_548)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_500),
.Y(n_628)
);

AOI21x1_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_531),
.B(n_626),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_528),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_L g626 ( 
.A(n_505),
.B(n_528),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_508),
.C(n_521),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_510),
.B(n_522),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_525),
.Y(n_681)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_586),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_533),
.A2(n_555),
.B(n_585),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_536),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_534),
.B(n_536),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_551),
.C(n_552),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_537),
.A2(n_582),
.B1(n_583),
.B2(n_584),
.Y(n_581)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_537),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_538),
.Y(n_594)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_541),
.Y(n_600)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_551),
.B(n_552),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_581),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_556),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_577),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_557),
.A2(n_577),
.B1(n_602),
.B2(n_603),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_557),
.Y(n_602)
);

AO221x1_ASAP7_75t_L g622 ( 
.A1(n_557),
.A2(n_577),
.B1(n_590),
.B2(n_602),
.C(n_603),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_558),
.A2(n_561),
.B(n_569),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_564),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_570),
.A2(n_573),
.B(n_575),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_577),
.Y(n_603)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_581),
.Y(n_624)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_582),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_585),
.B(n_587),
.C(n_623),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_588),
.A2(n_604),
.B(n_622),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_590),
.B(n_601),
.Y(n_589)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_591),
.Y(n_616)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_593),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_606),
.A2(n_612),
.B(n_621),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_607),
.B(n_608),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_607),
.B(n_608),
.Y(n_621)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_613),
.B(n_614),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_615),
.B(n_617),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_625),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g629 ( 
.A(n_630),
.B(n_688),
.C(n_702),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_631),
.B(n_661),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_632),
.B(n_633),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g707 ( 
.A(n_632),
.B(n_633),
.Y(n_707)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_634),
.B(n_658),
.Y(n_633)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_635),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_635),
.Y(n_685)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_636),
.B(n_647),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_636),
.Y(n_664)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_636),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_SL g669 ( 
.A1(n_637),
.A2(n_638),
.B1(n_670),
.B2(n_671),
.Y(n_669)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_641),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_642),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_648),
.A2(n_653),
.B1(n_654),
.B2(n_655),
.Y(n_647)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_648),
.Y(n_655)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_652),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_653),
.A2(n_654),
.B1(n_676),
.B2(n_683),
.Y(n_675)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_654),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_654),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_655),
.B(n_664),
.C(n_665),
.Y(n_663)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_656),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_658),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_661),
.A2(n_689),
.B(n_707),
.C(n_708),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_662),
.B(n_684),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_662),
.B(n_684),
.Y(n_708)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_663),
.B(n_666),
.Y(n_662)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_663),
.Y(n_701)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_665),
.Y(n_694)
);

XNOR2xp5_ASAP7_75t_L g666 ( 
.A(n_667),
.B(n_668),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g699 ( 
.A(n_667),
.B(n_700),
.C(n_701),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_668),
.Y(n_700)
);

XNOR2xp5_ASAP7_75t_L g668 ( 
.A(n_669),
.B(n_675),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_669),
.Y(n_692)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_673),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_674),
.Y(n_673)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_676),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_676),
.Y(n_693)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_678),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_678),
.Y(n_697)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_681),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g684 ( 
.A(n_685),
.B(n_686),
.C(n_687),
.Y(n_684)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_689),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_690),
.B(n_699),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_690),
.B(n_699),
.Y(n_705)
);

XNOR2xp5_ASAP7_75t_L g690 ( 
.A(n_691),
.B(n_695),
.Y(n_690)
);

MAJIxp5_ASAP7_75t_L g703 ( 
.A(n_691),
.B(n_696),
.C(n_698),
.Y(n_703)
);

MAJIxp5_ASAP7_75t_L g691 ( 
.A(n_692),
.B(n_693),
.C(n_694),
.Y(n_691)
);

XNOR2xp5_ASAP7_75t_L g695 ( 
.A(n_696),
.B(n_698),
.Y(n_695)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_702),
.A2(n_705),
.B(n_706),
.C(n_709),
.Y(n_704)
);


endmodule