module fake_jpeg_29779_n_452 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_452);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_452;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_6),
.B(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_5),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_64),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_51),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_0),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_43),
.Y(n_110)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_61),
.B(n_79),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_74),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_71),
.Y(n_105)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx11_ASAP7_75t_SL g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_16),
.B(n_1),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_77),
.Y(n_118)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_16),
.B(n_1),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_17),
.A2(n_14),
.B1(n_3),
.B2(n_4),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_75),
.A2(n_28),
.B1(n_46),
.B2(n_35),
.Y(n_114)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_26),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_26),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_18),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_87),
.Y(n_112)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_28),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_36),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_5),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_6),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_21),
.Y(n_138)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_33),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_40),
.B1(n_25),
.B2(n_45),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_98),
.A2(n_114),
.B1(n_131),
.B2(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_138),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_45),
.B1(n_25),
.B2(n_17),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_102),
.B(n_110),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_31),
.B1(n_17),
.B2(n_45),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_125),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_53),
.A2(n_31),
.B1(n_46),
.B2(n_22),
.Y(n_125)
);

NAND2x1_ASAP7_75t_L g126 ( 
.A(n_55),
.B(n_37),
.Y(n_126)
);

NAND2x1p5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_37),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_56),
.A2(n_37),
.B1(n_43),
.B2(n_20),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_128),
.A2(n_92),
.A3(n_69),
.B1(n_67),
.B2(n_12),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_31),
.B1(n_33),
.B2(n_26),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_83),
.A2(n_33),
.B1(n_42),
.B2(n_30),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_49),
.A2(n_33),
.B1(n_42),
.B2(n_30),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_63),
.B1(n_81),
.B2(n_73),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_57),
.A2(n_22),
.B1(n_35),
.B2(n_34),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_141),
.Y(n_161)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_50),
.B(n_34),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_143),
.Y(n_186)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx4_ASAP7_75t_SL g229 ( 
.A(n_147),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_170),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_150),
.B(n_153),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_112),
.B(n_70),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_151),
.B(n_111),
.Y(n_232)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_106),
.A2(n_37),
.B(n_82),
.C(n_93),
.Y(n_153)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_39),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_156),
.B(n_164),
.Y(n_202)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_110),
.A2(n_54),
.B(n_37),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_159),
.A2(n_124),
.B(n_10),
.Y(n_228)
);

NOR2x1_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_29),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_162),
.B(n_134),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_101),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

BUFx24_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_168),
.A2(n_195),
.B1(n_10),
.B2(n_11),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_103),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_170),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_82),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_95),
.B(n_29),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_185),
.Y(n_203)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_33),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_178),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_119),
.B(n_144),
.C(n_126),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_187),
.C(n_193),
.Y(n_235)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_66),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_190),
.Y(n_225)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_102),
.B(n_62),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_121),
.B(n_76),
.C(n_86),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_127),
.B(n_60),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_127),
.B(n_78),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_96),
.B(n_66),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_98),
.B1(n_131),
.B2(n_94),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_96),
.B(n_92),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_9),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_121),
.B(n_9),
.C(n_10),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_145),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_197),
.B(n_210),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_132),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_200),
.B(n_227),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_211),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_169),
.A2(n_123),
.B(n_94),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_145),
.B1(n_104),
.B2(n_129),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_213),
.A2(n_226),
.B1(n_185),
.B2(n_187),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_130),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_224),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_161),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_221),
.B(n_222),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_154),
.B(n_122),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_237),
.B1(n_238),
.B2(n_149),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_130),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_158),
.A2(n_129),
.B1(n_122),
.B2(n_124),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_153),
.A2(n_123),
.B(n_111),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_228),
.A2(n_159),
.B(n_177),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_176),
.CI(n_149),
.CON(n_243),
.SN(n_243)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_147),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_167),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_158),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_148),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_241),
.A2(n_244),
.B1(n_266),
.B2(n_235),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_242),
.A2(n_248),
.B1(n_249),
.B2(n_253),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_215),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_191),
.B1(n_184),
.B2(n_161),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_225),
.A2(n_172),
.B1(n_155),
.B2(n_165),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_246),
.A2(n_276),
.B1(n_254),
.B2(n_271),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_221),
.A2(n_184),
.B1(n_189),
.B2(n_188),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_201),
.A2(n_193),
.B1(n_157),
.B2(n_160),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_267),
.B(n_228),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_152),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_261),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_203),
.A2(n_175),
.B1(n_182),
.B2(n_163),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_254),
.A2(n_229),
.B1(n_208),
.B2(n_206),
.Y(n_281)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_256),
.B(n_258),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_197),
.B(n_162),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_202),
.B(n_205),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_259),
.Y(n_293)
);

AOI32xp33_ASAP7_75t_L g260 ( 
.A1(n_199),
.A2(n_181),
.A3(n_166),
.B1(n_165),
.B2(n_183),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_262),
.Y(n_282)
);

AO22x1_ASAP7_75t_SL g261 ( 
.A1(n_200),
.A2(n_174),
.B1(n_179),
.B2(n_166),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_203),
.B(n_12),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_14),
.Y(n_263)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_263),
.Y(n_302)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_207),
.A2(n_238),
.B1(n_232),
.B2(n_237),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_207),
.B(n_211),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_214),
.Y(n_269)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_215),
.B(n_235),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_196),
.Y(n_291)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_208),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_196),
.Y(n_273)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_231),
.Y(n_274)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_274),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_224),
.B(n_218),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_275),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_227),
.A2(n_226),
.B1(n_213),
.B2(n_229),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_277),
.A2(n_292),
.B(n_295),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_300),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_240),
.A2(n_267),
.B(n_266),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_284),
.A2(n_290),
.B(n_245),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_291),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_242),
.A2(n_230),
.B1(n_220),
.B2(n_206),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_289),
.A2(n_298),
.B1(n_254),
.B2(n_273),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_240),
.A2(n_212),
.B(n_218),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_240),
.A2(n_212),
.B(n_231),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_231),
.B(n_216),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_257),
.A2(n_204),
.B(n_234),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_297),
.A2(n_304),
.B(n_308),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_248),
.A2(n_209),
.B1(n_220),
.B2(n_230),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_204),
.C(n_216),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_306),
.C(n_243),
.Y(n_328)
);

OA22x2_ASAP7_75t_L g300 ( 
.A1(n_244),
.A2(n_209),
.B1(n_231),
.B2(n_241),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_264),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_252),
.A2(n_251),
.B(n_247),
.C(n_258),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_247),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_249),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_239),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_314),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_315),
.B(n_319),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_303),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_321),
.Y(n_344)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_253),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_320),
.A2(n_326),
.B1(n_300),
.B2(n_290),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_295),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_281),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_324),
.Y(n_352)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_325),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_278),
.A2(n_300),
.B1(n_277),
.B2(n_285),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_292),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_327),
.B(n_331),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_338),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_334),
.B(n_297),
.Y(n_343)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_250),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_261),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_333),
.B(n_339),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_284),
.A2(n_261),
.B(n_274),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_268),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_335),
.B(n_308),
.Y(n_350)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_337),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_243),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_289),
.B(n_298),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_306),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_348),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_343),
.A2(n_360),
.B(n_336),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_323),
.A2(n_300),
.B1(n_282),
.B2(n_279),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_347),
.A2(n_356),
.B1(n_320),
.B2(n_339),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_338),
.B(n_279),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_349),
.A2(n_358),
.B1(n_361),
.B2(n_329),
.Y(n_378)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_350),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_316),
.B(n_288),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_331),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_311),
.A2(n_307),
.B1(n_296),
.B2(n_301),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_326),
.A2(n_312),
.B1(n_333),
.B2(n_320),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_309),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_332),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_334),
.A2(n_301),
.B(n_296),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_326),
.A2(n_307),
.B1(n_280),
.B2(n_283),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_344),
.B(n_314),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_370),
.Y(n_391)
);

XNOR2x1_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_328),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_373),
.C(n_379),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_374),
.Y(n_389)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_340),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_372),
.Y(n_392)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_352),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_345),
.C(n_342),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_335),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_376),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_315),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_377),
.A2(n_351),
.B(n_353),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_378),
.A2(n_347),
.B1(n_349),
.B2(n_346),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_332),
.C(n_336),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_351),
.B(n_332),
.Y(n_380)
);

NOR4xp25_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_385),
.C(n_362),
.D(n_317),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_364),
.A2(n_312),
.B1(n_322),
.B2(n_321),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_382),
.Y(n_402)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_353),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_384),
.C(n_358),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_318),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g385 ( 
.A(n_346),
.B(n_318),
.CI(n_327),
.CON(n_385),
.SN(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_365),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_395),
.Y(n_410)
);

INVx13_ASAP7_75t_L g387 ( 
.A(n_385),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_360),
.B(n_364),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_390),
.A2(n_394),
.B(n_370),
.Y(n_409)
);

AOI21x1_ASAP7_75t_L g394 ( 
.A1(n_384),
.A2(n_363),
.B(n_319),
.Y(n_394)
);

NAND4xp25_ASAP7_75t_SL g395 ( 
.A(n_378),
.B(n_356),
.C(n_255),
.D(n_354),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_375),
.Y(n_411)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_397),
.B(n_398),
.C(n_401),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_361),
.C(n_362),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_391),
.C(n_390),
.Y(n_408)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_366),
.Y(n_400)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_400),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_367),
.C(n_379),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_406),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_383),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_369),
.C(n_366),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_412),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_409),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_411),
.A2(n_410),
.B1(n_393),
.B2(n_395),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_369),
.C(n_381),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_391),
.Y(n_413)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_413),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_385),
.C(n_372),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_392),
.Y(n_424)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_414),
.B(n_401),
.CI(n_387),
.CON(n_416),
.SN(n_416)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_418),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_408),
.B(n_386),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_313),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_415),
.A2(n_402),
.B1(n_393),
.B2(n_400),
.Y(n_420)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_420),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_415),
.A2(n_402),
.B1(n_387),
.B2(n_396),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_424),
.Y(n_434)
);

NOR2x1_ASAP7_75t_SL g426 ( 
.A(n_403),
.B(n_394),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_426),
.A2(n_403),
.B(n_392),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_382),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_427),
.B(n_371),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_423),
.C(n_425),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_431),
.Y(n_439)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_430),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_417),
.B(n_283),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_L g440 ( 
.A1(n_433),
.A2(n_436),
.B(n_330),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_425),
.A2(n_352),
.B(n_325),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_435),
.A2(n_427),
.B1(n_337),
.B2(n_313),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_432),
.B(n_416),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_437),
.B(n_438),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_442),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_416),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_439),
.A2(n_434),
.B(n_430),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_444),
.Y(n_447)
);

AOI21xp33_ASAP7_75t_L g445 ( 
.A1(n_439),
.A2(n_422),
.B(n_420),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_445),
.B(n_441),
.Y(n_448)
);

NOR3xp33_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_443),
.C(n_446),
.Y(n_449)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_447),
.C(n_418),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_450),
.A2(n_324),
.B(n_265),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_269),
.Y(n_452)
);


endmodule