module fake_jpeg_10659_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_19),
.Y(n_50)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_43),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_22),
.B1(n_32),
.B2(n_30),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_26),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_60),
.Y(n_91)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_22),
.B1(n_32),
.B2(n_30),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_32),
.B1(n_25),
.B2(n_27),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_34),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_72),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_76),
.B1(n_84),
.B2(n_51),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_83),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_25),
.B1(n_16),
.B2(n_21),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_77),
.B1(n_91),
.B2(n_72),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_21),
.B1(n_20),
.B2(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_29),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_77),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_29),
.B(n_18),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_90),
.B(n_3),
.Y(n_101)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_28),
.B1(n_17),
.B2(n_29),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_28),
.B1(n_17),
.B2(n_18),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_56),
.B1(n_58),
.B2(n_65),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_18),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_3),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_56),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_101),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_18),
.B(n_28),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_66),
.B(n_86),
.Y(n_123)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_105),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_69),
.B1(n_88),
.B2(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_54),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_114),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_89),
.Y(n_112)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_49),
.B1(n_65),
.B2(n_53),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_49),
.B1(n_71),
.B2(n_80),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_4),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_81),
.C(n_80),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_126),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_123),
.B(n_101),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_113),
.B1(n_105),
.B2(n_112),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_71),
.B(n_5),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_4),
.C(n_5),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_128),
.B(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_4),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_134),
.B(n_7),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_139),
.B(n_148),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_151),
.B1(n_126),
.B2(n_116),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_13),
.A3(n_15),
.B1(n_14),
.B2(n_11),
.C1(n_9),
.C2(n_6),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_120),
.B(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_109),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_144),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_150),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_103),
.B1(n_106),
.B2(n_8),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_11),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_6),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_123),
.B(n_118),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_159),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_115),
.C(n_117),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_135),
.C(n_136),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_119),
.B(n_132),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_116),
.B1(n_124),
.B2(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_147),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_170),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_171),
.C(n_154),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_136),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_146),
.C(n_125),
.Y(n_171)
);

OAI322xp33_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_150),
.A3(n_146),
.B1(n_151),
.B2(n_148),
.C1(n_122),
.C2(n_125),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_174),
.A2(n_161),
.B1(n_164),
.B2(n_156),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_154),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_169),
.B(n_166),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_180),
.B(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_165),
.B(n_163),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_178),
.B(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_181),
.A2(n_167),
.B(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_184),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_172),
.B1(n_155),
.B2(n_170),
.Y(n_184)
);

XOR2x1_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_182),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.C(n_194),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_179),
.B1(n_131),
.B2(n_103),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_179),
.C(n_131),
.Y(n_194)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_188),
.B(n_8),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_7),
.B(n_8),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_195),
.Y(n_198)
);


endmodule