module real_jpeg_13923_n_17 (n_5, n_4, n_8, n_0, n_12, n_339, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_339;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_3),
.A2(n_34),
.B1(n_53),
.B2(n_54),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_3),
.A2(n_34),
.B1(n_64),
.B2(n_66),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_134),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_5),
.A2(n_64),
.B1(n_66),
.B2(n_134),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_134),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_6),
.A2(n_64),
.B1(n_66),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_6),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_6),
.B(n_54),
.C(n_69),
.Y(n_166)
);

NAND2x1_ASAP7_75t_SL g170 ( 
.A(n_6),
.B(n_90),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_6),
.A2(n_125),
.B(n_178),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_6),
.A2(n_24),
.B(n_89),
.C(n_205),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_162),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_6),
.B(n_21),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_6),
.B(n_31),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_7),
.A2(n_38),
.B1(n_64),
.B2(n_66),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_38),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_7),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_9),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_9),
.A2(n_64),
.B1(n_66),
.B2(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_92),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_10),
.A2(n_64),
.B1(n_66),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_10),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_174),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_174),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_174),
.Y(n_276)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_77),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_77),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_12),
.A2(n_64),
.B1(n_66),
.B2(n_77),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_64),
.B1(n_66),
.B2(n_81),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_81),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_81),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_15),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_63),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_63),
.Y(n_266)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_33),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_21),
.A2(n_28),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_21),
.A2(n_28),
.B1(n_37),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_22),
.A2(n_76),
.B(n_78),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_22),
.A2(n_29),
.B1(n_76),
.B2(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_22),
.B(n_80),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_22),
.A2(n_29),
.B1(n_110),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_22),
.A2(n_78),
.B(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_22),
.A2(n_29),
.B1(n_133),
.B2(n_276),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

NAND2xp33_ASAP7_75t_SL g262 ( 
.A(n_23),
.B(n_25),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_24),
.A2(n_25),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g261 ( 
.A1(n_24),
.A2(n_27),
.A3(n_32),
.B1(n_249),
.B2(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_28),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_29),
.A2(n_133),
.B(n_135),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_29),
.A2(n_32),
.B(n_162),
.C(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_35),
.B(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_36),
.B(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_333),
.B(n_335),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_321),
.B(n_332),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_150),
.B(n_318),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_137),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_112),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_46),
.B(n_112),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_82),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_47),
.B(n_83),
.C(n_98),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_75),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_48),
.A2(n_49),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_60),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_50),
.A2(n_51),
.B1(n_75),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_50),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_57),
.B(n_58),
.Y(n_51)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_52),
.A2(n_57),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_52),
.B(n_179),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_52),
.A2(n_57),
.B1(n_124),
.B2(n_266),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_53),
.B(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_57),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_57),
.B(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_59),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_72),
.B2(n_74),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_62),
.A2(n_67),
.B1(n_74),
.B2(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_64),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_66),
.B1(n_88),
.B2(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_64),
.B(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_66),
.A2(n_88),
.B(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_74),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_67),
.B(n_164),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_67),
.A2(n_74),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_67),
.A2(n_74),
.B1(n_129),
.B2(n_255),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_73),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_71),
.A2(n_173),
.B(n_175),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_71),
.B(n_162),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_71),
.A2(n_175),
.B(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_74),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_98),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_84),
.B(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_95),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_85),
.A2(n_91),
.B1(n_93),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_85),
.A2(n_93),
.B1(n_103),
.B2(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_85),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_85),
.A2(n_93),
.B1(n_225),
.B2(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_85),
.A2(n_211),
.B(n_252),
.Y(n_274)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_90),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_86),
.B(n_212),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_86),
.A2(n_90),
.B(n_325),
.Y(n_324)
);

NOR2x1_ASAP7_75t_R g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_90),
.B(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_93),
.A2(n_225),
.B(n_226),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_93),
.A2(n_131),
.B(n_226),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_96),
.A2(n_161),
.B(n_163),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_96),
.A2(n_163),
.B(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_SL g148 ( 
.A(n_100),
.B(n_105),
.C(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_105),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_105),
.B(n_142),
.C(n_146),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_109),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_109),
.B(n_141),
.C(n_148),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_119),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_118),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_119),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_130),
.C(n_132),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_120),
.A2(n_121),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_122),
.A2(n_127),
.B1(n_128),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_122),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_125),
.A2(n_126),
.B1(n_207),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_125),
.A2(n_126),
.B1(n_232),
.B2(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_126),
.A2(n_184),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_126),
.B(n_162),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_126),
.A2(n_192),
.B(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_130),
.B(n_132),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_136),
.B(n_247),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_L g318 ( 
.A1(n_137),
.A2(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_149),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_138),
.B(n_149),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_148),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_143),
.Y(n_327)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_147),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_312),
.B(n_317),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_300),
.B(n_311),
.Y(n_151)
);

OAI321xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_268),
.A3(n_293),
.B1(n_298),
.B2(n_299),
.C(n_339),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_241),
.B(n_267),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_219),
.B(n_240),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_200),
.B(n_218),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_180),
.B(n_199),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_167),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_158),
.B(n_167),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_160),
.B1(n_165),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_172),
.C(n_176),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_188),
.B(n_198),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_182),
.B(n_186),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_193),
.B(n_197),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_190),
.B(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_202),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_213),
.C(n_217),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_206),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_221),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_233),
.B2(n_234),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_236),
.C(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_228),
.C(n_231),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_243),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_257),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_258),
.C(n_259),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_250),
.B2(n_256),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_251),
.C(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_264),
.Y(n_278)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_283),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_283),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_279),
.C(n_282),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_270),
.A2(n_271),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_277),
.C(n_278),
.Y(n_292)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_279),
.B(n_282),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_281),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_292),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_287),
.C(n_292),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_290),
.C(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_310),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_310),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_305),
.C(n_306),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_331),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_331),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_330),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_326),
.B1(n_328),
.B2(n_329),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_326),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_328),
.C(n_330),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_334),
.Y(n_337)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);


endmodule