module real_jpeg_10378_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_244;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_1),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_61),
.B1(n_67),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_3),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_88),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_88),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_88),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_38),
.B(n_42),
.C(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_38),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_7),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_7),
.B(n_50),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_9),
.A2(n_61),
.B1(n_67),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_9),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_137),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_137),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_137),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_10),
.A2(n_40),
.B1(n_50),
.B2(n_51),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_56),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_11),
.A2(n_56),
.B1(n_61),
.B2(n_67),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_56),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_12),
.A2(n_61),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_70),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_70),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_13),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_15),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_15),
.A2(n_51),
.B(n_63),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_15),
.A2(n_61),
.B1(n_67),
.B2(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_15),
.B(n_164),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_15),
.A2(n_38),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_15),
.B(n_38),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_15),
.A2(n_26),
.B1(n_33),
.B2(n_215),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_15),
.A2(n_50),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_15),
.B(n_50),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_16),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_46),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_16),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_17),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_17),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_17),
.A2(n_50),
.B1(n_51),
.B2(n_68),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_68),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_17),
.A2(n_38),
.B1(n_39),
.B2(n_68),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_122),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_21),
.B(n_92),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.C(n_78),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_22),
.A2(n_23),
.B1(n_72),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_47),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_24),
.B(n_58),
.C(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_25),
.B(n_36),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_26),
.A2(n_33),
.B(n_34),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_26),
.A2(n_33),
.B1(n_81),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_26),
.A2(n_33),
.B1(n_198),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_26),
.A2(n_33),
.B1(n_200),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_26),
.A2(n_33),
.B1(n_231),
.B2(n_247),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_27),
.A2(n_28),
.B1(n_145),
.B2(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_27),
.A2(n_28),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_29),
.B(n_44),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_29),
.B(n_220),
.Y(n_219)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_30),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_33),
.B(n_141),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_37),
.A2(n_41),
.B1(n_43),
.B2(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_38),
.B(n_54),
.Y(n_244)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_39),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_41),
.A2(n_43),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_41),
.A2(n_43),
.B1(n_206),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_41),
.A2(n_43),
.B1(n_229),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_41),
.A2(n_43),
.B1(n_167),
.B2(n_237),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_42),
.Y(n_210)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_43),
.B(n_141),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_58),
.B1(n_59),
.B2(n_71),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_53),
.B1(n_55),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_49),
.A2(n_53),
.B1(n_91),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_49),
.A2(n_53),
.B1(n_132),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_49),
.A2(n_53),
.B1(n_160),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_49),
.A2(n_53),
.B1(n_184),
.B2(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_52),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_53),
.B(n_141),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_57),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_65),
.B1(n_66),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_60),
.A2(n_65),
.B1(n_69),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_60),
.A2(n_65),
.B1(n_87),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_60),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_62),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_61),
.A2(n_62),
.B(n_141),
.C(n_142),
.Y(n_140)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_65),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_72),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_74),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_75),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_78),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.C(n_89),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_82),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_84),
.A2(n_99),
.B1(n_102),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_118),
.B2(n_119),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_109),
.B2(n_110),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_103),
.B(n_108),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_103),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_113),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_118),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_149),
.B(n_271),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_146),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_124),
.B(n_146),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_128),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_127),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_128),
.A2(n_129),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_133),
.C(n_138),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_189),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_171),
.B(n_188),
.Y(n_151)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_152),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_168),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_168),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_157),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_165),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_159),
.B1(n_165),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_172),
.B(n_174),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_180),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_175),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_178),
.Y(n_267)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_186),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_182),
.A2(n_183),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_185),
.B(n_186),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_187),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_269),
.C(n_270),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_263),
.B(n_268),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_249),
.B(n_262),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_233),
.B(n_248),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_223),
.B(n_232),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_212),
.B(n_222),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_196),
.B(n_201),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_207),
.B2(n_211),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_211),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_205),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_207),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_217),
.B(n_221),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_225),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_228),
.C(n_230),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_235),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_235),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.CI(n_241),
.CON(n_235),
.SN(n_235)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_240),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_246),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_250),
.B(n_251),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_257),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_259),
.C(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_258),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_259),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);


endmodule