module fake_jpeg_24288_n_288 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx2_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_13),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_45),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_24),
.B1(n_17),
.B2(n_26),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_18),
.B1(n_15),
.B2(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_28),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_58),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_33),
.A2(n_24),
.B1(n_20),
.B2(n_18),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_15),
.B1(n_26),
.B2(n_22),
.Y(n_73)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_24),
.B1(n_20),
.B2(n_26),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_69),
.B1(n_78),
.B2(n_49),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_71),
.B1(n_73),
.B2(n_75),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_45),
.B1(n_39),
.B2(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_15),
.B1(n_26),
.B2(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_42),
.A2(n_15),
.B1(n_22),
.B2(n_16),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_51),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_27),
.B1(n_14),
.B2(n_19),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_43),
.B1(n_42),
.B2(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_86),
.B1(n_93),
.B2(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_87),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_43),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_97),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_50),
.C(n_48),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_94),
.C(n_65),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_95),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_56),
.B1(n_41),
.B2(n_40),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_0),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_21),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_56),
.B1(n_41),
.B2(n_40),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_67),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_76),
.B1(n_74),
.B2(n_59),
.Y(n_108)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_113),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_120),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_92),
.C(n_89),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_112),
.C(n_115),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_64),
.C(n_73),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_64),
.C(n_68),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_68),
.C(n_78),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_72),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_14),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_94),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_70),
.B1(n_72),
.B2(n_27),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_85),
.B1(n_55),
.B2(n_60),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_70),
.B1(n_41),
.B2(n_56),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_55),
.B1(n_85),
.B2(n_80),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_134),
.B(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_138),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_94),
.B(n_102),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_137),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_88),
.A3(n_84),
.B1(n_14),
.B2(n_27),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_76),
.B1(n_84),
.B2(n_88),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_141),
.B1(n_148),
.B2(n_85),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_103),
.B1(n_126),
.B2(n_76),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_91),
.B(n_101),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_112),
.B(n_125),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_117),
.C(n_96),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_109),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_166),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_139),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_156),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_147),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_157),
.C(n_163),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_114),
.B1(n_113),
.B2(n_107),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_131),
.B1(n_137),
.B2(n_142),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_120),
.A3(n_111),
.B1(n_114),
.B2(n_119),
.C1(n_115),
.C2(n_14),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_79),
.B(n_19),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_146),
.B(n_129),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_162),
.B1(n_13),
.B2(n_12),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_96),
.B1(n_16),
.B2(n_79),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_34),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_174),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_99),
.C(n_34),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_99),
.B(n_21),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_171),
.B(n_31),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_32),
.C(n_31),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_150),
.C(n_134),
.Y(n_170)
);

AOI21x1_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_21),
.B(n_32),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_128),
.B(n_21),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_132),
.C(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_0),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_165),
.B1(n_173),
.B2(n_170),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_178),
.B1(n_182),
.B2(n_192),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_196),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_187),
.B1(n_3),
.B2(n_4),
.Y(n_211)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_139),
.B1(n_136),
.B2(n_2),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_184),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_3),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_169),
.C(n_172),
.Y(n_201)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_190),
.B(n_198),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_166),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_193),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_11),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_154),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_159),
.B1(n_153),
.B2(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_159),
.B1(n_151),
.B2(n_11),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_186),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_0),
.C(n_1),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_189),
.C(n_191),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_211),
.B1(n_190),
.B2(n_187),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_3),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_198),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_216),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_177),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_4),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_4),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_5),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_223),
.C(n_229),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_193),
.C(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_188),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_224),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_227),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_216),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_177),
.C(n_180),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_232),
.B1(n_209),
.B2(n_199),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_194),
.C(n_6),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_217),
.C(n_8),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_194),
.B1(n_6),
.B2(n_8),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_201),
.B(n_208),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_245),
.C(n_246),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_247),
.Y(n_259)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_233),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_9),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_222),
.C(n_219),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_5),
.C(n_8),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_SL g247 ( 
.A(n_231),
.B(n_5),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_235),
.A2(n_243),
.B1(n_239),
.B2(n_242),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_261),
.C(n_10),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_234),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_233),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_260),
.Y(n_264)
);

BUFx4f_ASAP7_75t_SL g258 ( 
.A(n_242),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_258),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_9),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_249),
.B(n_238),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_258),
.B(n_241),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_268),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_244),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_267),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_246),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_9),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_250),
.B(n_10),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_256),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_274),
.B(n_251),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_264),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_273),
.B(n_253),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_272),
.B(n_259),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_285),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_283),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_276),
.Y(n_288)
);


endmodule