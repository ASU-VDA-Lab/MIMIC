module fake_jpeg_14293_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_6),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_15),
.B(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_68),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_74),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_45),
.B1(n_47),
.B2(n_54),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_48),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_48),
.C(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_4),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_45),
.B1(n_56),
.B2(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_52),
.B1(n_51),
.B2(n_49),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_3),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_75),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_20),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_72),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_10),
.C(n_11),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_12),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_66),
.A3(n_71),
.B1(n_6),
.B2(n_7),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_41),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_104),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_105),
.B1(n_109),
.B2(n_18),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_5),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_105)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_28),
.B1(n_37),
.B2(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_108),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_12),
.B1(n_13),
.B2(n_17),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_112),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_128)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_23),
.B(n_24),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_31),
.Y(n_120)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_34),
.A3(n_107),
.B1(n_121),
.B2(n_113),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_32),
.B(n_33),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_107),
.B1(n_106),
.B2(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_127),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_130),
.B(n_131),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_119),
.C(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_133),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_129),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_124),
.C(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_124),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_120),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_118),
.Y(n_140)
);


endmodule