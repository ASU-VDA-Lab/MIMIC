module fake_netlist_6_1316_n_796 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_796);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_796;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_758;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_631;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_49),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_24),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_0),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_45),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_33),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_78),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_10),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_35),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_18),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_109),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_40),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_32),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_80),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_68),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_84),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_127),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_41),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_42),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_76),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_108),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_29),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_34),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_30),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_97),
.Y(n_194)
);

BUFx2_ASAP7_75t_SL g195 ( 
.A(n_63),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_58),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_112),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_106),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_83),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_92),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_16),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_64),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_66),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_95),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_130),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_143),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_37),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_57),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_157),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_27),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_21),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_44),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_60),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_137),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_170),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_0),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_162),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_165),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_167),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_1),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_169),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_209),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_171),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_172),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_161),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_204),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_174),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_168),
.B(n_1),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_168),
.B(n_2),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_160),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_175),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_177),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_188),
.B(n_2),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_160),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_176),
.Y(n_259)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_193),
.B(n_213),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_179),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_221),
.B(n_215),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_180),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_166),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_225),
.B(n_205),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_211),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_231),
.B(n_181),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_241),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_237),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_208),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_219),
.B(n_179),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_228),
.B(n_182),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_236),
.B(n_179),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_218),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_240),
.B(n_207),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_223),
.B(n_183),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_223),
.B(n_185),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_235),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_189),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_238),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_R g314 ( 
.A(n_289),
.B(n_238),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_179),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_190),
.Y(n_316)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_280),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_273),
.B(n_229),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_195),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_307),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

NAND3x1_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_297),
.C(n_306),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_284),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_194),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_275),
.B(n_229),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_294),
.B(n_197),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_198),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g339 ( 
.A(n_294),
.B(n_295),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_294),
.B(n_200),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_307),
.Y(n_343)
);

INVx4_ASAP7_75t_SL g344 ( 
.A(n_268),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_265),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_297),
.B(n_202),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_280),
.B(n_206),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_265),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_265),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_265),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_280),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_3),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_296),
.B(n_20),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_276),
.B(n_233),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_276),
.B(n_233),
.C(n_4),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_279),
.Y(n_358)
);

NAND2xp33_ASAP7_75t_L g359 ( 
.A(n_295),
.B(n_3),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_304),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_264),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_270),
.B(n_22),
.Y(n_364)
);

AO21x2_ASAP7_75t_L g365 ( 
.A1(n_271),
.A2(n_85),
.B(n_156),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_286),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_262),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_299),
.B(n_291),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_266),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_291),
.B(n_4),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_266),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_281),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g373 ( 
.A1(n_281),
.A2(n_285),
.B1(n_301),
.B2(n_283),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_286),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_326),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

NAND2x1p5_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_290),
.Y(n_378)
);

AO22x2_ASAP7_75t_L g379 ( 
.A1(n_357),
.A2(n_301),
.B1(n_300),
.B2(n_298),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_307),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_309),
.Y(n_381)
);

OAI221xp5_ASAP7_75t_L g382 ( 
.A1(n_359),
.A2(n_292),
.B1(n_283),
.B2(n_290),
.C(n_282),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_339),
.A2(n_260),
.B1(n_290),
.B2(n_286),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_330),
.A2(n_260),
.B1(n_300),
.B2(n_298),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_346),
.B(n_302),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_309),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

NAND2x1p5_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_290),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_321),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_312),
.B(n_302),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_324),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_329),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_329),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_321),
.Y(n_400)
);

AO22x2_ASAP7_75t_L g401 ( 
.A1(n_356),
.A2(n_308),
.B1(n_6),
.B2(n_7),
.Y(n_401)
);

NAND2x1p5_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_292),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

AO22x2_ASAP7_75t_L g404 ( 
.A1(n_355),
.A2(n_308),
.B1(n_6),
.B2(n_7),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

NAND2x1p5_ASAP7_75t_L g406 ( 
.A(n_318),
.B(n_308),
.Y(n_406)
);

OR2x6_ASAP7_75t_SL g407 ( 
.A(n_354),
.B(n_308),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_351),
.Y(n_409)
);

AO22x2_ASAP7_75t_L g410 ( 
.A1(n_355),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_277),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

BUFx6f_ASAP7_75t_SL g414 ( 
.A(n_367),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_323),
.B(n_260),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_277),
.Y(n_417)
);

AO22x2_ASAP7_75t_L g418 ( 
.A1(n_327),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_316),
.B(n_260),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_268),
.Y(n_420)
);

AO22x2_ASAP7_75t_L g421 ( 
.A1(n_359),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_369),
.Y(n_422)
);

OAI221xp5_ASAP7_75t_L g423 ( 
.A1(n_316),
.A2(n_278),
.B1(n_286),
.B2(n_287),
.C(n_269),
.Y(n_423)
);

OAI221xp5_ASAP7_75t_L g424 ( 
.A1(n_338),
.A2(n_310),
.B1(n_346),
.B2(n_336),
.C(n_341),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

AO22x2_ASAP7_75t_L g426 ( 
.A1(n_373),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_325),
.B(n_278),
.Y(n_427)
);

AO22x2_ASAP7_75t_L g428 ( 
.A1(n_373),
.A2(n_332),
.B1(n_314),
.B2(n_364),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_338),
.B(n_286),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_L g430 ( 
.A(n_339),
.B(n_268),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_325),
.B(n_287),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

OAI221xp5_ASAP7_75t_L g433 ( 
.A1(n_310),
.A2(n_287),
.B1(n_269),
.B2(n_261),
.C(n_16),
.Y(n_433)
);

AO22x2_ASAP7_75t_L g434 ( 
.A1(n_314),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_320),
.Y(n_435)
);

AO22x2_ASAP7_75t_L g436 ( 
.A1(n_344),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_436)
);

NAND2x1p5_ASAP7_75t_L g437 ( 
.A(n_353),
.B(n_287),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_353),
.A2(n_287),
.B1(n_261),
.B2(n_96),
.Y(n_438)
);

AO22x2_ASAP7_75t_L g439 ( 
.A1(n_344),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_313),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_351),
.B(n_261),
.Y(n_441)
);

BUFx6f_ASAP7_75t_SL g442 ( 
.A(n_367),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g443 ( 
.A1(n_344),
.A2(n_19),
.B1(n_328),
.B2(n_347),
.Y(n_443)
);

AO22x2_ASAP7_75t_L g444 ( 
.A1(n_343),
.A2(n_261),
.B1(n_25),
.B2(n_26),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_411),
.B(n_361),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_411),
.B(n_361),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_384),
.B(n_320),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_385),
.B(n_320),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_409),
.B(n_343),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_415),
.B(n_320),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_417),
.B(n_317),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_380),
.B(n_365),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_417),
.B(n_375),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_376),
.B(n_317),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_377),
.B(n_317),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_386),
.B(n_317),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_388),
.B(n_391),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_392),
.B(n_366),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_402),
.B(n_366),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_414),
.B(n_365),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_393),
.B(n_395),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_408),
.B(n_311),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_378),
.B(n_311),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_389),
.B(n_374),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_394),
.B(n_319),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_427),
.B(n_374),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_406),
.B(n_339),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_427),
.B(n_335),
.Y(n_468)
);

NAND2x1p5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_441),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_442),
.B(n_339),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_315),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_407),
.B(n_348),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_431),
.B(n_335),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_419),
.B(n_335),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_383),
.B(n_335),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_413),
.B(n_422),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_425),
.B(n_396),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_397),
.B(n_345),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_398),
.B(n_315),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_399),
.B(n_345),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_403),
.B(n_345),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_405),
.B(n_345),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_412),
.B(n_349),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_416),
.B(n_350),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_SL g485 ( 
.A(n_438),
.B(n_315),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_SL g486 ( 
.A(n_404),
.B(n_315),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_SL g487 ( 
.A(n_404),
.B(n_315),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_379),
.B(n_23),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_379),
.B(n_28),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g490 ( 
.A(n_440),
.B(n_31),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_432),
.B(n_36),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_437),
.B(n_38),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_381),
.B(n_39),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_428),
.B(n_401),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_387),
.B(n_43),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_424),
.B(n_268),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_390),
.B(n_46),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_400),
.B(n_47),
.Y(n_498)
);

AO31x2_ASAP7_75t_L g499 ( 
.A1(n_496),
.A2(n_428),
.A3(n_382),
.B(n_433),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_475),
.A2(n_430),
.B(n_420),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_449),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_472),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_471),
.A2(n_435),
.B(n_423),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_444),
.B(n_439),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_461),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_465),
.Y(n_506)
);

AOI21x1_ASAP7_75t_SL g507 ( 
.A1(n_488),
.A2(n_443),
.B(n_421),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_479),
.A2(n_443),
.B(n_439),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_453),
.B(n_444),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_489),
.B(n_401),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_469),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_457),
.A2(n_410),
.B(n_421),
.C(n_418),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_477),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_450),
.A2(n_268),
.B(n_410),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_462),
.Y(n_515)
);

NOR2x1_ASAP7_75t_SL g516 ( 
.A(n_492),
.B(n_436),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_494),
.A2(n_426),
.B1(n_418),
.B2(n_436),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_469),
.B(n_426),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_470),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_448),
.B(n_434),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_447),
.A2(n_434),
.B1(n_50),
.B2(n_51),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_473),
.A2(n_268),
.B(n_52),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_452),
.A2(n_48),
.B(n_53),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_483),
.A2(n_54),
.B(n_55),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_446),
.Y(n_526)
);

A2O1A1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_485),
.A2(n_56),
.B(n_59),
.C(n_61),
.Y(n_527)
);

OA21x2_ASAP7_75t_L g528 ( 
.A1(n_484),
.A2(n_62),
.B(n_65),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_467),
.B(n_466),
.Y(n_529)
);

CKINVDCx8_ASAP7_75t_R g530 ( 
.A(n_486),
.Y(n_530)
);

OAI21x1_ASAP7_75t_SL g531 ( 
.A1(n_487),
.A2(n_67),
.B(n_69),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_468),
.A2(n_70),
.B(n_71),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_451),
.B(n_158),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_459),
.A2(n_72),
.B(n_73),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g535 ( 
.A1(n_478),
.A2(n_74),
.B(n_75),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_463),
.A2(n_77),
.B(n_79),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_476),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_490),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_497),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_458),
.B(n_82),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_480),
.A2(n_86),
.B(n_87),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_460),
.Y(n_542)
);

OA21x2_ASAP7_75t_L g543 ( 
.A1(n_524),
.A2(n_498),
.B(n_497),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_510),
.B(n_498),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_509),
.A2(n_491),
.B1(n_464),
.B2(n_495),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_500),
.A2(n_482),
.B(n_481),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_502),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_505),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_502),
.B(n_456),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_524),
.A2(n_493),
.B(n_455),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_511),
.B(n_454),
.Y(n_551)
);

AOI221xp5_ASAP7_75t_L g552 ( 
.A1(n_522),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.C(n_93),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_539),
.A2(n_94),
.B(n_98),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_506),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_529),
.B(n_99),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_503),
.A2(n_100),
.B(n_101),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_537),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_508),
.A2(n_102),
.B(n_103),
.Y(n_558)
);

OAI21x1_ASAP7_75t_SL g559 ( 
.A1(n_531),
.A2(n_104),
.B(n_107),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_504),
.B(n_110),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_502),
.B(n_155),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_513),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_515),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_530),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_512),
.B(n_115),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_499),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_525),
.A2(n_116),
.B(n_117),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_541),
.A2(n_118),
.B(n_119),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_536),
.A2(n_121),
.B(n_122),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_499),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_535),
.A2(n_507),
.B(n_534),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_520),
.B(n_123),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_499),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_528),
.Y(n_574)
);

O2A1O1Ixp33_ASAP7_75t_SL g575 ( 
.A1(n_527),
.A2(n_124),
.B(n_125),
.C(n_126),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_517),
.B(n_521),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_518),
.A2(n_542),
.B1(n_517),
.B2(n_520),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_538),
.A2(n_128),
.B(n_131),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_538),
.B(n_133),
.Y(n_579)
);

OAI21x1_ASAP7_75t_SL g580 ( 
.A1(n_516),
.A2(n_134),
.B(n_135),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_528),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_533),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_501),
.B(n_154),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_519),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_566),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_566),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_570),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_584),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_563),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_548),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_548),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_570),
.Y(n_592)
);

OA21x2_ASAP7_75t_L g593 ( 
.A1(n_573),
.A2(n_514),
.B(n_532),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_557),
.Y(n_594)
);

AOI31xp33_ASAP7_75t_L g595 ( 
.A1(n_552),
.A2(n_514),
.A3(n_540),
.B(n_523),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_557),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_556),
.A2(n_546),
.B(n_567),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_556),
.A2(n_526),
.B(n_520),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_569),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_562),
.Y(n_600)
);

NAND2x1p5_ASAP7_75t_L g601 ( 
.A(n_571),
.B(n_526),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_573),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_574),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_554),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_547),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_560),
.B(n_526),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_577),
.A2(n_136),
.B1(n_138),
.B2(n_142),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_572),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_544),
.B(n_151),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_558),
.Y(n_610)
);

OAI22xp33_ASAP7_75t_L g611 ( 
.A1(n_560),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_572),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_544),
.B(n_148),
.Y(n_613)
);

BUFx4f_ASAP7_75t_SL g614 ( 
.A(n_547),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_572),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_560),
.A2(n_565),
.B1(n_576),
.B2(n_582),
.Y(n_616)
);

AOI21x1_ASAP7_75t_L g617 ( 
.A1(n_574),
.A2(n_149),
.B(n_150),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_543),
.A2(n_582),
.B(n_553),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_576),
.B(n_584),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_546),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_558),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_581),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_560),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_551),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_549),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_551),
.B(n_579),
.Y(n_626)
);

OAI221xp5_ASAP7_75t_L g627 ( 
.A1(n_545),
.A2(n_555),
.B1(n_583),
.B2(n_564),
.C(n_575),
.Y(n_627)
);

O2A1O1Ixp5_ASAP7_75t_L g628 ( 
.A1(n_581),
.A2(n_561),
.B(n_551),
.C(n_580),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_581),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_558),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_569),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_568),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_578),
.B(n_543),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_578),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_543),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_550),
.B(n_580),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_559),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_609),
.B(n_550),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_615),
.B(n_559),
.Y(n_639)
);

CKINVDCx12_ASAP7_75t_R g640 ( 
.A(n_606),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_588),
.B(n_550),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_608),
.B(n_612),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_614),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_590),
.B(n_596),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_625),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_R g646 ( 
.A(n_623),
.B(n_619),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_R g647 ( 
.A(n_629),
.B(n_608),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_596),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_616),
.B(n_626),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_R g650 ( 
.A(n_623),
.B(n_606),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_626),
.B(n_608),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_591),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_600),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g654 ( 
.A(n_605),
.B(n_609),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_629),
.B(n_612),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_590),
.B(n_594),
.Y(n_656)
);

OR2x4_ASAP7_75t_L g657 ( 
.A(n_608),
.B(n_612),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_613),
.B(n_608),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_613),
.B(n_612),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_600),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_604),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_612),
.B(n_624),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_R g663 ( 
.A(n_606),
.B(n_626),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_618),
.B(n_585),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_589),
.B(n_611),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_606),
.B(n_598),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_585),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_598),
.B(n_601),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_601),
.B(n_637),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_R g670 ( 
.A(n_636),
.B(n_633),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_637),
.Y(n_671)
);

XOR2xp5_ASAP7_75t_L g672 ( 
.A(n_601),
.B(n_607),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_636),
.B(n_633),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_617),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_586),
.B(n_587),
.Y(n_675)
);

XOR2xp5_ASAP7_75t_L g676 ( 
.A(n_617),
.B(n_586),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_587),
.B(n_592),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_603),
.Y(n_678)
);

NAND2xp33_ASAP7_75t_R g679 ( 
.A(n_593),
.B(n_632),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_666),
.B(n_592),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_667),
.Y(n_681)
);

INVxp33_ASAP7_75t_L g682 ( 
.A(n_654),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_673),
.B(n_635),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_653),
.B(n_660),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_661),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_664),
.B(n_635),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_677),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_638),
.B(n_602),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_653),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_677),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_669),
.B(n_652),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_675),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_648),
.B(n_660),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_678),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_645),
.B(n_603),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_664),
.B(n_620),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_668),
.B(n_656),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_648),
.B(n_602),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_656),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_644),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_641),
.B(n_622),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_671),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_676),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_650),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_658),
.B(n_622),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_644),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_659),
.B(n_620),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_671),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_L g709 ( 
.A(n_665),
.B(n_627),
.C(n_595),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_674),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_643),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_681),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_683),
.B(n_649),
.Y(n_713)
);

AOI33xp33_ASAP7_75t_L g714 ( 
.A1(n_699),
.A2(n_639),
.A3(n_662),
.B1(n_621),
.B2(n_610),
.B3(n_646),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_683),
.B(n_651),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_680),
.B(n_670),
.Y(n_716)
);

AOI221xp5_ASAP7_75t_L g717 ( 
.A1(n_709),
.A2(n_703),
.B1(n_685),
.B2(n_695),
.C(n_699),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_681),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_689),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_706),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_697),
.Y(n_721)
);

AND4x1_ASAP7_75t_L g722 ( 
.A(n_701),
.B(n_628),
.C(n_640),
.D(n_655),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_693),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_680),
.B(n_691),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_680),
.B(n_670),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_697),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_691),
.B(n_639),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_693),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_724),
.B(n_701),
.Y(n_729)
);

NAND2x1p5_ASAP7_75t_L g730 ( 
.A(n_722),
.B(n_702),
.Y(n_730)
);

NAND2x1_ASAP7_75t_L g731 ( 
.A(n_716),
.B(n_702),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_718),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_724),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_721),
.B(n_686),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_720),
.B(n_719),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_719),
.B(n_682),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_712),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_716),
.B(n_704),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_718),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_738),
.B(n_726),
.Y(n_740)
);

NOR2x1_ASAP7_75t_L g741 ( 
.A(n_735),
.B(n_702),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_735),
.B(n_711),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_730),
.A2(n_717),
.B1(n_657),
.B2(n_736),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_739),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_730),
.A2(n_663),
.B1(n_725),
.B2(n_713),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_734),
.B(n_728),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_740),
.B(n_729),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_746),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_744),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_741),
.Y(n_750)
);

AOI222xp33_ASAP7_75t_L g751 ( 
.A1(n_748),
.A2(n_743),
.B1(n_742),
.B2(n_736),
.C1(n_713),
.C2(n_725),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_749),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_748),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_750),
.A2(n_745),
.B(n_731),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_751),
.B(n_747),
.Y(n_755)
);

OAI31xp33_ASAP7_75t_SL g756 ( 
.A1(n_754),
.A2(n_727),
.A3(n_715),
.B(n_733),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_753),
.B(n_737),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_757),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_755),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_756),
.Y(n_760)
);

INVx5_ASAP7_75t_L g761 ( 
.A(n_757),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_759),
.B(n_752),
.C(n_714),
.Y(n_762)
);

NAND4xp25_ASAP7_75t_L g763 ( 
.A(n_758),
.B(n_684),
.C(n_710),
.D(n_642),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_SL g764 ( 
.A(n_761),
.B(n_760),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_761),
.Y(n_765)
);

OAI221xp5_ASAP7_75t_L g766 ( 
.A1(n_759),
.A2(n_708),
.B1(n_732),
.B2(n_672),
.C(n_723),
.Y(n_766)
);

NAND5xp2_ASAP7_75t_L g767 ( 
.A(n_764),
.B(n_710),
.C(n_727),
.D(n_715),
.E(n_705),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_765),
.B(n_708),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_SL g769 ( 
.A(n_762),
.B(n_647),
.C(n_690),
.Y(n_769)
);

AOI221xp5_ASAP7_75t_L g770 ( 
.A1(n_766),
.A2(n_687),
.B1(n_690),
.B2(n_692),
.C(n_662),
.Y(n_770)
);

AOI221x1_ASAP7_75t_L g771 ( 
.A1(n_763),
.A2(n_687),
.B1(n_694),
.B2(n_692),
.C(n_634),
.Y(n_771)
);

NAND4xp25_ASAP7_75t_L g772 ( 
.A(n_764),
.B(n_642),
.C(n_705),
.D(n_707),
.Y(n_772)
);

NAND4xp75_ASAP7_75t_L g773 ( 
.A(n_768),
.B(n_698),
.C(n_688),
.D(n_707),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_771),
.B(n_688),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_769),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_772),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_767),
.B(n_694),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_SL g778 ( 
.A(n_775),
.B(n_770),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_776),
.B(n_777),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_777),
.B(n_700),
.C(n_696),
.Y(n_780)
);

AOI222xp33_ASAP7_75t_L g781 ( 
.A1(n_778),
.A2(n_774),
.B1(n_773),
.B2(n_674),
.C1(n_630),
.C2(n_634),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_779),
.B(n_700),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_780),
.A2(n_657),
.B1(n_698),
.B2(n_674),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_782),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_781),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_783),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_782),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_785),
.A2(n_631),
.B(n_599),
.Y(n_788)
);

AOI22x1_ASAP7_75t_L g789 ( 
.A1(n_786),
.A2(n_696),
.B1(n_631),
.B2(n_686),
.Y(n_789)
);

AOI31xp33_ASAP7_75t_L g790 ( 
.A1(n_788),
.A2(n_787),
.A3(n_784),
.B(n_610),
.Y(n_790)
);

AOI31xp33_ASAP7_75t_L g791 ( 
.A1(n_789),
.A2(n_621),
.A3(n_679),
.B(n_630),
.Y(n_791)
);

XOR2xp5_ASAP7_75t_L g792 ( 
.A(n_790),
.B(n_593),
.Y(n_792)
);

OA21x2_ASAP7_75t_L g793 ( 
.A1(n_792),
.A2(n_791),
.B(n_597),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_793),
.Y(n_794)
);

AOI221xp5_ASAP7_75t_L g795 ( 
.A1(n_794),
.A2(n_599),
.B1(n_632),
.B2(n_630),
.C(n_679),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_795),
.A2(n_599),
.B1(n_632),
.B2(n_593),
.Y(n_796)
);


endmodule