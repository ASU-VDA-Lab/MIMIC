module fake_jpeg_12261_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_16),
.B1(n_38),
.B2(n_36),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_54),
.B1(n_50),
.B2(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_50),
.B1(n_61),
.B2(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_49),
.B1(n_44),
.B2(n_55),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_61),
.B1(n_66),
.B2(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_80),
.B1(n_84),
.B2(n_62),
.Y(n_97)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_85),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_104),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_59),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_94),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_56),
.B1(n_46),
.B2(n_45),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_97),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_103),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_58),
.B(n_48),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_17),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_102),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_58),
.B1(n_48),
.B2(n_15),
.Y(n_101)
);

NAND2x1p5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_58),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_1),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_22),
.C(n_40),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_111),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_2),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_110),
.C(n_5),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_120),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_2),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_14),
.B1(n_34),
.B2(n_31),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_108),
.B1(n_116),
.B2(n_106),
.Y(n_133)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_35),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_93),
.B(n_3),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_4),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_133),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_96),
.C(n_23),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_128),
.C(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_5),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_28),
.C(n_27),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_136),
.A2(n_107),
.B(n_25),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_112),
.B1(n_122),
.B2(n_124),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_107),
.B(n_7),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_135),
.B1(n_129),
.B2(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_130),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_125),
.C(n_24),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_146),
.B(n_143),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_6),
.B(n_7),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_150),
.B(n_6),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_8),
.Y(n_152)
);


endmodule