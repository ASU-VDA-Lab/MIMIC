module fake_jpeg_20169_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_19),
.B1(n_20),
.B2(n_28),
.Y(n_71)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_30),
.B1(n_27),
.B2(n_31),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_23),
.B1(n_34),
.B2(n_29),
.Y(n_82)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_30),
.B1(n_27),
.B2(n_37),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_19),
.B1(n_32),
.B2(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_57),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_79),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_39),
.B(n_16),
.C(n_32),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_21),
.B1(n_38),
.B2(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_21),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_38),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_71),
.B1(n_74),
.B2(n_45),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_17),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_17),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_29),
.Y(n_79)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_83),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_84),
.B1(n_0),
.B2(n_1),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_34),
.B1(n_24),
.B2(n_2),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_73),
.Y(n_104)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_91),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_60),
.B1(n_67),
.B2(n_69),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_96),
.B1(n_108),
.B2(n_64),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_44),
.B1(n_24),
.B2(n_3),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_89),
.B1(n_92),
.B2(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_24),
.C(n_15),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_79),
.C(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_59),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_3),
.C(n_4),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_81),
.B(n_59),
.C(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_104),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_89),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_96),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_107),
.B1(n_80),
.B2(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_66),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_119),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_93),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_97),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_86),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_133),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_66),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_83),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_99),
.B1(n_61),
.B2(n_7),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_64),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_75),
.B1(n_68),
.B2(n_6),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_105),
.B(n_98),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_142),
.B(n_147),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_103),
.B(n_100),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_145),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_103),
.B1(n_75),
.B2(n_107),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_115),
.B1(n_126),
.B2(n_119),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_132),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_88),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_155),
.C(n_124),
.Y(n_165)
);

AOI21x1_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_91),
.B(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_123),
.B(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_128),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_152),
.B1(n_117),
.B2(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_99),
.B1(n_61),
.B2(n_7),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_4),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_134),
.B(n_118),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_61),
.C(n_7),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_161),
.B1(n_171),
.B2(n_174),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_162),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_172),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_167),
.B(n_168),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_130),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_150),
.B(n_135),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_173),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_133),
.B(n_111),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_171),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_133),
.C(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_133),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_153),
.A2(n_116),
.B(n_115),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_13),
.C(n_8),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_187),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_184),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_146),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_158),
.B1(n_170),
.B2(n_169),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_149),
.B1(n_152),
.B2(n_139),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_140),
.B1(n_176),
.B2(n_159),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_165),
.C(n_164),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_196),
.C(n_201),
.Y(n_206)
);

BUFx12_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_190),
.B(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

XOR2x2_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_164),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_181),
.B1(n_182),
.B2(n_138),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_139),
.C(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_167),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_183),
.B1(n_188),
.B2(n_185),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_160),
.C(n_143),
.Y(n_201)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_209),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_201),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_175),
.B(n_140),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_200),
.C(n_191),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_212),
.Y(n_220)
);

AOI211xp5_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_194),
.B(n_192),
.C(n_196),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_200),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_217),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_180),
.C(n_192),
.Y(n_217)
);

AOI211xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_204),
.B(n_209),
.C(n_205),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_218),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_210),
.B1(n_207),
.B2(n_9),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_225),
.Y(n_227)
);

OAI22x1_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_212),
.B1(n_216),
.B2(n_9),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_220),
.C(n_219),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_219),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_227),
.C(n_10),
.Y(n_229)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_5),
.B(n_12),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_5),
.Y(n_231)
);


endmodule