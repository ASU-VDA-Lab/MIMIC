module fake_jpeg_14331_n_474 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_474);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_474;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_48),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_87),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_75),
.Y(n_140)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_79),
.Y(n_142)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_24),
.B(n_8),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_18),
.B(n_8),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_89),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_46),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_91),
.Y(n_108)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_18),
.B(n_8),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_95),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_16),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_52),
.A2(n_47),
.B1(n_46),
.B2(n_43),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_102),
.A2(n_115),
.B1(n_119),
.B2(n_133),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_47),
.B1(n_46),
.B2(n_37),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_104),
.A2(n_40),
.B1(n_35),
.B2(n_42),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_117),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_59),
.A2(n_47),
.B1(n_35),
.B2(n_32),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_34),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_47),
.B1(n_16),
.B2(n_43),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_44),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_58),
.B(n_44),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_61),
.A2(n_19),
.B1(n_22),
.B2(n_42),
.Y(n_133)
);

NAND2x1_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_43),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_135),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_57),
.A2(n_45),
.B1(n_36),
.B2(n_34),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_50),
.B(n_22),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_145),
.B(n_22),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_158),
.Y(n_201)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_65),
.B1(n_55),
.B2(n_73),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_96),
.Y(n_152)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_96),
.A2(n_91),
.B1(n_71),
.B2(n_40),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_154),
.B(n_195),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_62),
.B1(n_86),
.B2(n_82),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_155),
.A2(n_165),
.B1(n_138),
.B2(n_124),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_122),
.A2(n_67),
.B1(n_36),
.B2(n_31),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_111),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_108),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_182),
.Y(n_213)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_49),
.Y(n_164)
);

NAND2x1_ASAP7_75t_L g232 ( 
.A(n_164),
.B(n_166),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_49),
.Y(n_166)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_23),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_170),
.B(n_171),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_116),
.B(n_23),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_174),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_112),
.A2(n_33),
.B(n_36),
.C(n_34),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_185),
.B(n_31),
.C(n_27),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_87),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_140),
.C(n_142),
.Y(n_204)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_97),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_191),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_104),
.A2(n_93),
.B1(n_70),
.B2(n_81),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_183),
.B1(n_189),
.B2(n_102),
.Y(n_203)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_105),
.B(n_19),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_188),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_23),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_135),
.A2(n_66),
.B1(n_77),
.B2(n_63),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_110),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_187),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_98),
.B(n_76),
.CI(n_87),
.CON(n_185),
.SN(n_185)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_129),
.B(n_19),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_41),
.Y(n_225)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_97),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_118),
.Y(n_202)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_21),
.B1(n_31),
.B2(n_33),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_42),
.B(n_41),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_121),
.B(n_40),
.Y(n_195)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g270 ( 
.A1(n_203),
.A2(n_106),
.B1(n_168),
.B2(n_163),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_211),
.C(n_230),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_148),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_195),
.Y(n_250)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_154),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_140),
.C(n_142),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_212),
.A2(n_21),
.B(n_27),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_152),
.B1(n_165),
.B2(n_181),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_225),
.B(n_234),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_103),
.B1(n_99),
.B2(n_137),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_233),
.B1(n_152),
.B2(n_176),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_166),
.B(n_141),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_149),
.B(n_100),
.C(n_72),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_235),
.C(n_169),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_137),
.B1(n_132),
.B2(n_107),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_158),
.B(n_100),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_169),
.B(n_139),
.C(n_136),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_153),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_240),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_237),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_239),
.B(n_250),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_249),
.B1(n_257),
.B2(n_260),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_164),
.B1(n_161),
.B2(n_184),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_199),
.A2(n_164),
.B1(n_192),
.B2(n_175),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_246),
.A2(n_220),
.B(n_212),
.Y(n_273)
);

AO21x2_ASAP7_75t_L g247 ( 
.A1(n_207),
.A2(n_154),
.B(n_180),
.Y(n_247)
);

INVxp33_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_248),
.B(n_254),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_203),
.A2(n_195),
.B1(n_157),
.B2(n_107),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_252),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_235),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_259),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_191),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_215),
.A2(n_177),
.B(n_185),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_255),
.A2(n_210),
.B(n_228),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_201),
.B(n_178),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_256),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_215),
.A2(n_127),
.B1(n_136),
.B2(n_139),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_216),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_127),
.B1(n_143),
.B2(n_176),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_202),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_263),
.Y(n_286)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_209),
.B(n_173),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_200),
.A2(n_193),
.B1(n_185),
.B2(n_186),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_270),
.B1(n_265),
.B2(n_260),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_200),
.A2(n_143),
.B1(n_118),
.B2(n_167),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_265),
.A2(n_218),
.B1(n_168),
.B2(n_162),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_177),
.C(n_160),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_239),
.C(n_238),
.Y(n_279)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_232),
.B(n_230),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_213),
.B(n_150),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_271),
.Y(n_277)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_272),
.A2(n_219),
.B1(n_229),
.B2(n_218),
.Y(n_299)
);

A2O1A1O1Ixp25_ASAP7_75t_L g312 ( 
.A1(n_273),
.A2(n_301),
.B(n_294),
.C(n_276),
.D(n_291),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_249),
.A2(n_206),
.B1(n_204),
.B2(n_231),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_275),
.A2(n_276),
.B(n_294),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_246),
.A2(n_206),
.B(n_227),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_243),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_278),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_247),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_237),
.A2(n_232),
.B1(n_211),
.B2(n_222),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_281),
.A2(n_292),
.B1(n_257),
.B2(n_247),
.Y(n_324)
);

OA22x2_ASAP7_75t_L g334 ( 
.A1(n_288),
.A2(n_304),
.B1(n_247),
.B2(n_196),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_262),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_251),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_208),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_295),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_247),
.A2(n_222),
.B1(n_226),
.B2(n_208),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_246),
.A2(n_226),
.B(n_210),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_241),
.B(n_221),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_263),
.A2(n_238),
.B(n_245),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_297),
.B(n_305),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_299),
.A2(n_229),
.B1(n_214),
.B2(n_267),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_221),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_302),
.C(n_266),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_250),
.B(n_223),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_244),
.A2(n_223),
.B(n_229),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_241),
.B(n_228),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_252),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_308),
.B(n_300),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_266),
.C(n_255),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_315),
.C(n_326),
.Y(n_347)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_312),
.A2(n_331),
.B(n_280),
.Y(n_342)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_287),
.Y(n_314)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_240),
.C(n_259),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_278),
.A2(n_275),
.B1(n_284),
.B2(n_282),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_317),
.A2(n_336),
.B1(n_301),
.B2(n_282),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_258),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_322),
.C(n_323),
.Y(n_344)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_321),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_274),
.B(n_258),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_277),
.B(n_214),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_324),
.A2(n_288),
.B1(n_304),
.B2(n_307),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_325),
.B(n_328),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_285),
.B(n_268),
.C(n_242),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_302),
.C(n_305),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_295),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_329),
.A2(n_304),
.B1(n_299),
.B2(n_303),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_289),
.A2(n_292),
.B1(n_281),
.B2(n_286),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_330),
.A2(n_324),
.B1(n_331),
.B2(n_320),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_289),
.A2(n_247),
.B1(n_269),
.B2(n_272),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_274),
.B(n_196),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_333),
.B(n_290),
.Y(n_366)
);

INVx3_ASAP7_75t_SL g354 ( 
.A(n_334),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_286),
.B(n_272),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_335),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_275),
.A2(n_196),
.B1(n_162),
.B2(n_120),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_338),
.Y(n_363)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_340),
.A2(n_351),
.B1(n_355),
.B2(n_330),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_285),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_348),
.Y(n_370)
);

AOI21xp33_ASAP7_75t_L g350 ( 
.A1(n_319),
.A2(n_301),
.B(n_293),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_336),
.B1(n_328),
.B2(n_309),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_339),
.A2(n_273),
.B(n_293),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_300),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_357),
.C(n_358),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_309),
.A2(n_307),
.B1(n_302),
.B2(n_284),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_297),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_360),
.A2(n_362),
.B1(n_367),
.B2(n_334),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_321),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_366),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_296),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_364),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_303),
.C(n_298),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_332),
.C(n_298),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_369),
.A2(n_356),
.B1(n_343),
.B2(n_358),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_371),
.A2(n_384),
.B1(n_386),
.B2(n_389),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_313),
.Y(n_372)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_359),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_378),
.Y(n_406)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_363),
.Y(n_376)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_354),
.A2(n_313),
.B1(n_325),
.B2(n_314),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_359),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_379),
.B(n_383),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_352),
.A2(n_312),
.B(n_339),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_21),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_354),
.A2(n_335),
.B1(n_316),
.B2(n_337),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_354),
.A2(n_319),
.B1(n_334),
.B2(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_368),
.Y(n_385)
);

AO221x1_ASAP7_75t_L g411 ( 
.A1(n_385),
.A2(n_390),
.B1(n_0),
.B2(n_1),
.C(n_2),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_362),
.A2(n_341),
.B1(n_343),
.B2(n_367),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_392),
.C(n_348),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_334),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_388),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_341),
.A2(n_75),
.B1(n_35),
.B2(n_41),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_174),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_347),
.B(n_174),
.C(n_33),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_SL g417 ( 
.A(n_394),
.B(n_404),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_347),
.C(n_346),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_405),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_370),
.B(n_357),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_370),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_400),
.A2(n_408),
.B1(n_409),
.B2(n_389),
.Y(n_418)
);

BUFx12f_ASAP7_75t_SL g401 ( 
.A(n_380),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_391),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_377),
.A2(n_351),
.B(n_355),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g414 ( 
.A(n_402),
.B(n_384),
.Y(n_414)
);

OAI322xp33_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_344),
.A3(n_353),
.B1(n_342),
.B2(n_365),
.C1(n_368),
.C2(n_340),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_174),
.C(n_27),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_372),
.C(n_385),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_369),
.A2(n_37),
.B1(n_32),
.B2(n_2),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_379),
.A2(n_37),
.B1(n_32),
.B2(n_2),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_0),
.C(n_1),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_0),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_411),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_403),
.A2(n_373),
.B1(n_377),
.B2(n_388),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_412),
.A2(n_406),
.B1(n_398),
.B2(n_393),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_419),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_414),
.A2(n_403),
.B1(n_406),
.B2(n_394),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_373),
.C(n_392),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_416),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_395),
.B(n_376),
.Y(n_416)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_418),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_421),
.A2(n_427),
.B(n_395),
.Y(n_430)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_401),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_424),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_R g425 ( 
.A(n_399),
.B(n_374),
.C(n_381),
.Y(n_425)
);

INVx11_ASAP7_75t_L g428 ( 
.A(n_425),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_386),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_426),
.B(n_407),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_402),
.A2(n_371),
.B(n_9),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_425),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_429),
.B(n_430),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_414),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_436),
.Y(n_453)
);

OAI21xp33_ASAP7_75t_L g452 ( 
.A1(n_434),
.A2(n_6),
.B(n_12),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_397),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_423),
.B(n_405),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_437),
.B(n_438),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_412),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_427),
.A2(n_408),
.B1(n_409),
.B2(n_410),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_440),
.B(n_6),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_439),
.B(n_420),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_443),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_435),
.C(n_434),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_436),
.B(n_417),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_448),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_445),
.A2(n_446),
.B1(n_450),
.B2(n_433),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_428),
.B(n_419),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_428),
.B(n_414),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_431),
.A2(n_413),
.B(n_6),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_449),
.A2(n_452),
.B(n_5),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_451),
.B(n_441),
.Y(n_454)
);

NAND3xp33_ASAP7_75t_SL g463 ( 
.A(n_454),
.B(n_461),
.C(n_455),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_430),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_457),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_445),
.B(n_433),
.C(n_440),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_460),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_5),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_459),
.B(n_446),
.C(n_452),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_463),
.Y(n_469)
);

OAI31xp67_ASAP7_75t_L g466 ( 
.A1(n_454),
.A2(n_5),
.A3(n_11),
.B(n_2),
.Y(n_466)
);

A2O1A1O1Ixp25_ASAP7_75t_L g468 ( 
.A1(n_466),
.A2(n_3),
.B(n_10),
.C(n_11),
.D(n_15),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_457),
.C(n_3),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_467),
.A2(n_468),
.B(n_0),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_464),
.C(n_10),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_470),
.A2(n_471),
.B(n_1),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_472),
.A2(n_11),
.B(n_1),
.Y(n_473)
);

HAxp5_ASAP7_75t_SL g474 ( 
.A(n_473),
.B(n_11),
.CON(n_474),
.SN(n_474)
);


endmodule