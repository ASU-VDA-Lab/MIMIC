module real_jpeg_2087_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_28),
.B1(n_32),
.B2(n_37),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_1),
.A2(n_28),
.B1(n_50),
.B2(n_51),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_1),
.A2(n_28),
.B1(n_63),
.B2(n_67),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_2),
.A2(n_63),
.B1(n_67),
.B2(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_2),
.A2(n_32),
.B1(n_37),
.B2(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_3),
.B(n_25),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_3),
.B(n_166),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_3),
.A2(n_37),
.B(n_47),
.C(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_3),
.B(n_49),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_3),
.A2(n_32),
.B1(n_37),
.B2(n_216),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_3),
.B(n_63),
.C(n_66),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_216),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_3),
.B(n_88),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_3),
.B(n_61),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_5),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_5),
.A2(n_32),
.B1(n_37),
.B2(n_98),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_98),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_5),
.A2(n_63),
.B1(n_67),
.B2(n_98),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_6),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_6),
.A2(n_32),
.B1(n_37),
.B2(n_137),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_137),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_6),
.A2(n_63),
.B1(n_67),
.B2(n_137),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_32),
.B1(n_37),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_58),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_7),
.A2(n_58),
.B1(n_63),
.B2(n_67),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_9),
.A2(n_32),
.B1(n_37),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_55),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_9),
.A2(n_55),
.B1(n_63),
.B2(n_67),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_14),
.A2(n_32),
.B1(n_37),
.B2(n_41),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_14),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_14),
.A2(n_41),
.B1(n_63),
.B2(n_67),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_15),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_15),
.A2(n_32),
.B1(n_37),
.B2(n_165),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_15),
.A2(n_50),
.B1(n_51),
.B2(n_165),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_15),
.A2(n_63),
.B1(n_67),
.B2(n_165),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_112),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_110),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_99),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_20),
.B(n_99),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_80),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_21),
.B(n_74),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_42),
.B2(n_73),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_22),
.A2(n_23),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_23),
.B(n_43),
.C(n_60),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_31),
.B2(n_40),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_24),
.A2(n_31),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_26),
.B1(n_35),
.B2(n_38),
.Y(n_39)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_26),
.A2(n_35),
.A3(n_37),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_26),
.A2(n_29),
.B(n_216),
.C(n_225),
.Y(n_224)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_29),
.A2(n_31),
.B1(n_40),
.B2(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_29),
.A2(n_135),
.B(n_138),
.Y(n_134)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_30),
.A2(n_136),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_31),
.B(n_97),
.Y(n_139)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_31),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_31),
.A2(n_95),
.B(n_180),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_32),
.B(n_38),
.Y(n_188)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_47),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_59),
.B2(n_60),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_54),
.B1(n_56),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_45),
.A2(n_56),
.B1(n_57),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_45),
.A2(n_56),
.B1(n_76),
.B2(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_45),
.A2(n_182),
.B(n_184),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_45),
.A2(n_184),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_46),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_46),
.A2(n_49),
.B1(n_183),
.B2(n_200),
.Y(n_228)
);

AO22x2_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_49)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_49),
.B(n_162),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_51),
.B1(n_65),
.B2(n_66),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_50),
.A2(n_53),
.B(n_216),
.Y(n_215)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_51),
.B(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_56),
.A2(n_133),
.B(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_56),
.A2(n_161),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_60),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_68),
.B(n_70),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_61),
.A2(n_68),
.B1(n_93),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_61),
.A2(n_68),
.B1(n_131),
.B2(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_61),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_71),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_78),
.B1(n_79),
.B2(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_62),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_62),
.A2(n_232),
.B(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_62),
.A2(n_78),
.B1(n_209),
.B2(n_243),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_63),
.B(n_272),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_68),
.A2(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_68),
.B(n_212),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_74),
.A2(n_75),
.B(n_77),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_78),
.A2(n_211),
.B(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B(n_94),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_82),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_91),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_84),
.B1(n_94),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_83),
.A2(n_84),
.B1(n_91),
.B2(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_88),
.B(n_89),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_88),
.B1(n_128),
.B2(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_85),
.A2(n_216),
.B(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_86),
.A2(n_87),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_86),
.A2(n_87),
.B1(n_191),
.B2(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_86),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_86),
.A2(n_247),
.B(n_248),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_86),
.A2(n_87),
.B1(n_247),
.B2(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_87),
.A2(n_206),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_87),
.B(n_220),
.Y(n_249)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_88),
.A2(n_219),
.B(n_276),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_91),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_140),
.B(n_313),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_114),
.B(n_116),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.C(n_123),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_132),
.C(n_134),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_125),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_134),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_139),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_167),
.B(n_312),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_143),
.B(n_146),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.C(n_163),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_154),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_155),
.B(n_157),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_156),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

OAI21x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_193),
.B(n_311),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_169),
.B(n_171),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_178),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_172),
.B(n_176),
.Y(n_296)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_178),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_185),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_179),
.B(n_181),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_185),
.B(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_186),
.A2(n_189),
.B1(n_190),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI31xp33_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_293),
.A3(n_303),
.B(n_308),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_237),
.B(n_292),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_221),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_196),
.B(n_221),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_207),
.C(n_213),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_197),
.B(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_202),
.C(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_207),
.B(n_213),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_217),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_233),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_222),
.B(n_234),
.C(n_236),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_223),
.B(n_228),
.C(n_229),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_287),
.B(n_291),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_256),
.B(n_286),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_250),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_240),
.B(n_250),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_246),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_255),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_254),
.C(n_255),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_268),
.B(n_285),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_264),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_264),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_279),
.B(n_284),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_274),
.B(n_278),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_277),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_282),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_297),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_307),
.Y(n_309)
);


endmodule