module fake_jpeg_6415_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx24_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_3),
.B(n_0),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_12),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_12),
.B1(n_7),
.B2(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_17),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_0),
.Y(n_16)
);

AO21x1_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_11),
.B(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_19),
.Y(n_25)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_21),
.B(n_28),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_4),
.B1(n_9),
.B2(n_16),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_16),
.C(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_21),
.B1(n_20),
.B2(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NAND4xp25_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_24),
.C(n_28),
.D(n_20),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_38),
.B(n_34),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_37),
.B(n_36),
.C(n_42),
.Y(n_43)
);

AOI32xp33_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_44),
.A3(n_22),
.B1(n_41),
.B2(n_30),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_29),
.B(n_18),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_R g47 ( 
.A(n_46),
.B(n_19),
.Y(n_47)
);


endmodule