module fake_netlist_5_751_n_1946 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1946);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1946;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_192;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_46),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_126),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_153),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_53),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_184),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_91),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_85),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_45),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_27),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_77),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_129),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_4),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_39),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_1),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_31),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_28),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_8),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_101),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_15),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_17),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_100),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_39),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_119),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_161),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_61),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_159),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_109),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_10),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_17),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_41),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_58),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_55),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_81),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_40),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_54),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_124),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_105),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_136),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_45),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_78),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_36),
.Y(n_245)
);

BUFx8_ASAP7_75t_SL g246 ( 
.A(n_139),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_18),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_165),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_71),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_154),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_93),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_148),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_57),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_64),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_67),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_96),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_75),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_177),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_110),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_88),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_170),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_2),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_82),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_13),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_44),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_157),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_160),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_121),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_12),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_103),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_34),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_54),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_186),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_174),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_125),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_46),
.Y(n_276)
);

BUFx8_ASAP7_75t_SL g277 ( 
.A(n_72),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_123),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_94),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_40),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_144),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_65),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_112),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_21),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_27),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_117),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_9),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_52),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_26),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_116),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_49),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_149),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_92),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_5),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_135),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_18),
.Y(n_296)
);

BUFx8_ASAP7_75t_SL g297 ( 
.A(n_95),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_34),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_80),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_5),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_86),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_138),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_180),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_26),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_127),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_63),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_120),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_147),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_179),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_104),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_143),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_21),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_146),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_58),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_131),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_150),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_83),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_108),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_3),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_32),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_66),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_6),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_69),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_158),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_97),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_140),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_189),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_166),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_115),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_8),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_141),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_98),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_169),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_74),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_152),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_137),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_79),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_76),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_173),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_52),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_24),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_182),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_156),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_33),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_57),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_128),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_4),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_11),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_183),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_118),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_23),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_41),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_1),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_106),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_19),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_44),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_178),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_107),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_22),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_188),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_35),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_32),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_19),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_2),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_60),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_35),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_167),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_23),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_0),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_30),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_16),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_175),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_99),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_33),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_90),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_53),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_51),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_10),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_56),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_246),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_256),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_288),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_277),
.Y(n_384)
);

INVxp33_ASAP7_75t_SL g385 ( 
.A(n_192),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_297),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_215),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_236),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_239),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_232),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_240),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_215),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_204),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_380),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_379),
.Y(n_396)
);

INVxp33_ASAP7_75t_SL g397 ( 
.A(n_192),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_241),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_272),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_228),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_213),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_230),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_245),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_242),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_303),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_194),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_196),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_244),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_196),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_194),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_264),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_269),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_249),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_248),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_250),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_271),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_280),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_299),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_263),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_284),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_365),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_294),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_281),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_251),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_339),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_344),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_371),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_298),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_252),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_347),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_300),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_321),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_299),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_342),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_255),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_370),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_258),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_201),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_330),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_362),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_259),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_267),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_275),
.Y(n_448)
);

INVxp33_ASAP7_75t_SL g449 ( 
.A(n_201),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_275),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_283),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_283),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_217),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_292),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_205),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_292),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_310),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_203),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_203),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_310),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_292),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_191),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_200),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_202),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_214),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_219),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_366),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_272),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_268),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_274),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_278),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_221),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_227),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_282),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_256),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_382),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_475),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_475),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_330),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_382),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_382),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_422),
.B(n_205),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_383),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_403),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_403),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_381),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_456),
.B(n_193),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_406),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_448),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_393),
.A2(n_315),
.B1(n_323),
.B2(n_262),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_444),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_450),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_422),
.B(n_205),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_450),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_451),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_452),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_452),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_453),
.A2(n_369),
.B1(n_364),
.B2(n_253),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_461),
.B(n_229),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_390),
.A2(n_352),
.B1(n_375),
.B2(n_207),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_444),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_457),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_457),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_388),
.B(n_220),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_399),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_460),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_460),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_387),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_396),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_387),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_401),
.A2(n_420),
.B1(n_424),
.B2(n_415),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g518 ( 
.A(n_441),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_392),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_458),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_392),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_468),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_396),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_389),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_394),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_394),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_400),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_402),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_462),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_426),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_427),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_462),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_L g534 ( 
.A(n_391),
.B(n_398),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_402),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_412),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_463),
.B(n_235),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_463),
.B(n_254),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_464),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_412),
.Y(n_540)
);

BUFx6f_ASAP7_75t_SL g541 ( 
.A(n_455),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_428),
.B(n_257),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_419),
.B(n_193),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_464),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_407),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_407),
.B(n_257),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_404),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_431),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_466),
.B(n_195),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_467),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_466),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_472),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_533),
.Y(n_555)
);

NOR2x1p5_ASAP7_75t_L g556 ( 
.A(n_524),
.B(n_384),
.Y(n_556)
);

AOI21x1_ASAP7_75t_L g557 ( 
.A1(n_481),
.A2(n_473),
.B(n_472),
.Y(n_557)
);

INVxp67_ASAP7_75t_SL g558 ( 
.A(n_546),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_546),
.B(n_407),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_547),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_547),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_486),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_428),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_533),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_486),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_480),
.B(n_409),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_505),
.A2(n_405),
.B(n_302),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_486),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_480),
.B(n_414),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_476),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_546),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_505),
.B(n_256),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_505),
.B(n_473),
.C(n_417),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_486),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_507),
.B(n_416),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_507),
.B(n_425),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_476),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_476),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_507),
.B(n_430),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_533),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_533),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_533),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_533),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_486),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_533),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_531),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_477),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_476),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_477),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_480),
.B(n_411),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_505),
.B(n_417),
.C(n_413),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_480),
.B(n_438),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_545),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_545),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_477),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_478),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_545),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_549),
.B(n_440),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_530),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_478),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_497),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_478),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_484),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_518),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_490),
.B(n_441),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_490),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_481),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_516),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_537),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_543),
.B(n_446),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_497),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_530),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_543),
.B(n_447),
.Y(n_617)
);

NAND2x1p5_ASAP7_75t_L g618 ( 
.A(n_537),
.B(n_260),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_532),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_537),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_481),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_537),
.A2(n_408),
.B1(n_410),
.B2(n_385),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_516),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_538),
.B(n_418),
.C(n_413),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_530),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_482),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_516),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_520),
.B(n_471),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_516),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_491),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_516),
.Y(n_632)
);

INVxp67_ASAP7_75t_SL g633 ( 
.A(n_482),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_539),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_520),
.B(n_397),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_516),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_519),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_491),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_483),
.B(n_449),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_539),
.Y(n_640)
);

NOR2x1p5_ASAP7_75t_L g641 ( 
.A(n_551),
.B(n_386),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_482),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_539),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_544),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_519),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_497),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_497),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_498),
.B(n_470),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_544),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_519),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_551),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_519),
.Y(n_652)
);

INVx11_ASAP7_75t_L g653 ( 
.A(n_489),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_544),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_485),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_519),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_511),
.B(n_474),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_496),
.B(n_411),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_511),
.B(n_455),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_534),
.B(n_459),
.Y(n_660)
);

CKINVDCx11_ASAP7_75t_R g661 ( 
.A(n_550),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_519),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_497),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_519),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_521),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_521),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_496),
.B(n_411),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_497),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_548),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_496),
.B(n_434),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_496),
.B(n_538),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_496),
.B(n_434),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_522),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_504),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_521),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_496),
.B(n_538),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_522),
.B(n_444),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_506),
.B(n_444),
.Y(n_678)
);

OAI21xp33_ASAP7_75t_SL g679 ( 
.A1(n_542),
.A2(n_445),
.B(n_443),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_538),
.A2(n_434),
.B1(n_279),
.B2(n_359),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_504),
.A2(n_233),
.B1(n_378),
.B2(n_375),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_552),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_521),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_548),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_548),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_515),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_506),
.B(n_257),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_553),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_521),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_553),
.A2(n_256),
.B1(n_261),
.B2(n_350),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_496),
.B(n_305),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_541),
.B(n_443),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_521),
.Y(n_693)
);

AND2x6_ASAP7_75t_L g694 ( 
.A(n_553),
.B(n_256),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_521),
.Y(n_695)
);

AND2x2_ASAP7_75t_SL g696 ( 
.A(n_494),
.B(n_261),
.Y(n_696)
);

XOR2xp5_ASAP7_75t_L g697 ( 
.A(n_495),
.B(n_206),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_554),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_503),
.B(n_309),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_554),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_493),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_493),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_554),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_493),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_515),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_523),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_705),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_696),
.B(n_195),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_610),
.A2(n_306),
.B1(n_376),
.B2(n_373),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_651),
.A2(n_541),
.B1(n_301),
.B2(n_308),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_585),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_557),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_610),
.B(n_261),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_557),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_651),
.B(n_503),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_L g716 ( 
.A1(n_639),
.A2(n_445),
.B(n_421),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_705),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_614),
.B(n_503),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_696),
.B(n_197),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_560),
.A2(n_562),
.B1(n_571),
.B2(n_567),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_706),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_706),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_594),
.B(n_503),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_572),
.Y(n_724)
);

OR2x2_ASAP7_75t_SL g725 ( 
.A(n_564),
.B(n_495),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_560),
.A2(n_541),
.B1(n_290),
.B2(n_314),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_608),
.B(n_494),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_596),
.A2(n_541),
.B1(n_324),
.B2(n_319),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_594),
.B(n_525),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_577),
.B(n_197),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_686),
.B(n_525),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_686),
.B(n_568),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_572),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_638),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_701),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_L g736 ( 
.A1(n_674),
.A2(n_609),
.B1(n_595),
.B2(n_575),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_673),
.B(n_677),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_572),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_701),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_699),
.B(n_559),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_559),
.B(n_525),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_609),
.B(n_198),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_572),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_673),
.B(n_631),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_559),
.B(n_525),
.Y(n_745)
);

AND2x6_ASAP7_75t_L g746 ( 
.A(n_613),
.B(n_261),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_559),
.B(n_501),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_574),
.A2(n_261),
.B1(n_350),
.B2(n_359),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_629),
.B(n_198),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_702),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_631),
.B(n_517),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_613),
.B(n_501),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_580),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_660),
.B(n_199),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_580),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_702),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_574),
.A2(n_687),
.B1(n_613),
.B2(n_620),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_620),
.B(n_501),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_580),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_561),
.B(n_622),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_617),
.B(n_199),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_564),
.B(n_517),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_704),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_620),
.B(n_508),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_704),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_661),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_638),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_558),
.A2(n_326),
.B1(n_318),
.B2(n_332),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_561),
.B(n_212),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_573),
.B(n_508),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_589),
.B(n_508),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_589),
.B(n_509),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_603),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_574),
.A2(n_350),
.B1(n_359),
.B2(n_295),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_595),
.B(n_523),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_597),
.B(n_509),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_603),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_597),
.B(n_509),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_561),
.B(n_212),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_678),
.B(n_222),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_598),
.B(n_497),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_598),
.B(n_512),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_561),
.B(n_222),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_578),
.B(n_582),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_601),
.B(n_512),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_616),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_L g787 ( 
.A(n_574),
.B(n_333),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_575),
.A2(n_601),
.B(n_679),
.C(n_625),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_580),
.B(n_512),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_616),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_626),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_590),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_581),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_581),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_581),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_626),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_634),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_634),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_679),
.A2(n_336),
.B1(n_340),
.B2(n_338),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_581),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_592),
.B(n_350),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_691),
.A2(n_540),
.B(n_536),
.C(n_535),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_635),
.B(n_528),
.C(n_527),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_592),
.B(n_350),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_592),
.B(n_512),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_659),
.B(n_223),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_592),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_680),
.B(n_512),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_633),
.B(n_574),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_574),
.B(n_512),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_657),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_641),
.Y(n_812)
);

NAND2x1_ASAP7_75t_L g813 ( 
.A(n_584),
.B(n_485),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_574),
.A2(n_359),
.B1(n_343),
.B2(n_312),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_618),
.B(n_512),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_618),
.B(n_334),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_618),
.B(n_513),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_SL g818 ( 
.A1(n_648),
.A2(n_305),
.B1(n_374),
.B2(n_272),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_602),
.B(n_223),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_692),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_607),
.B(n_224),
.Y(n_821)
);

INVx8_ASAP7_75t_L g822 ( 
.A(n_590),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_640),
.B(n_513),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_640),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_L g825 ( 
.A(n_641),
.B(n_359),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_697),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_619),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_643),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_644),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_644),
.B(n_513),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_619),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_625),
.B(n_224),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_649),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_649),
.B(n_513),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_654),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_654),
.Y(n_836)
);

NOR2x1p5_ASAP7_75t_L g837 ( 
.A(n_682),
.B(n_206),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_669),
.B(n_513),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_669),
.B(n_513),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_681),
.B(n_225),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_681),
.B(n_684),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_682),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_556),
.A2(n_225),
.B1(n_286),
.B2(n_361),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_684),
.A2(n_293),
.B1(n_335),
.B2(n_368),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_671),
.B(n_676),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_685),
.B(n_492),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_685),
.B(n_492),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_688),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_653),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_688),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_698),
.B(n_499),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_698),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_556),
.B(n_528),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_700),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_700),
.B(n_286),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_703),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_L g857 ( 
.A(n_658),
.B(n_529),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_703),
.B(n_555),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_611),
.B(n_529),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_591),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_555),
.B(n_499),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_L g862 ( 
.A(n_667),
.B(n_351),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_565),
.B(n_500),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_565),
.A2(n_266),
.B(n_270),
.C(n_273),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_583),
.B(n_500),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_583),
.B(n_502),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_588),
.A2(n_361),
.B1(n_358),
.B2(n_355),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_588),
.B(n_311),
.Y(n_868)
);

BUFx6f_ASAP7_75t_SL g869 ( 
.A(n_653),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_584),
.B(n_502),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_670),
.B(n_351),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_563),
.A2(n_316),
.B(n_317),
.C(n_322),
.Y(n_872)
);

NOR3xp33_ASAP7_75t_L g873 ( 
.A(n_672),
.B(n_536),
.C(n_535),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_591),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_584),
.B(n_355),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_853),
.B(n_540),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_732),
.B(n_611),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_734),
.B(n_767),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_850),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_850),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_718),
.B(n_611),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_812),
.B(n_418),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_715),
.B(n_707),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_775),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_744),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_749),
.A2(n_630),
.B1(n_612),
.B2(n_693),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_717),
.B(n_611),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_721),
.B(n_621),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_749),
.A2(n_695),
.B1(n_612),
.B2(n_693),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_737),
.B(n_358),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_811),
.B(n_231),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_775),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_724),
.Y(n_893)
);

OR2x2_ASAP7_75t_SL g894 ( 
.A(n_762),
.B(n_325),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_722),
.B(n_621),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_727),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_733),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_738),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_SL g899 ( 
.A(n_818),
.B(n_208),
.C(n_207),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_784),
.A2(n_636),
.B1(n_689),
.B2(n_683),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_736),
.B(n_585),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_803),
.B(n_421),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_784),
.B(n_585),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_740),
.B(n_621),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_723),
.B(n_621),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_720),
.B(n_423),
.Y(n_906)
);

OR2x2_ASAP7_75t_SL g907 ( 
.A(n_725),
.B(n_337),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_820),
.B(n_585),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_845),
.A2(n_584),
.B(n_615),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_743),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_742),
.B(n_627),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_742),
.B(n_627),
.Y(n_912)
);

OR2x6_ASAP7_75t_L g913 ( 
.A(n_822),
.B(n_423),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_821),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_757),
.B(n_585),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_841),
.A2(n_780),
.B1(n_719),
.B2(n_708),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_753),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_729),
.B(n_859),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_755),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_751),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_821),
.Y(n_921)
);

NOR3xp33_ASAP7_75t_SL g922 ( 
.A(n_760),
.B(n_209),
.C(n_208),
.Y(n_922)
);

NOR3xp33_ASAP7_75t_SL g923 ( 
.A(n_840),
.B(n_210),
.C(n_209),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_759),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_793),
.Y(n_925)
);

NAND2x1p5_ASAP7_75t_L g926 ( 
.A(n_794),
.B(n_627),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_841),
.B(n_627),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_795),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_819),
.B(n_429),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_761),
.B(n_586),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_819),
.B(n_429),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_712),
.B(n_642),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_855),
.B(n_642),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_751),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_827),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_773),
.Y(n_936)
);

AND2x6_ASAP7_75t_SL g937 ( 
.A(n_751),
.B(n_432),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_780),
.A2(n_642),
.B1(n_655),
.B2(n_695),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_800),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_807),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_761),
.B(n_432),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_773),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_873),
.A2(n_642),
.B1(n_655),
.B2(n_689),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_855),
.B(n_757),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_875),
.B(n_655),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_806),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_792),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_806),
.B(n_433),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_831),
.B(n_842),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_777),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_788),
.A2(n_566),
.B(n_563),
.Y(n_951)
);

INVx5_ASAP7_75t_L g952 ( 
.A(n_746),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_741),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_766),
.Y(n_954)
);

CKINVDCx8_ASAP7_75t_R g955 ( 
.A(n_822),
.Y(n_955)
);

AND2x6_ASAP7_75t_L g956 ( 
.A(n_712),
.B(n_566),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_714),
.B(n_655),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_769),
.B(n_234),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_745),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_714),
.B(n_569),
.Y(n_960)
);

NAND3xp33_ASAP7_75t_SL g961 ( 
.A(n_843),
.B(n_211),
.C(n_210),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_777),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_786),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_709),
.A2(n_630),
.B1(n_623),
.B2(n_683),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_786),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_858),
.B(n_569),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_710),
.B(n_586),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_754),
.B(n_435),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_790),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_790),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_791),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_791),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_796),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_796),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_858),
.B(n_570),
.Y(n_975)
);

AO22x2_ASAP7_75t_L g976 ( 
.A1(n_779),
.A2(n_435),
.B1(n_436),
.B2(n_437),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_797),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_783),
.B(n_237),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_869),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_SL g980 ( 
.A1(n_826),
.A2(n_345),
.B1(n_216),
.B2(n_218),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_875),
.B(n_570),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_730),
.B(n_238),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_798),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_828),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_828),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_822),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_869),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_837),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_836),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_836),
.B(n_576),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_770),
.B(n_576),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_799),
.B(n_586),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_845),
.A2(n_587),
.B(n_579),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_848),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_848),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_849),
.B(n_436),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_824),
.A2(n_624),
.B1(n_628),
.B2(n_675),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_854),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_854),
.B(n_579),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_856),
.B(n_587),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_867),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_856),
.B(n_829),
.Y(n_1002)
);

INVx5_ASAP7_75t_L g1003 ( 
.A(n_746),
.Y(n_1003)
);

BUFx4f_ASAP7_75t_L g1004 ( 
.A(n_746),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_833),
.B(n_624),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_735),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_728),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_835),
.B(n_628),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_852),
.B(n_632),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_861),
.Y(n_1010)
);

BUFx4f_ASAP7_75t_L g1011 ( 
.A(n_746),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_SL g1012 ( 
.A1(n_825),
.A2(n_305),
.B1(n_374),
.B2(n_218),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_863),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_865),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_816),
.A2(n_662),
.B1(n_645),
.B2(n_675),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_746),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_726),
.Y(n_1017)
);

CKINVDCx16_ASAP7_75t_R g1018 ( 
.A(n_768),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_752),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_731),
.B(n_713),
.Y(n_1020)
);

BUFx12f_ASAP7_75t_L g1021 ( 
.A(n_716),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_L g1022 ( 
.A(n_832),
.B(n_285),
.C(n_296),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_747),
.B(n_437),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_866),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_713),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_758),
.B(n_632),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_860),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_860),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_871),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_735),
.B(n_739),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_SL g1031 ( 
.A(n_802),
.B(n_374),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_748),
.A2(n_690),
.B1(n_226),
.B2(n_216),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_857),
.B(n_586),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_764),
.A2(n_652),
.B1(n_666),
.B2(n_665),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_711),
.B(n_636),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_808),
.B(n_846),
.Y(n_1036)
);

BUFx8_ASAP7_75t_L g1037 ( 
.A(n_739),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_847),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_874),
.Y(n_1039)
);

AO22x1_ASAP7_75t_L g1040 ( 
.A1(n_809),
.A2(n_211),
.B1(n_226),
.B2(n_345),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_750),
.B(n_637),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_R g1042 ( 
.A(n_862),
.B(n_787),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_851),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_756),
.B(n_637),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_756),
.B(n_439),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_SL g1046 ( 
.A1(n_748),
.A2(n_349),
.B1(n_346),
.B2(n_348),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_763),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_870),
.A2(n_662),
.B1(n_666),
.B2(n_665),
.Y(n_1048)
);

AND2x2_ASAP7_75t_SL g1049 ( 
.A(n_774),
.B(n_439),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_765),
.B(n_771),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_844),
.B(n_442),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_765),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_868),
.B(n_442),
.C(n_307),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_813),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_772),
.B(n_645),
.Y(n_1055)
);

NOR3xp33_ASAP7_75t_L g1056 ( 
.A(n_868),
.B(n_291),
.C(n_243),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_844),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_776),
.B(n_650),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_778),
.B(n_650),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_815),
.B(n_487),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_789),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_914),
.B(n_817),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_SL g1063 ( 
.A(n_916),
.B(n_348),
.C(n_346),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_993),
.A2(n_805),
.B(n_781),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_946),
.A2(n_864),
.B(n_872),
.C(n_801),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_878),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_944),
.A2(n_982),
.B(n_978),
.C(n_958),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_918),
.A2(n_774),
.B(n_646),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_1037),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_921),
.B(n_814),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_1057),
.A2(n_782),
.B(n_785),
.C(n_810),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_884),
.A2(n_814),
.B1(n_804),
.B2(n_801),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_896),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1010),
.B(n_823),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_929),
.B(n_487),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_884),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_890),
.A2(n_804),
.B(n_838),
.C(n_834),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_974),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_884),
.B(n_830),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_SL g1080 ( 
.A(n_899),
.B(n_349),
.C(n_352),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_915),
.A2(n_615),
.B(n_646),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_904),
.A2(n_615),
.B(n_646),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1013),
.B(n_839),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_904),
.A2(n_615),
.B(n_646),
.Y(n_1084)
);

CKINVDCx14_ASAP7_75t_R g1085 ( 
.A(n_954),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_931),
.B(n_586),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_961),
.A2(n_664),
.B(n_656),
.C(n_652),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1001),
.A2(n_664),
.B1(n_656),
.B2(n_488),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_983),
.B(n_605),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_876),
.A2(n_1023),
.B1(n_1017),
.B2(n_941),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_945),
.A2(n_981),
.B(n_881),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_942),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1029),
.A2(n_488),
.B1(n_663),
.B2(n_647),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_881),
.A2(n_605),
.B(n_663),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_905),
.A2(n_605),
.B(n_663),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_901),
.A2(n_479),
.B(n_604),
.C(n_600),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_930),
.A2(n_903),
.B(n_927),
.Y(n_1097)
);

AND3x1_ASAP7_75t_SL g1098 ( 
.A(n_937),
.B(n_372),
.C(n_360),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_974),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_983),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_963),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_905),
.A2(n_605),
.B(n_663),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_983),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_876),
.B(n_479),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1006),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_948),
.B(n_247),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1018),
.B(n_605),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1006),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_995),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_927),
.A2(n_975),
.B(n_966),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_L g1111 ( 
.A(n_953),
.B(n_647),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_891),
.B(n_265),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_996),
.B(n_647),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_885),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_986),
.B(n_514),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1023),
.A2(n_694),
.B1(n_514),
.B2(n_526),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1014),
.B(n_593),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_960),
.A2(n_647),
.B(n_663),
.Y(n_1118)
);

INVxp67_ASAP7_75t_SL g1119 ( 
.A(n_995),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_972),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_996),
.B(n_647),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_SL g1122 ( 
.A(n_955),
.B(n_353),
.Y(n_1122)
);

BUFx8_ASAP7_75t_SL g1123 ( 
.A(n_979),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_936),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1038),
.B(n_276),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_960),
.A2(n_668),
.B(n_599),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1037),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_909),
.A2(n_668),
.B(n_599),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1007),
.A2(n_514),
.B1(n_526),
.B2(n_606),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1024),
.B(n_593),
.Y(n_1130)
);

AND2x6_ASAP7_75t_L g1131 ( 
.A(n_1036),
.B(n_600),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_883),
.A2(n_287),
.B(n_289),
.C(n_304),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1043),
.B(n_947),
.Y(n_1133)
);

BUFx4f_ASAP7_75t_L g1134 ( 
.A(n_913),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_995),
.B(n_668),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_947),
.B(n_313),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_892),
.A2(n_694),
.B1(n_526),
.B2(n_320),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_894),
.B(n_341),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_932),
.A2(n_668),
.B(n_606),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_935),
.B(n_331),
.Y(n_1140)
);

BUFx12f_ASAP7_75t_L g1141 ( 
.A(n_987),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_968),
.A2(n_604),
.B1(n_694),
.B2(n_372),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_883),
.B(n_485),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1053),
.A2(n_360),
.B(n_357),
.C(n_356),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_988),
.B(n_122),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_SL g1146 ( 
.A(n_1049),
.B(n_357),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_953),
.B(n_694),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_932),
.A2(n_668),
.B(n_694),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1022),
.A2(n_694),
.B1(n_356),
.B2(n_353),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_950),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_949),
.B(n_882),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_920),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_R g1153 ( 
.A(n_987),
.B(n_185),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_998),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_957),
.A2(n_668),
.B(n_694),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1025),
.A2(n_0),
.B(n_6),
.C(n_7),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_957),
.A2(n_181),
.B(n_172),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_877),
.A2(n_164),
.B(n_155),
.Y(n_1158)
);

INVxp67_ASAP7_75t_SL g1159 ( 
.A(n_998),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_973),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_879),
.B(n_142),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_L g1162 ( 
.A(n_980),
.B(n_934),
.C(n_1040),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_906),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_966),
.A2(n_134),
.B(n_130),
.Y(n_1164)
);

OAI22x1_ASAP7_75t_L g1165 ( 
.A1(n_906),
.A2(n_902),
.B1(n_907),
.B2(n_1025),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_953),
.B(n_113),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_962),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1051),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_959),
.B(n_1019),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_880),
.B(n_111),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_965),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_975),
.A2(n_102),
.B(n_89),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_998),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_959),
.B(n_87),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1056),
.A2(n_14),
.B(n_20),
.C(n_22),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_959),
.B(n_73),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_933),
.A2(n_70),
.B(n_68),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1019),
.B(n_62),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_902),
.A2(n_20),
.B(n_24),
.C(n_25),
.Y(n_1179)
);

INVx5_ASAP7_75t_L g1180 ( 
.A(n_956),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1002),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1021),
.B(n_29),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_913),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_913),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1060),
.B(n_30),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1050),
.A2(n_31),
.B(n_36),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_919),
.Y(n_1187)
);

AO21x1_ASAP7_75t_L g1188 ( 
.A1(n_1031),
.A2(n_37),
.B(n_38),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_1045),
.Y(n_1189)
);

AND2x2_ASAP7_75t_SL g1190 ( 
.A(n_1031),
.B(n_37),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1019),
.B(n_38),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_922),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1045),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_R g1194 ( 
.A(n_919),
.B(n_42),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_925),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_984),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_969),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1050),
.A2(n_42),
.B(n_43),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1061),
.B(n_911),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_912),
.B(n_43),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1002),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_L g1202 ( 
.A(n_1012),
.B(n_1046),
.C(n_1032),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_923),
.B(n_47),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_925),
.B(n_48),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_994),
.Y(n_1205)
);

AOI22x1_ASAP7_75t_L g1206 ( 
.A1(n_976),
.A2(n_977),
.B1(n_985),
.B2(n_971),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_926),
.Y(n_1207)
);

BUFx8_ASAP7_75t_SL g1208 ( 
.A(n_1004),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_956),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_970),
.B(n_989),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_893),
.B(n_50),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_897),
.B(n_50),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1047),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_976),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_898),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_992),
.A2(n_51),
.B(n_55),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1032),
.A2(n_56),
.B(n_59),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_910),
.B(n_59),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1035),
.A2(n_991),
.B(n_1020),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_908),
.A2(n_967),
.B(n_939),
.C(n_917),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1055),
.A2(n_1058),
.B(n_1026),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1067),
.A2(n_1112),
.B(n_1200),
.C(n_1202),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1091),
.A2(n_1008),
.A3(n_1005),
.B(n_1009),
.Y(n_1223)
);

NOR2xp67_ASAP7_75t_L g1224 ( 
.A(n_1114),
.B(n_900),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1075),
.B(n_1055),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1064),
.A2(n_951),
.B(n_999),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1128),
.A2(n_951),
.B(n_999),
.Y(n_1227)
);

INVx8_ASAP7_75t_L g1228 ( 
.A(n_1141),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1221),
.A2(n_1058),
.B(n_1059),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1090),
.B(n_1011),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1081),
.A2(n_990),
.B(n_1000),
.Y(n_1231)
);

INVx5_ASAP7_75t_L g1232 ( 
.A(n_1209),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1066),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1092),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1151),
.B(n_1011),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1074),
.B(n_940),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_SL g1237 ( 
.A1(n_1071),
.A2(n_1060),
.B(n_1033),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1094),
.A2(n_1000),
.B(n_990),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1074),
.B(n_924),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1083),
.B(n_928),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1133),
.B(n_1125),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1189),
.B(n_1060),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_SL g1243 ( 
.A(n_1190),
.B(n_1004),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1213),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1101),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1219),
.A2(n_886),
.B(n_889),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1120),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1073),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1077),
.A2(n_1048),
.B(n_1044),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1110),
.A2(n_1009),
.B(n_1008),
.Y(n_1250)
);

AO21x1_ASAP7_75t_L g1251 ( 
.A1(n_1216),
.A2(n_1005),
.B(n_888),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1111),
.A2(n_1016),
.B(n_1003),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1199),
.B(n_1030),
.Y(n_1253)
);

AO21x2_ASAP7_75t_L g1254 ( 
.A1(n_1097),
.A2(n_1015),
.B(n_1042),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1095),
.A2(n_887),
.B(n_888),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1189),
.B(n_1039),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1193),
.B(n_1104),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1068),
.A2(n_1044),
.B(n_1041),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1199),
.B(n_1030),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1146),
.B(n_1134),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1082),
.A2(n_1016),
.B(n_1003),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1104),
.B(n_1076),
.Y(n_1262)
);

AOI221xp5_ASAP7_75t_L g1263 ( 
.A1(n_1138),
.A2(n_1052),
.B1(n_895),
.B2(n_887),
.C(n_938),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1102),
.A2(n_895),
.B(n_926),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1084),
.A2(n_1003),
.B(n_952),
.Y(n_1265)
);

INVx5_ASAP7_75t_L g1266 ( 
.A(n_1209),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1083),
.A2(n_1003),
.B(n_952),
.Y(n_1267)
);

INVxp67_ASAP7_75t_SL g1268 ( 
.A(n_1187),
.Y(n_1268)
);

AO32x2_ASAP7_75t_L g1269 ( 
.A1(n_1181),
.A2(n_1201),
.A3(n_1168),
.B1(n_1214),
.B2(n_1109),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1118),
.A2(n_1034),
.B(n_997),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1152),
.B(n_1028),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1139),
.A2(n_1027),
.B(n_964),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1126),
.A2(n_943),
.B(n_956),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1169),
.B(n_956),
.Y(n_1274)
);

AND3x1_ASAP7_75t_L g1275 ( 
.A(n_1080),
.B(n_952),
.C(n_1016),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1152),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1160),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1169),
.B(n_1054),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1187),
.Y(n_1279)
);

AOI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1086),
.A2(n_1079),
.B(n_1143),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1144),
.A2(n_1054),
.B(n_1063),
.C(n_1146),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1076),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1123),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1206),
.A2(n_1054),
.B(n_1096),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1062),
.B(n_1215),
.Y(n_1285)
);

BUFx8_ASAP7_75t_L g1286 ( 
.A(n_1183),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1180),
.A2(n_1220),
.B(n_1130),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1065),
.A2(n_1217),
.B(n_1175),
.C(n_1132),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1087),
.A2(n_1155),
.B(n_1148),
.Y(n_1289)
);

NOR4xp25_ASAP7_75t_L g1290 ( 
.A(n_1168),
.B(n_1201),
.C(n_1181),
.D(n_1179),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_SL g1291 ( 
.A(n_1180),
.B(n_1069),
.Y(n_1291)
);

AOI21xp33_ASAP7_75t_L g1292 ( 
.A1(n_1165),
.A2(n_1188),
.B(n_1070),
.Y(n_1292)
);

OAI21xp33_ASAP7_75t_L g1293 ( 
.A1(n_1140),
.A2(n_1163),
.B(n_1212),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1085),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1187),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1196),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1180),
.A2(n_1130),
.B(n_1117),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1205),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1166),
.A2(n_1174),
.B(n_1207),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1162),
.A2(n_1192),
.B1(n_1107),
.B2(n_1136),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1134),
.B(n_1122),
.Y(n_1301)
);

INVx5_ASAP7_75t_L g1302 ( 
.A(n_1209),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1072),
.A2(n_1113),
.B1(n_1121),
.B2(n_1117),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1124),
.B(n_1171),
.Y(n_1304)
);

AOI211x1_ASAP7_75t_L g1305 ( 
.A1(n_1203),
.A2(n_1198),
.B(n_1186),
.C(n_1204),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1210),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1150),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1167),
.B(n_1197),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1119),
.A2(n_1159),
.B(n_1177),
.Y(n_1309)
);

OAI21xp33_ASAP7_75t_L g1310 ( 
.A1(n_1211),
.A2(n_1182),
.B(n_1122),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1210),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1078),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1164),
.A2(n_1172),
.B(n_1158),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1157),
.A2(n_1178),
.B(n_1176),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1129),
.A2(n_1131),
.B(n_1191),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1076),
.B(n_1195),
.Y(n_1316)
);

AOI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1161),
.A2(n_1170),
.B(n_1147),
.Y(n_1317)
);

AO21x1_ASAP7_75t_L g1318 ( 
.A1(n_1147),
.A2(n_1089),
.B(n_1093),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1099),
.B(n_1103),
.Y(n_1319)
);

NOR2x1_ASAP7_75t_SL g1320 ( 
.A(n_1195),
.B(n_1173),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1115),
.A2(n_1105),
.B(n_1108),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1195),
.B(n_1194),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1100),
.B(n_1154),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1218),
.B(n_1145),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1218),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1184),
.B(n_1145),
.Y(n_1326)
);

INVx5_ASAP7_75t_L g1327 ( 
.A(n_1208),
.Y(n_1327)
);

AO21x1_ASAP7_75t_L g1328 ( 
.A1(n_1109),
.A2(n_1154),
.B(n_1135),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1131),
.B(n_1088),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1173),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1156),
.A2(n_1116),
.B(n_1142),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1131),
.A2(n_1185),
.A3(n_1137),
.B(n_1149),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1185),
.B(n_1127),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1131),
.B(n_1173),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1185),
.A2(n_1153),
.B(n_1098),
.Y(n_1335)
);

INVxp67_ASAP7_75t_SL g1336 ( 
.A(n_1111),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1075),
.B(n_929),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1064),
.A2(n_993),
.B(n_1128),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1064),
.A2(n_993),
.B(n_1128),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1066),
.Y(n_1340)
);

AOI221x1_ASAP7_75t_L g1341 ( 
.A1(n_1067),
.A2(n_1202),
.B1(n_1217),
.B2(n_1216),
.C(n_1165),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1064),
.A2(n_993),
.B(n_1128),
.Y(n_1342)
);

AO32x2_ASAP7_75t_L g1343 ( 
.A1(n_1181),
.A2(n_1201),
.A3(n_1168),
.B1(n_709),
.B2(n_651),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1106),
.B(n_1151),
.Y(n_1344)
);

AOI21xp33_ASAP7_75t_L g1345 ( 
.A1(n_1067),
.A2(n_1112),
.B(n_916),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1064),
.A2(n_993),
.B(n_1128),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1213),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1067),
.A2(n_1112),
.B(n_916),
.C(n_749),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1112),
.B(n_393),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1067),
.A2(n_1091),
.B(n_1221),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1066),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1066),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1091),
.A2(n_1221),
.B(n_1219),
.Y(n_1353)
);

AOI221xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1217),
.A2(n_1067),
.B1(n_1168),
.B2(n_916),
.C(n_1181),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1213),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_SL g1356 ( 
.A1(n_1217),
.A2(n_1067),
.B1(n_1168),
.B2(n_916),
.C(n_1181),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1067),
.A2(n_1112),
.B(n_916),
.C(n_749),
.Y(n_1357)
);

AOI31xp67_ASAP7_75t_L g1358 ( 
.A1(n_1086),
.A2(n_901),
.A3(n_992),
.B(n_930),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1064),
.A2(n_993),
.B(n_1128),
.Y(n_1359)
);

NOR4xp25_ASAP7_75t_L g1360 ( 
.A(n_1067),
.B(n_1217),
.C(n_1175),
.D(n_1168),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1067),
.B(n_1010),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1091),
.A2(n_1221),
.B(n_1219),
.Y(n_1362)
);

NOR2xp67_ASAP7_75t_L g1363 ( 
.A(n_1114),
.B(n_827),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1064),
.A2(n_993),
.B(n_1128),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1067),
.A2(n_1091),
.B(n_1221),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_SL g1366 ( 
.A1(n_1188),
.A2(n_1206),
.B(n_1174),
.Y(n_1366)
);

OAI22x1_ASAP7_75t_L g1367 ( 
.A1(n_1214),
.A2(n_697),
.B1(n_1192),
.B2(n_1112),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1067),
.A2(n_1112),
.B(n_916),
.C(n_749),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1067),
.A2(n_1091),
.B(n_1221),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1123),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1067),
.B(n_1010),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1091),
.A2(n_1221),
.B(n_1219),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1213),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1091),
.A2(n_1221),
.B(n_1219),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1067),
.B(n_1010),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1064),
.A2(n_993),
.B(n_1128),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1091),
.A2(n_1221),
.B(n_1219),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1064),
.A2(n_993),
.B(n_1128),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1293),
.A2(n_1360),
.B1(n_1345),
.B2(n_1222),
.C(n_1290),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1235),
.B(n_1242),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1340),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1353),
.A2(n_1372),
.B(n_1362),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1348),
.A2(n_1368),
.B(n_1357),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1234),
.Y(n_1384)
);

BUFx12f_ASAP7_75t_L g1385 ( 
.A(n_1370),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1245),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1233),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_SL g1388 ( 
.A1(n_1345),
.A2(n_1288),
.B(n_1281),
.C(n_1375),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1350),
.A2(n_1369),
.B(n_1365),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1276),
.B(n_1325),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1294),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1351),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1310),
.A2(n_1367),
.B1(n_1349),
.B2(n_1241),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1374),
.A2(n_1377),
.B(n_1289),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1352),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1337),
.B(n_1344),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1276),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1306),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_SL g1399 ( 
.A1(n_1366),
.A2(n_1315),
.B(n_1318),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1346),
.A2(n_1364),
.B(n_1359),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1282),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1325),
.A2(n_1336),
.B1(n_1300),
.B2(n_1260),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1292),
.A2(n_1375),
.B1(n_1371),
.B2(n_1361),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_SL g1404 ( 
.A(n_1283),
.B(n_1327),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1376),
.A2(n_1378),
.B(n_1226),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1244),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1354),
.A2(n_1356),
.B(n_1361),
.C(n_1371),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1232),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1264),
.A2(n_1238),
.B(n_1231),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1255),
.A2(n_1272),
.B(n_1227),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1285),
.B(n_1243),
.Y(n_1411)
);

OR2x6_ASAP7_75t_L g1412 ( 
.A(n_1305),
.B(n_1237),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1311),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1315),
.B(n_1230),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1247),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1278),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1277),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1243),
.B(n_1322),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1258),
.A2(n_1284),
.B(n_1229),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1248),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1246),
.A2(n_1249),
.B(n_1287),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1292),
.A2(n_1360),
.B(n_1301),
.C(n_1290),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1236),
.A2(n_1240),
.B1(n_1239),
.B2(n_1224),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1278),
.Y(n_1424)
);

OAI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1354),
.A2(n_1356),
.B1(n_1335),
.B2(n_1326),
.C(n_1333),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1253),
.B(n_1259),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1304),
.B(n_1308),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1246),
.A2(n_1225),
.B(n_1249),
.C(n_1236),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1271),
.B(n_1256),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1242),
.A2(n_1331),
.B1(n_1239),
.B2(n_1240),
.Y(n_1430)
);

INVx5_ASAP7_75t_L g1431 ( 
.A(n_1282),
.Y(n_1431)
);

AOI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1303),
.A2(n_1263),
.B1(n_1257),
.B2(n_1355),
.C(n_1347),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1258),
.A2(n_1299),
.B(n_1273),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1331),
.A2(n_1373),
.B1(n_1298),
.B2(n_1296),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1257),
.B(n_1341),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1297),
.A2(n_1261),
.B(n_1265),
.Y(n_1436)
);

AO32x2_ASAP7_75t_L g1437 ( 
.A1(n_1343),
.A2(n_1269),
.A3(n_1358),
.B1(n_1295),
.B2(n_1330),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1307),
.A2(n_1251),
.B1(n_1312),
.B2(n_1314),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1286),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_R g1440 ( 
.A(n_1327),
.B(n_1228),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1314),
.A2(n_1286),
.B1(n_1327),
.B2(n_1313),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1319),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1232),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1270),
.A2(n_1280),
.B(n_1309),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1250),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1317),
.A2(n_1267),
.B(n_1274),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1321),
.A2(n_1313),
.B(n_1252),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1319),
.Y(n_1448)
);

AO21x2_ASAP7_75t_L g1449 ( 
.A1(n_1254),
.A2(n_1334),
.B(n_1328),
.Y(n_1449)
);

NAND2x1p5_ASAP7_75t_L g1450 ( 
.A(n_1291),
.B(n_1266),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1363),
.A2(n_1262),
.B1(n_1268),
.B2(n_1279),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1316),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1254),
.A2(n_1320),
.B(n_1232),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1223),
.A2(n_1343),
.B(n_1269),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1223),
.A2(n_1343),
.B(n_1269),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1223),
.A2(n_1332),
.B(n_1275),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1282),
.B(n_1295),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1232),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1323),
.A2(n_1332),
.B(n_1266),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1266),
.A2(n_1302),
.B(n_1330),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1332),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1266),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1302),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1302),
.A2(n_1348),
.B(n_1368),
.C(n_1357),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1302),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1228),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1348),
.A2(n_1067),
.B(n_1357),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1234),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1282),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1276),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1235),
.B(n_1242),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1276),
.B(n_1325),
.Y(n_1472)
);

AOI21xp33_ASAP7_75t_L g1473 ( 
.A1(n_1222),
.A2(n_1293),
.B(n_1112),
.Y(n_1473)
);

AND2x6_ASAP7_75t_L g1474 ( 
.A(n_1329),
.B(n_1209),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1340),
.Y(n_1475)
);

OR2x6_ASAP7_75t_L g1476 ( 
.A(n_1305),
.B(n_1237),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1338),
.A2(n_1342),
.B(n_1339),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1233),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1222),
.A2(n_1057),
.B1(n_1067),
.B2(n_1348),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1234),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_SL g1481 ( 
.A1(n_1348),
.A2(n_1357),
.B(n_1368),
.C(n_1222),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1337),
.A2(n_1146),
.B1(n_1057),
.B2(n_1168),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1234),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1337),
.B(n_1349),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1337),
.B(n_1349),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1233),
.Y(n_1486)
);

BUFx4f_ASAP7_75t_L g1487 ( 
.A(n_1228),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1350),
.A2(n_1369),
.B(n_1365),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1350),
.A2(n_1369),
.B(n_1365),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1337),
.B(n_1349),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1338),
.A2(n_1342),
.B(n_1339),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_SL g1492 ( 
.A1(n_1366),
.A2(n_1188),
.B(n_1315),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1233),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1234),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1234),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1234),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1337),
.B(n_1349),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1338),
.A2(n_1342),
.B(n_1339),
.Y(n_1498)
);

AO32x2_ASAP7_75t_L g1499 ( 
.A1(n_1303),
.A2(n_1181),
.A3(n_1201),
.B1(n_1168),
.B2(n_1343),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1233),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1344),
.B(n_1324),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1338),
.A2(n_1342),
.B(n_1339),
.Y(n_1502)
);

AO22x2_ASAP7_75t_L g1503 ( 
.A1(n_1341),
.A2(n_1305),
.B1(n_1202),
.B2(n_1366),
.Y(n_1503)
);

O2A1O1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1222),
.A2(n_1357),
.B(n_1368),
.C(n_1348),
.Y(n_1504)
);

BUFx12f_ASAP7_75t_L g1505 ( 
.A(n_1370),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1338),
.A2(n_1342),
.B(n_1339),
.Y(n_1506)
);

NAND2x1p5_ASAP7_75t_L g1507 ( 
.A(n_1291),
.B(n_1180),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1338),
.A2(n_1342),
.B(n_1339),
.Y(n_1508)
);

INVx3_ASAP7_75t_SL g1509 ( 
.A(n_1294),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1340),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1338),
.A2(n_1342),
.B(n_1339),
.Y(n_1511)
);

NAND2x1p5_ASAP7_75t_L g1512 ( 
.A(n_1291),
.B(n_1180),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1348),
.A2(n_1067),
.B(n_1357),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1233),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1233),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1420),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1415),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1415),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1428),
.A2(n_1479),
.B(n_1504),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1426),
.B(n_1429),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1462),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1501),
.B(n_1411),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1393),
.A2(n_1379),
.B1(n_1482),
.B2(n_1403),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1393),
.A2(n_1482),
.B1(n_1403),
.B2(n_1490),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1411),
.B(n_1396),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1428),
.A2(n_1450),
.B(n_1464),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1427),
.B(n_1484),
.Y(n_1527)
);

AOI211xp5_ASAP7_75t_L g1528 ( 
.A1(n_1473),
.A2(n_1513),
.B(n_1467),
.C(n_1481),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1485),
.A2(n_1497),
.B1(n_1418),
.B2(n_1425),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1390),
.B(n_1472),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1392),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1406),
.Y(n_1532)
);

CKINVDCx11_ASAP7_75t_R g1533 ( 
.A(n_1385),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1407),
.A2(n_1383),
.B1(n_1414),
.B2(n_1422),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1417),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1397),
.B(n_1470),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1470),
.B(n_1442),
.Y(n_1537)
);

O2A1O1Ixp5_ASAP7_75t_L g1538 ( 
.A1(n_1423),
.A2(n_1464),
.B(n_1446),
.C(n_1407),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1381),
.Y(n_1539)
);

O2A1O1Ixp5_ASAP7_75t_L g1540 ( 
.A1(n_1453),
.A2(n_1402),
.B(n_1451),
.C(n_1380),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1481),
.A2(n_1388),
.B(n_1492),
.C(n_1414),
.Y(n_1541)
);

OA21x2_ASAP7_75t_L g1542 ( 
.A1(n_1419),
.A2(n_1410),
.B(n_1447),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1450),
.A2(n_1507),
.B(n_1512),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1414),
.A2(n_1503),
.B1(n_1430),
.B2(n_1413),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1433),
.A2(n_1409),
.B(n_1400),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1388),
.A2(n_1399),
.B(n_1510),
.C(n_1475),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1503),
.A2(n_1430),
.B1(n_1398),
.B2(n_1413),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1448),
.B(n_1398),
.Y(n_1548)
);

AOI31xp33_ASAP7_75t_L g1549 ( 
.A1(n_1432),
.A2(n_1441),
.A3(n_1507),
.B(n_1512),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1503),
.A2(n_1434),
.B1(n_1488),
.B2(n_1489),
.Y(n_1550)
);

OA21x2_ASAP7_75t_L g1551 ( 
.A1(n_1400),
.A2(n_1498),
.B(n_1511),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1468),
.B(n_1496),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1412),
.A2(n_1476),
.B(n_1424),
.C(n_1416),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1424),
.B(n_1496),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_SL g1555 ( 
.A1(n_1462),
.A2(n_1460),
.B(n_1443),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1384),
.B(n_1386),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1466),
.B(n_1392),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1385),
.Y(n_1558)
);

O2A1O1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1412),
.A2(n_1476),
.B(n_1421),
.C(n_1466),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1478),
.B(n_1514),
.Y(n_1560)
);

NOR2xp67_ASAP7_75t_L g1561 ( 
.A(n_1395),
.B(n_1493),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1480),
.B(n_1483),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1505),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1434),
.A2(n_1488),
.B1(n_1489),
.B2(n_1389),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1389),
.A2(n_1488),
.B1(n_1489),
.B2(n_1495),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1514),
.B(n_1458),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1494),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1387),
.B(n_1515),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1412),
.A2(n_1476),
.B(n_1421),
.C(n_1500),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1486),
.B(n_1452),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1437),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1474),
.B(n_1463),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1461),
.B(n_1449),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1461),
.A2(n_1438),
.B1(n_1439),
.B2(n_1455),
.C(n_1404),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1401),
.B(n_1469),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1437),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1401),
.B(n_1469),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1454),
.A2(n_1487),
.B1(n_1431),
.B2(n_1465),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1408),
.B(n_1431),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1457),
.B(n_1431),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1449),
.B(n_1455),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1437),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1477),
.A2(n_1502),
.B(n_1491),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1474),
.B(n_1431),
.Y(n_1584)
);

OA21x2_ASAP7_75t_L g1585 ( 
.A1(n_1506),
.A2(n_1508),
.B(n_1436),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1459),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_SL g1587 ( 
.A1(n_1440),
.A2(n_1394),
.B(n_1391),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1454),
.A2(n_1509),
.B1(n_1499),
.B2(n_1391),
.Y(n_1588)
);

O2A1O1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1456),
.A2(n_1444),
.B(n_1445),
.C(n_1394),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1394),
.A2(n_1444),
.B(n_1456),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1474),
.B(n_1454),
.Y(n_1591)
);

AO21x1_ASAP7_75t_L g1592 ( 
.A1(n_1499),
.A2(n_1474),
.B(n_1405),
.Y(n_1592)
);

O2A1O1Ixp5_ASAP7_75t_L g1593 ( 
.A1(n_1499),
.A2(n_1345),
.B(n_1473),
.C(n_1222),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1505),
.A2(n_1190),
.B1(n_1057),
.B2(n_1222),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1405),
.B(n_1426),
.Y(n_1595)
);

AOI221x1_ASAP7_75t_SL g1596 ( 
.A1(n_1405),
.A2(n_1310),
.B1(n_1473),
.B2(n_1482),
.C(n_1168),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1473),
.A2(n_1222),
.B(n_1357),
.C(n_1348),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1385),
.Y(n_1598)
);

OR2x2_ASAP7_75t_SL g1599 ( 
.A(n_1466),
.B(n_899),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1393),
.A2(n_1190),
.B1(n_1057),
.B2(n_1222),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1392),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1473),
.A2(n_1222),
.B(n_1357),
.C(n_1348),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1428),
.A2(n_1357),
.B(n_1348),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1420),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1473),
.A2(n_1222),
.B(n_1293),
.C(n_1348),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1419),
.A2(n_1410),
.B(n_1467),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1393),
.A2(n_818),
.B1(n_1349),
.B2(n_1190),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_SL g1608 ( 
.A1(n_1435),
.A2(n_1203),
.B(n_1361),
.Y(n_1608)
);

OA22x2_ASAP7_75t_L g1609 ( 
.A1(n_1402),
.A2(n_1310),
.B1(n_1260),
.B2(n_1300),
.Y(n_1609)
);

O2A1O1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1473),
.A2(n_1222),
.B(n_1357),
.C(n_1348),
.Y(n_1610)
);

OA22x2_ASAP7_75t_L g1611 ( 
.A1(n_1402),
.A2(n_1310),
.B1(n_1260),
.B2(n_1300),
.Y(n_1611)
);

O2A1O1Ixp5_ASAP7_75t_L g1612 ( 
.A1(n_1473),
.A2(n_1345),
.B(n_1222),
.C(n_1467),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1380),
.B(n_1471),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1393),
.A2(n_1190),
.B1(n_1057),
.B2(n_1222),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1420),
.Y(n_1615)
);

O2A1O1Ixp5_ASAP7_75t_L g1616 ( 
.A1(n_1473),
.A2(n_1345),
.B(n_1222),
.C(n_1467),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1382),
.A2(n_1357),
.B(n_1348),
.Y(n_1617)
);

O2A1O1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1473),
.A2(n_1222),
.B(n_1357),
.C(n_1348),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1391),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1382),
.A2(n_1357),
.B(n_1348),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1517),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1587),
.B(n_1603),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1518),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1551),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1591),
.B(n_1565),
.Y(n_1625)
);

OR2x6_ASAP7_75t_L g1626 ( 
.A(n_1569),
.B(n_1526),
.Y(n_1626)
);

OR2x6_ASAP7_75t_L g1627 ( 
.A(n_1559),
.B(n_1617),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1565),
.B(n_1595),
.Y(n_1628)
);

OAI211xp5_ASAP7_75t_L g1629 ( 
.A1(n_1528),
.A2(n_1605),
.B(n_1519),
.C(n_1614),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1525),
.B(n_1522),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1532),
.B(n_1535),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1554),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1586),
.Y(n_1633)
);

OAI211xp5_ASAP7_75t_L g1634 ( 
.A1(n_1600),
.A2(n_1614),
.B(n_1597),
.C(n_1618),
.Y(n_1634)
);

INVx5_ASAP7_75t_L g1635 ( 
.A(n_1552),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1589),
.A2(n_1590),
.B(n_1620),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1567),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1545),
.Y(n_1638)
);

AO21x2_ASAP7_75t_L g1639 ( 
.A1(n_1564),
.A2(n_1550),
.B(n_1592),
.Y(n_1639)
);

AO21x2_ASAP7_75t_L g1640 ( 
.A1(n_1564),
.A2(n_1550),
.B(n_1578),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1588),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1581),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1588),
.B(n_1571),
.Y(n_1643)
);

AOI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1602),
.A2(n_1610),
.B(n_1612),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1536),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1576),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1583),
.Y(n_1647)
);

AO21x2_ASAP7_75t_L g1648 ( 
.A1(n_1547),
.A2(n_1544),
.B(n_1534),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1573),
.B(n_1530),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1547),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1544),
.B(n_1582),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1520),
.B(n_1527),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1585),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1538),
.A2(n_1593),
.B(n_1616),
.Y(n_1654)
);

AO21x2_ASAP7_75t_L g1655 ( 
.A1(n_1534),
.A2(n_1523),
.B(n_1549),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1613),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1542),
.A2(n_1606),
.B(n_1608),
.Y(n_1657)
);

OR2x6_ASAP7_75t_L g1658 ( 
.A(n_1553),
.B(n_1543),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1606),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1533),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1548),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1555),
.B(n_1541),
.Y(n_1662)
);

AO21x2_ASAP7_75t_L g1663 ( 
.A1(n_1523),
.A2(n_1549),
.B(n_1524),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1537),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1556),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1562),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1524),
.A2(n_1600),
.B(n_1611),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1540),
.A2(n_1574),
.B(n_1572),
.Y(n_1668)
);

AO21x2_ASAP7_75t_L g1669 ( 
.A1(n_1529),
.A2(n_1584),
.B(n_1594),
.Y(n_1669)
);

AO21x2_ASAP7_75t_L g1670 ( 
.A1(n_1594),
.A2(n_1546),
.B(n_1596),
.Y(n_1670)
);

CKINVDCx14_ASAP7_75t_R g1671 ( 
.A(n_1619),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1607),
.A2(n_1611),
.B1(n_1609),
.B2(n_1599),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1568),
.B(n_1539),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1672),
.B(n_1609),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1624),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1663),
.A2(n_1539),
.B1(n_1570),
.B2(n_1601),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1628),
.B(n_1566),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1672),
.B(n_1566),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1638),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1621),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1639),
.B(n_1575),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1639),
.B(n_1640),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1624),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1640),
.B(n_1577),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1640),
.B(n_1557),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1633),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1621),
.Y(n_1687)
);

OR2x6_ASAP7_75t_L g1688 ( 
.A(n_1627),
.B(n_1521),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1623),
.Y(n_1689)
);

AOI222xp33_ASAP7_75t_L g1690 ( 
.A1(n_1629),
.A2(n_1598),
.B1(n_1563),
.B2(n_1558),
.C1(n_1561),
.C2(n_1560),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1640),
.B(n_1557),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1664),
.B(n_1580),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1629),
.A2(n_1604),
.B1(n_1531),
.B2(n_1615),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1635),
.Y(n_1694)
);

NOR2xp67_ASAP7_75t_L g1695 ( 
.A(n_1635),
.B(n_1579),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1642),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1645),
.B(n_1531),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1649),
.Y(n_1698)
);

AND2x4_ASAP7_75t_SL g1699 ( 
.A(n_1622),
.B(n_1658),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1628),
.B(n_1516),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1646),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1686),
.Y(n_1702)
);

NAND3xp33_ASAP7_75t_L g1703 ( 
.A(n_1674),
.B(n_1644),
.C(n_1667),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1701),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1674),
.A2(n_1667),
.B(n_1644),
.Y(n_1705)
);

AO21x2_ASAP7_75t_L g1706 ( 
.A1(n_1682),
.A2(n_1695),
.B(n_1647),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1676),
.A2(n_1655),
.B1(n_1663),
.B2(n_1670),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1675),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1682),
.A2(n_1634),
.B1(n_1641),
.B2(n_1655),
.C(n_1663),
.Y(n_1709)
);

AOI21xp33_ASAP7_75t_L g1710 ( 
.A1(n_1690),
.A2(n_1655),
.B(n_1663),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_L g1711 ( 
.A(n_1682),
.B(n_1634),
.C(n_1627),
.Y(n_1711)
);

INVx5_ASAP7_75t_L g1712 ( 
.A(n_1688),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1698),
.B(n_1649),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1698),
.B(n_1656),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1697),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1677),
.B(n_1625),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1692),
.B(n_1666),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1676),
.A2(n_1622),
.B1(n_1626),
.B2(n_1662),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1701),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1682),
.A2(n_1655),
.B1(n_1650),
.B2(n_1652),
.C(n_1648),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1697),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1693),
.Y(n_1722)
);

NAND2xp33_ASAP7_75t_R g1723 ( 
.A(n_1694),
.B(n_1622),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_L g1724 ( 
.A(n_1690),
.B(n_1627),
.C(n_1668),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1690),
.A2(n_1622),
.B1(n_1669),
.B2(n_1648),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1686),
.Y(n_1726)
);

NAND3xp33_ASAP7_75t_SL g1727 ( 
.A(n_1693),
.B(n_1660),
.C(n_1673),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1680),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1683),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1687),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1687),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1678),
.A2(n_1670),
.B1(n_1648),
.B2(n_1622),
.Y(n_1732)
);

OAI21x1_ASAP7_75t_L g1733 ( 
.A1(n_1679),
.A2(n_1657),
.B(n_1636),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1695),
.B(n_1694),
.Y(n_1734)
);

OAI33xp33_ASAP7_75t_L g1735 ( 
.A1(n_1689),
.A2(n_1665),
.A3(n_1632),
.B1(n_1651),
.B2(n_1625),
.B3(n_1637),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1699),
.A2(n_1627),
.B(n_1626),
.Y(n_1736)
);

AOI33xp33_ASAP7_75t_L g1737 ( 
.A1(n_1685),
.A2(n_1643),
.A3(n_1661),
.B1(n_1637),
.B2(n_1630),
.B3(n_1631),
.Y(n_1737)
);

NOR3xp33_ASAP7_75t_L g1738 ( 
.A(n_1700),
.B(n_1636),
.C(n_1650),
.Y(n_1738)
);

INVx4_ASAP7_75t_L g1739 ( 
.A(n_1700),
.Y(n_1739)
);

INVx5_ASAP7_75t_L g1740 ( 
.A(n_1712),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1712),
.B(n_1695),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1734),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1702),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1722),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1734),
.B(n_1684),
.Y(n_1745)
);

OA21x2_ASAP7_75t_L g1746 ( 
.A1(n_1733),
.A2(n_1659),
.B(n_1653),
.Y(n_1746)
);

CKINVDCx16_ASAP7_75t_R g1747 ( 
.A(n_1727),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1704),
.B(n_1696),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1734),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1728),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1720),
.B(n_1654),
.C(n_1626),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1712),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1702),
.Y(n_1753)
);

AND2x6_ASAP7_75t_SL g1754 ( 
.A(n_1714),
.B(n_1658),
.Y(n_1754)
);

INVx4_ASAP7_75t_SL g1755 ( 
.A(n_1719),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1706),
.B(n_1684),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1726),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1730),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1709),
.B(n_1694),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1706),
.B(n_1684),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1731),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1716),
.B(n_1708),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1739),
.B(n_1685),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1713),
.Y(n_1764)
);

INVx2_ASAP7_75t_SL g1765 ( 
.A(n_1712),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1750),
.Y(n_1766)
);

AND2x4_ASAP7_75t_SL g1767 ( 
.A(n_1741),
.B(n_1658),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1764),
.B(n_1737),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1750),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1740),
.B(n_1738),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1758),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1756),
.B(n_1760),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1740),
.B(n_1685),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1756),
.B(n_1685),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1756),
.B(n_1691),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1760),
.B(n_1691),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1740),
.B(n_1691),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1746),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1758),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1760),
.B(n_1691),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1747),
.B(n_1705),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1740),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1740),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1746),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1745),
.B(n_1737),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1746),
.Y(n_1786)
);

AND2x4_ASAP7_75t_SL g1787 ( 
.A(n_1741),
.B(n_1658),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1764),
.B(n_1721),
.Y(n_1788)
);

A2O1A1Ixp33_ASAP7_75t_L g1789 ( 
.A1(n_1751),
.A2(n_1703),
.B(n_1711),
.C(n_1710),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1761),
.Y(n_1790)
);

INVx3_ASAP7_75t_R g1791 ( 
.A(n_1742),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1762),
.B(n_1729),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1754),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1743),
.B(n_1715),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1762),
.B(n_1729),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1740),
.B(n_1679),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1741),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1761),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1757),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1762),
.B(n_1717),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1746),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1757),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1740),
.B(n_1679),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1788),
.B(n_1759),
.Y(n_1804)
);

OAI21xp33_ASAP7_75t_L g1805 ( 
.A1(n_1781),
.A2(n_1751),
.B(n_1759),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1785),
.B(n_1742),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1789),
.B(n_1747),
.Y(n_1807)
);

NOR2xp67_ASAP7_75t_L g1808 ( 
.A(n_1782),
.B(n_1749),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1793),
.A2(n_1732),
.B1(n_1707),
.B2(n_1725),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1799),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1768),
.B(n_1743),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1768),
.B(n_1753),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1793),
.B(n_1740),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1799),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1785),
.B(n_1742),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1770),
.A2(n_1724),
.B(n_1707),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1766),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1766),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1769),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1785),
.B(n_1749),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1772),
.B(n_1749),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1800),
.B(n_1753),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1788),
.B(n_1744),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1794),
.B(n_1722),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1800),
.B(n_1748),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1794),
.B(n_1763),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1792),
.Y(n_1827)
);

AOI21xp33_ASAP7_75t_L g1828 ( 
.A1(n_1770),
.A2(n_1765),
.B(n_1752),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1802),
.B(n_1763),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1769),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1771),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1800),
.B(n_1748),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1791),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1802),
.B(n_1681),
.Y(n_1834)
);

INVxp67_ASAP7_75t_L g1835 ( 
.A(n_1771),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1772),
.B(n_1755),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1779),
.B(n_1681),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1779),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1767),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1772),
.B(n_1755),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1811),
.B(n_1790),
.Y(n_1841)
);

INVx2_ASAP7_75t_SL g1842 ( 
.A(n_1821),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1833),
.B(n_1790),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1807),
.B(n_1798),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1805),
.A2(n_1732),
.B1(n_1718),
.B2(n_1787),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1823),
.B(n_1671),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1810),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1824),
.B(n_1798),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1839),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1817),
.Y(n_1850)
);

INVx4_ASAP7_75t_L g1851 ( 
.A(n_1813),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1806),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1806),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1836),
.B(n_1797),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1836),
.B(n_1797),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1818),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1821),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1819),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1811),
.B(n_1792),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1814),
.B(n_1774),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1840),
.B(n_1797),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1820),
.B(n_1774),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1840),
.B(n_1797),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1838),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1830),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1813),
.B(n_1797),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1853),
.B(n_1835),
.Y(n_1867)
);

OAI32xp33_ASAP7_75t_L g1868 ( 
.A1(n_1852),
.A2(n_1804),
.A3(n_1809),
.B1(n_1816),
.B2(n_1812),
.Y(n_1868)
);

AOI222xp33_ASAP7_75t_L g1869 ( 
.A1(n_1844),
.A2(n_1815),
.B1(n_1813),
.B2(n_1820),
.C1(n_1831),
.C2(n_1735),
.Y(n_1869)
);

A2O1A1Ixp33_ASAP7_75t_L g1870 ( 
.A1(n_1845),
.A2(n_1812),
.B(n_1815),
.C(n_1828),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1859),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1849),
.A2(n_1787),
.B1(n_1767),
.B2(n_1808),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1846),
.B(n_1851),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1866),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1859),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1854),
.Y(n_1876)
);

AOI221xp5_ASAP7_75t_L g1877 ( 
.A1(n_1843),
.A2(n_1829),
.B1(n_1826),
.B2(n_1834),
.C(n_1770),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1841),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1857),
.B(n_1842),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1860),
.B(n_1822),
.Y(n_1880)
);

AOI211xp5_ASAP7_75t_L g1881 ( 
.A1(n_1848),
.A2(n_1770),
.B(n_1822),
.C(n_1783),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1851),
.B(n_1825),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1841),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1854),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1842),
.B(n_1827),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1857),
.A2(n_1767),
.B1(n_1787),
.B2(n_1773),
.Y(n_1886)
);

AOI222xp33_ASAP7_75t_L g1887 ( 
.A1(n_1868),
.A2(n_1847),
.B1(n_1865),
.B2(n_1864),
.C1(n_1856),
.C2(n_1850),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1871),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1875),
.B(n_1847),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1876),
.B(n_1855),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1878),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1884),
.B(n_1855),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1883),
.B(n_1850),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1873),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1880),
.B(n_1862),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1874),
.B(n_1851),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1879),
.B(n_1861),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1885),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1867),
.B(n_1825),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1889),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1887),
.A2(n_1870),
.B(n_1869),
.Y(n_1901)
);

NAND3xp33_ASAP7_75t_SL g1902 ( 
.A(n_1887),
.B(n_1869),
.C(n_1881),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1897),
.B(n_1882),
.Y(n_1903)
);

OAI31xp33_ASAP7_75t_L g1904 ( 
.A1(n_1896),
.A2(n_1867),
.A3(n_1863),
.B(n_1861),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1890),
.B(n_1892),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1899),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1894),
.A2(n_1872),
.B1(n_1886),
.B2(n_1863),
.Y(n_1907)
);

OAI22xp33_ASAP7_75t_SL g1908 ( 
.A1(n_1888),
.A2(n_1783),
.B1(n_1782),
.B2(n_1858),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1898),
.B(n_1877),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1889),
.A2(n_1858),
.B(n_1783),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1905),
.Y(n_1911)
);

A2O1A1Ixp33_ASAP7_75t_SL g1912 ( 
.A1(n_1901),
.A2(n_1891),
.B(n_1893),
.C(n_1782),
.Y(n_1912)
);

XNOR2xp5_ASAP7_75t_L g1913 ( 
.A(n_1907),
.B(n_1895),
.Y(n_1913)
);

A2O1A1Ixp33_ASAP7_75t_L g1914 ( 
.A1(n_1902),
.A2(n_1893),
.B(n_1770),
.C(n_1783),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_SL g1915 ( 
.A(n_1900),
.Y(n_1915)
);

AOI322xp5_ASAP7_75t_L g1916 ( 
.A1(n_1902),
.A2(n_1909),
.A3(n_1906),
.B1(n_1903),
.B2(n_1775),
.C1(n_1780),
.C2(n_1776),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1916),
.B(n_1904),
.Y(n_1917)
);

NOR3xp33_ASAP7_75t_L g1918 ( 
.A(n_1911),
.B(n_1908),
.C(n_1910),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1915),
.Y(n_1919)
);

XNOR2xp5_ASAP7_75t_L g1920 ( 
.A(n_1913),
.B(n_1782),
.Y(n_1920)
);

INVx1_ASAP7_75t_SL g1921 ( 
.A(n_1912),
.Y(n_1921)
);

OAI21xp33_ASAP7_75t_SL g1922 ( 
.A1(n_1914),
.A2(n_1827),
.B(n_1791),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1911),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1919),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1923),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1921),
.B(n_1918),
.Y(n_1926)
);

NAND2xp33_ASAP7_75t_SL g1927 ( 
.A(n_1920),
.B(n_1832),
.Y(n_1927)
);

AND4x2_ASAP7_75t_L g1928 ( 
.A(n_1922),
.B(n_1736),
.C(n_1832),
.D(n_1754),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1917),
.A2(n_1837),
.B(n_1803),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1924),
.Y(n_1930)
);

NAND4xp25_ASAP7_75t_L g1931 ( 
.A(n_1926),
.B(n_1752),
.C(n_1773),
.D(n_1777),
.Y(n_1931)
);

XNOR2xp5_ASAP7_75t_L g1932 ( 
.A(n_1927),
.B(n_1752),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1930),
.B(n_1925),
.Y(n_1933)
);

AOI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1933),
.A2(n_1932),
.B1(n_1931),
.B2(n_1929),
.C(n_1928),
.Y(n_1934)
);

NOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1934),
.B(n_1752),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1934),
.Y(n_1936)
);

OAI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1935),
.A2(n_1936),
.B(n_1803),
.Y(n_1937)
);

OAI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1936),
.A2(n_1795),
.B1(n_1792),
.B2(n_1803),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1937),
.Y(n_1939)
);

OAI321xp33_ASAP7_75t_L g1940 ( 
.A1(n_1938),
.A2(n_1765),
.A3(n_1784),
.B1(n_1786),
.B2(n_1778),
.C(n_1801),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1939),
.B(n_1803),
.Y(n_1941)
);

AO21x2_ASAP7_75t_L g1942 ( 
.A1(n_1941),
.A2(n_1940),
.B(n_1784),
.Y(n_1942)
);

OAI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1942),
.A2(n_1803),
.B(n_1796),
.Y(n_1943)
);

OAI221xp5_ASAP7_75t_R g1944 ( 
.A1(n_1943),
.A2(n_1723),
.B1(n_1778),
.B2(n_1784),
.C(n_1801),
.Y(n_1944)
);

OAI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1944),
.A2(n_1778),
.B1(n_1786),
.B2(n_1801),
.Y(n_1945)
);

AOI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1945),
.A2(n_1796),
.B(n_1786),
.C(n_1773),
.Y(n_1946)
);


endmodule