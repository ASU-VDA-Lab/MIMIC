module real_aes_2631_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g531 ( .A(n_0), .B(n_228), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_1), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g162 ( .A(n_2), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_3), .B(n_534), .Y(n_553) );
NAND2xp33_ASAP7_75t_SL g524 ( .A(n_4), .B(n_183), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_5), .B(n_196), .Y(n_219) );
INVx1_ASAP7_75t_L g516 ( .A(n_6), .Y(n_516) );
INVx1_ASAP7_75t_L g253 ( .A(n_7), .Y(n_253) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_8), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_9), .Y(n_270) );
AND2x2_ASAP7_75t_L g551 ( .A(n_10), .B(n_152), .Y(n_551) );
INVx2_ASAP7_75t_L g153 ( .A(n_11), .Y(n_153) );
AND3x1_ASAP7_75t_L g111 ( .A(n_12), .B(n_34), .C(n_112), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g125 ( .A(n_12), .Y(n_125) );
INVx1_ASAP7_75t_L g229 ( .A(n_13), .Y(n_229) );
AOI221x1_ASAP7_75t_L g519 ( .A1(n_14), .A2(n_185), .B1(n_520), .B2(n_522), .C(n_523), .Y(n_519) );
OAI22xp5_ASAP7_75t_SL g805 ( .A1(n_14), .A2(n_58), .B1(n_806), .B2(n_807), .Y(n_805) );
INVxp67_ASAP7_75t_L g807 ( .A(n_14), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_15), .B(n_534), .Y(n_587) );
INVx1_ASAP7_75t_L g110 ( .A(n_16), .Y(n_110) );
INVx1_ASAP7_75t_L g226 ( .A(n_17), .Y(n_226) );
INVx1_ASAP7_75t_SL g174 ( .A(n_18), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_19), .B(n_177), .Y(n_199) );
AOI33xp33_ASAP7_75t_L g244 ( .A1(n_20), .A2(n_48), .A3(n_159), .B1(n_170), .B2(n_245), .B3(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_21), .A2(n_522), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_22), .B(n_228), .Y(n_556) );
AOI221xp5_ASAP7_75t_SL g596 ( .A1(n_23), .A2(n_39), .B1(n_522), .B2(n_534), .C(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g263 ( .A(n_24), .Y(n_263) );
OR2x2_ASAP7_75t_L g154 ( .A(n_25), .B(n_93), .Y(n_154) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_25), .A2(n_93), .B(n_153), .Y(n_187) );
INVxp67_ASAP7_75t_L g518 ( .A(n_26), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_27), .B(n_231), .Y(n_591) );
AND2x2_ASAP7_75t_L g545 ( .A(n_28), .B(n_151), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_29), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_30), .B(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_31), .A2(n_522), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_32), .B(n_231), .Y(n_598) );
AND2x2_ASAP7_75t_L g164 ( .A(n_33), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g169 ( .A(n_33), .Y(n_169) );
AND2x2_ASAP7_75t_L g183 ( .A(n_33), .B(n_162), .Y(n_183) );
OR2x6_ASAP7_75t_L g126 ( .A(n_34), .B(n_127), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_35), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_36), .B(n_157), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_37), .A2(n_186), .B1(n_192), .B2(n_196), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_38), .B(n_201), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_40), .A2(n_85), .B1(n_167), .B2(n_522), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_41), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_42), .B(n_228), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_43), .B(n_203), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_44), .B(n_177), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_45), .Y(n_195) );
AND2x2_ASAP7_75t_L g535 ( .A(n_46), .B(n_151), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_47), .B(n_151), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_49), .B(n_177), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_50), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_50), .A2(n_63), .B1(n_442), .B2(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_51), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g160 ( .A(n_52), .Y(n_160) );
INVx1_ASAP7_75t_L g179 ( .A(n_52), .Y(n_179) );
AOI22x1_ASAP7_75t_L g132 ( .A1(n_53), .A2(n_133), .B1(n_134), .B2(n_135), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_53), .Y(n_133) );
AND2x2_ASAP7_75t_L g295 ( .A(n_54), .B(n_151), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_55), .A2(n_77), .B1(n_157), .B2(n_167), .C(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_56), .B(n_157), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_57), .B(n_534), .Y(n_544) );
INVx1_ASAP7_75t_L g806 ( .A(n_58), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_59), .B(n_186), .Y(n_272) );
AOI21xp5_ASAP7_75t_SL g208 ( .A1(n_60), .A2(n_167), .B(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g572 ( .A(n_61), .B(n_151), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_62), .B(n_231), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_63), .Y(n_818) );
INVx1_ASAP7_75t_L g222 ( .A(n_64), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_65), .B(n_228), .Y(n_570) );
AND2x2_ASAP7_75t_SL g592 ( .A(n_66), .B(n_152), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_67), .A2(n_522), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g293 ( .A(n_68), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_69), .B(n_231), .Y(n_557) );
AND2x2_ASAP7_75t_SL g564 ( .A(n_70), .B(n_203), .Y(n_564) );
XOR2xp5_ASAP7_75t_L g131 ( .A(n_71), .B(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_72), .A2(n_104), .B1(n_136), .B2(n_137), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_72), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_73), .A2(n_167), .B(n_292), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_74), .A2(n_816), .B1(n_817), .B2(n_819), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_74), .Y(n_816) );
INVx1_ASAP7_75t_L g165 ( .A(n_75), .Y(n_165) );
INVx1_ASAP7_75t_L g181 ( .A(n_75), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_76), .B(n_157), .Y(n_247) );
AND2x2_ASAP7_75t_L g184 ( .A(n_78), .B(n_185), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_79), .A2(n_106), .B1(n_115), .B2(n_828), .Y(n_105) );
INVx1_ASAP7_75t_L g223 ( .A(n_80), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_81), .A2(n_167), .B(n_173), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_82), .A2(n_167), .B(n_198), .C(n_202), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_83), .A2(n_88), .B1(n_157), .B2(n_534), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_84), .B(n_534), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_86), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g128 ( .A(n_86), .Y(n_128) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_87), .B(n_185), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_89), .A2(n_167), .B1(n_242), .B2(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_90), .B(n_228), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_91), .B(n_228), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_92), .A2(n_522), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g210 ( .A(n_94), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_95), .B(n_231), .Y(n_569) );
AND2x2_ASAP7_75t_L g248 ( .A(n_96), .B(n_185), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_97), .A2(n_261), .B(n_262), .C(n_264), .Y(n_260) );
INVxp67_ASAP7_75t_L g521 ( .A(n_98), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_99), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_100), .B(n_231), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_101), .A2(n_522), .B(n_589), .Y(n_588) );
BUFx2_ASAP7_75t_L g120 ( .A(n_102), .Y(n_120) );
INVx1_ASAP7_75t_SL g803 ( .A(n_102), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_103), .B(n_177), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_104), .Y(n_137) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g829 ( .A(n_107), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_111), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_110), .B(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_801), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_129), .Y(n_121) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
AND2x6_ASAP7_75t_SL g506 ( .A(n_125), .B(n_126), .Y(n_506) );
OR2x6_ASAP7_75t_SL g797 ( .A(n_125), .B(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_125), .B(n_798), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_126), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B1(n_138), .B2(n_799), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22x1_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_505), .B1(n_507), .B2(n_795), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_140), .A2(n_505), .B1(n_508), .B2(n_800), .Y(n_799) );
AND3x1_ASAP7_75t_L g140 ( .A(n_141), .B(n_499), .C(n_502), .Y(n_140) );
NAND5xp2_ASAP7_75t_L g141 ( .A(n_142), .B(n_399), .C(n_429), .D(n_443), .E(n_469), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OAI21xp33_ASAP7_75t_L g499 ( .A1(n_143), .A2(n_442), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g812 ( .A(n_143), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_348), .Y(n_143) );
NOR3xp33_ASAP7_75t_SL g144 ( .A(n_145), .B(n_296), .C(n_330), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_213), .B(n_235), .C(n_274), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_188), .Y(n_146) );
BUFx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_148), .B(n_286), .Y(n_351) );
AND2x2_ASAP7_75t_L g438 ( .A(n_148), .B(n_216), .Y(n_438) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g234 ( .A(n_149), .B(n_205), .Y(n_234) );
INVx1_ASAP7_75t_L g276 ( .A(n_149), .Y(n_276) );
INVx2_ASAP7_75t_L g281 ( .A(n_149), .Y(n_281) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_149), .Y(n_309) );
INVx1_ASAP7_75t_L g323 ( .A(n_149), .Y(n_323) );
AND2x2_ASAP7_75t_L g327 ( .A(n_149), .B(n_218), .Y(n_327) );
AND2x2_ASAP7_75t_L g408 ( .A(n_149), .B(n_217), .Y(n_408) );
AO21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_155), .B(n_184), .Y(n_149) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_150), .A2(n_539), .B(n_545), .Y(n_538) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_150), .A2(n_566), .B(n_572), .Y(n_565) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_150), .A2(n_539), .B(n_545), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_151), .Y(n_150) );
OA21x2_ASAP7_75t_L g595 ( .A1(n_151), .A2(n_596), .B(n_600), .Y(n_595) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x4_ASAP7_75t_L g196 ( .A(n_153), .B(n_154), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_166), .Y(n_155) );
INVx1_ASAP7_75t_L g273 ( .A(n_157), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_157), .A2(n_167), .B1(n_515), .B2(n_517), .Y(n_514) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_163), .Y(n_157) );
INVx1_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_161), .Y(n_158) );
OR2x6_ASAP7_75t_L g175 ( .A(n_159), .B(n_171), .Y(n_175) );
INVxp33_ASAP7_75t_L g245 ( .A(n_159), .Y(n_245) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g172 ( .A(n_160), .B(n_162), .Y(n_172) );
AND2x4_ASAP7_75t_L g231 ( .A(n_160), .B(n_180), .Y(n_231) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x6_ASAP7_75t_L g522 ( .A(n_164), .B(n_172), .Y(n_522) );
INVx2_ASAP7_75t_L g171 ( .A(n_165), .Y(n_171) );
AND2x6_ASAP7_75t_L g228 ( .A(n_165), .B(n_178), .Y(n_228) );
INVxp67_ASAP7_75t_L g271 ( .A(n_167), .Y(n_271) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_172), .Y(n_167) );
NOR2x1p5_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
INVx1_ASAP7_75t_L g246 ( .A(n_170), .Y(n_246) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_182), .Y(n_173) );
INVx2_ASAP7_75t_L g201 ( .A(n_175), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_175), .A2(n_182), .B(n_210), .C(n_211), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_175), .A2(n_222), .B1(n_223), .B2(n_224), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_SL g252 ( .A1(n_175), .A2(n_182), .B(n_253), .C(n_254), .Y(n_252) );
INVxp67_ASAP7_75t_L g261 ( .A(n_175), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g292 ( .A1(n_175), .A2(n_182), .B(n_293), .C(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g224 ( .A(n_177), .Y(n_224) );
AND2x4_ASAP7_75t_L g534 ( .A(n_177), .B(n_183), .Y(n_534) );
AND2x4_ASAP7_75t_L g177 ( .A(n_178), .B(n_180), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_182), .A2(n_199), .B(n_200), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_182), .B(n_196), .Y(n_232) );
INVx1_ASAP7_75t_L g242 ( .A(n_182), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_182), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_182), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_182), .A2(n_556), .B(n_557), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_182), .A2(n_569), .B(n_570), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_182), .A2(n_590), .B(n_591), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_182), .A2(n_598), .B(n_599), .Y(n_597) );
INVx5_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_183), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_185), .A2(n_260), .B1(n_265), .B2(n_266), .Y(n_259) );
INVx3_ASAP7_75t_L g266 ( .A(n_185), .Y(n_266) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_186), .B(n_269), .Y(n_268) );
AOI21x1_ASAP7_75t_L g527 ( .A1(n_186), .A2(n_528), .B(n_535), .Y(n_527) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx4f_ASAP7_75t_L g203 ( .A(n_187), .Y(n_203) );
AND2x4_ASAP7_75t_SL g188 ( .A(n_189), .B(n_204), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g233 ( .A(n_190), .Y(n_233) );
AND2x2_ASAP7_75t_L g277 ( .A(n_190), .B(n_218), .Y(n_277) );
AND2x2_ASAP7_75t_L g298 ( .A(n_190), .B(n_205), .Y(n_298) );
INVx1_ASAP7_75t_L g321 ( .A(n_190), .Y(n_321) );
AND2x4_ASAP7_75t_L g388 ( .A(n_190), .B(n_217), .Y(n_388) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_197), .Y(n_190) );
NOR3xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .C(n_195), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_196), .A2(n_208), .B(n_212), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_196), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_196), .B(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_196), .B(n_521), .Y(n_520) );
NOR3xp33_ASAP7_75t_L g523 ( .A(n_196), .B(n_224), .C(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_196), .A2(n_553), .B(n_554), .Y(n_552) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_202), .A2(n_240), .B(n_248), .Y(n_239) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_202), .A2(n_240), .B(n_248), .Y(n_303) );
AOI21x1_ASAP7_75t_L g560 ( .A1(n_202), .A2(n_561), .B(n_564), .Y(n_560) );
INVx2_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_203), .A2(n_251), .B(n_255), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_203), .A2(n_587), .B(n_588), .Y(n_586) );
AND2x4_ASAP7_75t_L g404 ( .A(n_204), .B(n_321), .Y(n_404) );
OR2x2_ASAP7_75t_L g445 ( .A(n_204), .B(n_446), .Y(n_445) );
NOR2xp67_ASAP7_75t_SL g464 ( .A(n_204), .B(n_337), .Y(n_464) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_204), .B(n_396), .Y(n_482) );
INVx4_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2x1_ASAP7_75t_SL g282 ( .A(n_205), .B(n_218), .Y(n_282) );
AND2x4_ASAP7_75t_L g320 ( .A(n_205), .B(n_321), .Y(n_320) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_205), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_205), .B(n_280), .Y(n_358) );
INVx2_ASAP7_75t_L g372 ( .A(n_205), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_205), .B(n_324), .Y(n_394) );
AND2x2_ASAP7_75t_L g486 ( .A(n_205), .B(n_344), .Y(n_486) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2x1_ASAP7_75t_L g214 ( .A(n_215), .B(n_234), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_216), .B(n_323), .Y(n_337) );
AND2x2_ASAP7_75t_SL g346 ( .A(n_216), .B(n_326), .Y(n_346) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_233), .Y(n_216) );
INVx1_ASAP7_75t_L g324 ( .A(n_217), .Y(n_324) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g344 ( .A(n_218), .Y(n_344) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_225), .B(n_232), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_224), .B(n_263), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B1(n_229), .B2(n_230), .Y(n_225) );
INVxp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g377 ( .A(n_233), .Y(n_377) );
INVx2_ASAP7_75t_SL g422 ( .A(n_234), .Y(n_422) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_256), .Y(n_236) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_237), .B(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g368 ( .A(n_237), .Y(n_368) );
AND2x2_ASAP7_75t_L g492 ( .A(n_237), .B(n_317), .Y(n_492) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_249), .Y(n_237) );
AND2x4_ASAP7_75t_L g305 ( .A(n_238), .B(n_287), .Y(n_305) );
INVx1_ASAP7_75t_L g316 ( .A(n_238), .Y(n_316) );
AND2x2_ASAP7_75t_L g347 ( .A(n_238), .B(n_302), .Y(n_347) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_239), .B(n_250), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_239), .B(n_288), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_241), .B(n_247), .Y(n_240) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g285 ( .A(n_250), .Y(n_285) );
AND2x4_ASAP7_75t_L g353 ( .A(n_250), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g365 ( .A(n_250), .Y(n_365) );
INVx1_ASAP7_75t_L g407 ( .A(n_250), .Y(n_407) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_250), .Y(n_419) );
AND2x2_ASAP7_75t_L g435 ( .A(n_250), .B(n_258), .Y(n_435) );
BUFx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g382 ( .A(n_257), .B(n_340), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_257), .Y(n_384) );
AND2x2_ASAP7_75t_L g405 ( .A(n_257), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g284 ( .A(n_258), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g312 ( .A(n_258), .Y(n_312) );
INVx2_ASAP7_75t_L g318 ( .A(n_258), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_258), .B(n_288), .Y(n_333) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_267), .Y(n_258) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_266), .A2(n_289), .B(n_295), .Y(n_288) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_266), .A2(n_289), .B(n_295), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B1(n_272), .B2(n_273), .Y(n_267) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI21xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_278), .B(n_283), .Y(n_274) );
INVx1_ASAP7_75t_L g414 ( .A(n_275), .Y(n_414) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx2_ASAP7_75t_L g334 ( .A(n_277), .Y(n_334) );
AND2x2_ASAP7_75t_L g390 ( .A(n_277), .B(n_326), .Y(n_390) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
INVx1_ASAP7_75t_L g304 ( .A(n_279), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_279), .B(n_320), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_279), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g411 ( .A(n_279), .B(n_404), .Y(n_411) );
AND2x2_ASAP7_75t_L g485 ( .A(n_279), .B(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_280), .Y(n_473) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_281), .Y(n_393) );
AND2x2_ASAP7_75t_L g306 ( .A(n_282), .B(n_307), .Y(n_306) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_282), .A2(n_495), .B(n_497), .Y(n_494) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx3_ASAP7_75t_L g380 ( .A(n_284), .Y(n_380) );
NAND2x1_ASAP7_75t_SL g424 ( .A(n_284), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g427 ( .A(n_284), .B(n_305), .Y(n_427) );
AND2x2_ASAP7_75t_L g339 ( .A(n_286), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g476 ( .A(n_286), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g487 ( .A(n_286), .B(n_435), .Y(n_487) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_287), .B(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g418 ( .A(n_288), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
OAI21xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_310), .B(n_313), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_305), .B2(n_306), .Y(n_297) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_298), .Y(n_355) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_304), .Y(n_299) );
AND2x2_ASAP7_75t_L g328 ( .A(n_300), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g434 ( .A(n_300), .B(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_300), .A2(n_453), .B1(n_454), .B2(n_455), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_300), .B(n_461), .Y(n_460) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g317 ( .A(n_302), .B(n_318), .Y(n_317) );
NOR2xp67_ASAP7_75t_L g398 ( .A(n_302), .B(n_318), .Y(n_398) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_302), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g354 ( .A(n_303), .Y(n_354) );
AND2x2_ASAP7_75t_L g362 ( .A(n_303), .B(n_318), .Y(n_362) );
INVx1_ASAP7_75t_L g425 ( .A(n_303), .Y(n_425) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2x1_ASAP7_75t_L g343 ( .A(n_308), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g455 ( .A(n_311), .B(n_340), .Y(n_455) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g329 ( .A(n_312), .Y(n_329) );
AND2x2_ASAP7_75t_L g352 ( .A(n_312), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g440 ( .A(n_312), .B(n_347), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_319), .B1(n_325), .B2(n_328), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g448 ( .A(n_315), .B(n_449), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g478 ( .A(n_318), .B(n_365), .Y(n_478) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx2_ASAP7_75t_L g345 ( .A(n_320), .Y(n_345) );
OAI21xp33_ASAP7_75t_SL g491 ( .A1(n_320), .A2(n_492), .B(n_493), .Y(n_491) );
AND2x4_ASAP7_75t_SL g322 ( .A(n_323), .B(n_324), .Y(n_322) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_323), .Y(n_481) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_SL g423 ( .A1(n_326), .A2(n_424), .B(n_426), .C(n_428), .Y(n_423) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_327), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g428 ( .A(n_327), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_327), .B(n_404), .Y(n_468) );
INVx1_ASAP7_75t_SL g335 ( .A(n_328), .Y(n_335) );
AND2x2_ASAP7_75t_L g416 ( .A(n_329), .B(n_353), .Y(n_416) );
INVx1_ASAP7_75t_L g461 ( .A(n_329), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B1(n_335), .B2(n_336), .C(n_338), .Y(n_330) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_331), .Y(n_450) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g498 ( .A(n_333), .B(n_341), .Y(n_498) );
OR2x2_ASAP7_75t_L g357 ( .A(n_334), .B(n_358), .Y(n_357) );
NOR2x1_ASAP7_75t_L g370 ( .A(n_334), .B(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_334), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g496 ( .A(n_334), .B(n_393), .Y(n_496) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI32xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .A3(n_345), .B1(n_346), .B2(n_347), .Y(n_338) );
INVx1_ASAP7_75t_L g359 ( .A(n_340), .Y(n_359) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_342), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g454 ( .A(n_343), .Y(n_454) );
OAI22xp33_ASAP7_75t_SL g436 ( .A1(n_345), .A2(n_437), .B1(n_439), .B2(n_441), .Y(n_436) );
INVx1_ASAP7_75t_L g467 ( .A(n_346), .Y(n_467) );
AOI211x1_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_355), .B(n_356), .C(n_373), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_350), .B(n_435), .Y(n_441) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g397 ( .A(n_353), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g463 ( .A(n_353), .Y(n_463) );
OAI222xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B1(n_360), .B2(n_366), .C1(n_367), .C2(n_369), .Y(n_356) );
INVxp67_ASAP7_75t_L g453 ( .A(n_357), .Y(n_453) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_361), .B(n_446), .Y(n_493) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g409 ( .A(n_362), .B(n_406), .Y(n_409) );
INVx3_ASAP7_75t_L g449 ( .A(n_364), .Y(n_449) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g387 ( .A(n_372), .B(n_388), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B1(n_381), .B2(n_386), .C(n_389), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_375), .A2(n_432), .B(n_434), .Y(n_431) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g385 ( .A(n_379), .Y(n_385) );
OR2x2_ASAP7_75t_L g489 ( .A(n_380), .B(n_425), .Y(n_489) );
NOR2xp67_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_383), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_386), .A2(n_415), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_387), .A2(n_459), .B(n_466), .Y(n_465) );
INVx4_ASAP7_75t_L g396 ( .A(n_388), .Y(n_396) );
OAI31xp33_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_391), .A3(n_395), .B(n_397), .Y(n_389) );
INVx1_ASAP7_75t_L g447 ( .A(n_391), .Y(n_447) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g421 ( .A(n_396), .Y(n_421) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_412), .Y(n_399) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_400), .B(n_412), .C(n_431), .D(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_410), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B1(n_408), .B2(n_409), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g472 ( .A(n_404), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_405), .B(n_425), .Y(n_433) );
INVx1_ASAP7_75t_SL g446 ( .A(n_408), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_423), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_417), .B2(n_420), .Y(n_413) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2x1_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_422), .A2(n_485), .B1(n_487), .B2(n_488), .Y(n_484) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NOR3xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_436), .C(n_442), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g501 ( .A(n_436), .Y(n_501) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI21xp33_ASAP7_75t_L g502 ( .A1(n_442), .A2(n_503), .B(n_504), .Y(n_502) );
INVxp33_ASAP7_75t_L g503 ( .A(n_443), .Y(n_503) );
AND2x2_ASAP7_75t_L g811 ( .A(n_443), .B(n_469), .Y(n_811) );
NOR2xp67_ASAP7_75t_L g443 ( .A(n_444), .B(n_451), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_447), .B1(n_448), .B2(n_450), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_448), .A2(n_471), .B(n_474), .Y(n_470) );
INVx2_ASAP7_75t_L g458 ( .A(n_449), .Y(n_458) );
NAND3xp33_ASAP7_75t_SL g451 ( .A(n_452), .B(n_456), .C(n_465), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_462), .B2(n_464), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVxp33_ASAP7_75t_SL g504 ( .A(n_469), .Y(n_504) );
NOR3x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_483), .C(n_490), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_491), .B(n_494), .Y(n_490) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g813 ( .A(n_500), .Y(n_813) );
CKINVDCx11_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_672), .Y(n_508) );
NOR4xp25_ASAP7_75t_L g509 ( .A(n_510), .B(n_615), .C(n_654), .D(n_661), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_536), .B1(n_573), .B2(n_582), .C(n_601), .Y(n_510) );
OR2x2_ASAP7_75t_L g745 ( .A(n_511), .B(n_607), .Y(n_745) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g660 ( .A(n_512), .B(n_585), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_512), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_SL g725 ( .A(n_512), .B(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_525), .Y(n_512) );
AND2x4_ASAP7_75t_SL g584 ( .A(n_513), .B(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g606 ( .A(n_513), .Y(n_606) );
AND2x2_ASAP7_75t_L g641 ( .A(n_513), .B(n_614), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_513), .B(n_526), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_513), .B(n_608), .Y(n_693) );
OR2x2_ASAP7_75t_L g771 ( .A(n_513), .B(n_585), .Y(n_771) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .Y(n_513) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g593 ( .A(n_526), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_526), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g619 ( .A(n_526), .Y(n_619) );
OR2x2_ASAP7_75t_L g624 ( .A(n_526), .B(n_608), .Y(n_624) );
AND2x2_ASAP7_75t_L g637 ( .A(n_526), .B(n_595), .Y(n_637) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_526), .Y(n_640) );
INVx1_ASAP7_75t_L g652 ( .A(n_526), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_526), .B(n_606), .Y(n_717) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_537), .B(n_546), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g581 ( .A(n_538), .B(n_565), .Y(n_581) );
AND2x4_ASAP7_75t_L g611 ( .A(n_538), .B(n_550), .Y(n_611) );
INVx2_ASAP7_75t_L g645 ( .A(n_538), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_538), .B(n_565), .Y(n_703) );
AND2x2_ASAP7_75t_L g750 ( .A(n_538), .B(n_579), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_544), .Y(n_539) );
AOI222xp33_ASAP7_75t_L g738 ( .A1(n_546), .A2(n_610), .B1(n_653), .B2(n_713), .C1(n_739), .C2(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_558), .Y(n_547) );
AND2x2_ASAP7_75t_L g657 ( .A(n_548), .B(n_577), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_548), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g786 ( .A(n_548), .B(n_626), .Y(n_786) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_549), .A2(n_617), .B(n_621), .Y(n_616) );
AND2x2_ASAP7_75t_L g697 ( .A(n_549), .B(n_580), .Y(n_697) );
OR2x2_ASAP7_75t_L g722 ( .A(n_549), .B(n_581), .Y(n_722) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx5_ASAP7_75t_L g576 ( .A(n_550), .Y(n_576) );
AND2x2_ASAP7_75t_L g663 ( .A(n_550), .B(n_645), .Y(n_663) );
AND2x2_ASAP7_75t_L g689 ( .A(n_550), .B(n_565), .Y(n_689) );
OR2x2_ASAP7_75t_L g692 ( .A(n_550), .B(n_579), .Y(n_692) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_550), .Y(n_710) );
AND2x4_ASAP7_75t_SL g767 ( .A(n_550), .B(n_644), .Y(n_767) );
OR2x2_ASAP7_75t_L g776 ( .A(n_550), .B(n_603), .Y(n_776) );
OR2x6_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g609 ( .A(n_558), .Y(n_609) );
AOI221xp5_ASAP7_75t_SL g727 ( .A1(n_558), .A2(n_611), .B1(n_728), .B2(n_730), .C(n_731), .Y(n_727) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_565), .Y(n_558) );
OR2x2_ASAP7_75t_L g666 ( .A(n_559), .B(n_636), .Y(n_666) );
OR2x2_ASAP7_75t_L g676 ( .A(n_559), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g702 ( .A(n_559), .B(n_703), .Y(n_702) );
AND2x4_ASAP7_75t_L g708 ( .A(n_559), .B(n_627), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_559), .B(n_691), .Y(n_720) );
INVx2_ASAP7_75t_L g733 ( .A(n_559), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_559), .B(n_611), .Y(n_754) );
AND2x2_ASAP7_75t_L g758 ( .A(n_559), .B(n_580), .Y(n_758) );
AND2x2_ASAP7_75t_L g766 ( .A(n_559), .B(n_767), .Y(n_766) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g579 ( .A(n_560), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_565), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g610 ( .A(n_565), .B(n_579), .Y(n_610) );
INVx2_ASAP7_75t_L g627 ( .A(n_565), .Y(n_627) );
AND2x4_ASAP7_75t_L g644 ( .A(n_565), .B(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_565), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_571), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g756 ( .A(n_575), .B(n_578), .Y(n_756) );
AND2x4_ASAP7_75t_L g602 ( .A(n_576), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g643 ( .A(n_576), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g670 ( .A(n_576), .B(n_610), .Y(n_670) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
AND2x2_ASAP7_75t_L g774 ( .A(n_578), .B(n_775), .Y(n_774) );
BUFx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g626 ( .A(n_579), .B(n_627), .Y(n_626) );
OAI21xp5_ASAP7_75t_SL g646 ( .A1(n_580), .A2(n_647), .B(n_653), .Y(n_646) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_593), .Y(n_583) );
INVx1_ASAP7_75t_SL g700 ( .A(n_584), .Y(n_700) );
AND2x2_ASAP7_75t_L g730 ( .A(n_584), .B(n_640), .Y(n_730) );
AND2x4_ASAP7_75t_L g741 ( .A(n_584), .B(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g607 ( .A(n_585), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g614 ( .A(n_585), .Y(n_614) );
AND2x4_ASAP7_75t_L g620 ( .A(n_585), .B(n_606), .Y(n_620) );
INVx2_ASAP7_75t_L g631 ( .A(n_585), .Y(n_631) );
INVx1_ASAP7_75t_L g680 ( .A(n_585), .Y(n_680) );
OR2x2_ASAP7_75t_L g701 ( .A(n_585), .B(n_685), .Y(n_701) );
OR2x2_ASAP7_75t_L g715 ( .A(n_585), .B(n_595), .Y(n_715) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_585), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_585), .B(n_637), .Y(n_787) );
OR2x6_ASAP7_75t_L g585 ( .A(n_586), .B(n_592), .Y(n_585) );
INVx1_ASAP7_75t_L g632 ( .A(n_593), .Y(n_632) );
AND2x2_ASAP7_75t_L g765 ( .A(n_593), .B(n_631), .Y(n_765) );
AND2x2_ASAP7_75t_L g790 ( .A(n_593), .B(n_620), .Y(n_790) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g608 ( .A(n_595), .Y(n_608) );
BUFx3_ASAP7_75t_L g650 ( .A(n_595), .Y(n_650) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_595), .Y(n_677) );
INVx1_ASAP7_75t_L g686 ( .A(n_595), .Y(n_686) );
AOI33xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_604), .A3(n_609), .B1(n_610), .B2(n_611), .B3(n_612), .Y(n_601) );
AOI21x1_ASAP7_75t_SL g704 ( .A1(n_602), .A2(n_626), .B(n_688), .Y(n_704) );
INVx2_ASAP7_75t_L g734 ( .A(n_602), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_602), .B(n_733), .Y(n_740) );
AND2x2_ASAP7_75t_L g688 ( .A(n_603), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
AND2x2_ASAP7_75t_L g651 ( .A(n_606), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g752 ( .A(n_607), .Y(n_752) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_608), .Y(n_742) );
OAI32xp33_ASAP7_75t_L g791 ( .A1(n_609), .A2(n_611), .A3(n_787), .B1(n_792), .B2(n_794), .Y(n_791) );
AND2x2_ASAP7_75t_L g709 ( .A(n_610), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g699 ( .A(n_611), .Y(n_699) );
AND2x2_ASAP7_75t_L g764 ( .A(n_611), .B(n_708), .Y(n_764) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_625), .B1(n_628), .B2(n_642), .C(n_646), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_619), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_620), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_620), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_620), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g669 ( .A(n_624), .Y(n_669) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_633), .C(n_638), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_630), .A2(n_692), .B1(n_732), .B2(n_735), .Y(n_731) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g635 ( .A(n_631), .Y(n_635) );
NOR2x1p5_ASAP7_75t_L g649 ( .A(n_631), .B(n_650), .Y(n_649) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_631), .Y(n_671) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI322xp33_ASAP7_75t_L g698 ( .A1(n_634), .A2(n_676), .A3(n_699), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_704), .Y(n_698) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_636), .A2(n_655), .B(n_656), .C(n_658), .Y(n_654) );
OR2x2_ASAP7_75t_L g746 ( .A(n_636), .B(n_700), .Y(n_746) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g653 ( .A(n_637), .B(n_641), .Y(n_653) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g659 ( .A(n_643), .B(n_660), .Y(n_659) );
INVx3_ASAP7_75t_SL g691 ( .A(n_644), .Y(n_691) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_648), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_SL g695 ( .A(n_651), .Y(n_695) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_652), .Y(n_737) );
OR2x6_ASAP7_75t_SL g792 ( .A(n_655), .B(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI211xp5_ASAP7_75t_L g782 ( .A1(n_660), .A2(n_783), .B(n_784), .C(n_791), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_664), .B(n_667), .C(n_671), .Y(n_661) );
OAI211xp5_ASAP7_75t_SL g673 ( .A1(n_662), .A2(n_674), .B(n_681), .C(n_705), .Y(n_673) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_718), .C(n_762), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_678), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_677), .Y(n_769) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g724 ( .A(n_680), .Y(n_724) );
NOR3xp33_ASAP7_75t_SL g681 ( .A(n_682), .B(n_694), .C(n_698), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_687), .B1(n_690), .B2(n_693), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g726 ( .A(n_686), .Y(n_726) );
INVxp67_ASAP7_75t_SL g793 ( .A(n_686), .Y(n_793) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_SL g779 ( .A(n_692), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
OR2x2_ASAP7_75t_L g729 ( .A(n_695), .B(n_715), .Y(n_729) );
OR2x2_ASAP7_75t_L g780 ( .A(n_695), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g778 ( .A(n_703), .Y(n_778) );
OR2x2_ASAP7_75t_L g794 ( .A(n_703), .B(n_733), .Y(n_794) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B(n_711), .Y(n_705) );
OAI31xp33_ASAP7_75t_L g719 ( .A1(n_706), .A2(n_720), .A3(n_721), .B(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g751 ( .A(n_716), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND4xp25_ASAP7_75t_SL g718 ( .A(n_719), .B(n_727), .C(n_738), .D(n_743), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_726), .Y(n_761) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_747), .B1(n_751), .B2(n_753), .C(n_755), .Y(n_743) );
NAND2xp33_ASAP7_75t_SL g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g788 ( .A(n_747), .Y(n_788) );
AND2x2_ASAP7_75t_SL g747 ( .A(n_748), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AOI21xp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B(n_759), .Y(n_755) );
INVx1_ASAP7_75t_L g783 ( .A(n_757), .Y(n_783) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_763), .B(n_782), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_766), .B2(n_768), .C(n_772), .Y(n_763) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVx1_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
AOI21xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_777), .B(n_780), .Y(n_772) );
INVxp33_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_796), .Y(n_800) );
CKINVDCx11_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
OAI21xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_804), .B(n_825), .Y(n_801) );
INVx2_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_808), .B(n_820), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_805), .A2(n_821), .B(n_822), .Y(n_820) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g821 ( .A(n_809), .Y(n_821) );
XNOR2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_814), .Y(n_809) );
NAND3x1_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .C(n_813), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g819 ( .A(n_817), .Y(n_819) );
CKINVDCx11_ASAP7_75t_R g827 ( .A(n_822), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_823), .Y(n_822) );
BUFx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
endmodule