module real_jpeg_31335_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_0),
.Y(n_242)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_0),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_1),
.Y(n_115)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_3),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_4),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_4),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_4),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_4),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_4),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_4),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_5),
.B(n_63),
.Y(n_62)
);

NAND2x1p5_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_5),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_5),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_5),
.B(n_49),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_5),
.B(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_6),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_6),
.Y(n_132)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_7),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_7),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_7),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_7),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_7),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_7),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_8),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_8),
.B(n_95),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_10),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_49),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_10),
.B(n_74),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_12),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_13),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_13),
.B(n_68),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g142 ( 
.A(n_13),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_13),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_13),
.B(n_31),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_14),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_14),
.B(n_180),
.Y(n_179)
);

BUFx24_ASAP7_75t_L g208 ( 
.A(n_14),
.Y(n_208)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_14),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_15),
.B(n_44),
.Y(n_43)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_15),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_15),
.B(n_49),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_15),
.B(n_25),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_15),
.B(n_44),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_189),
.Y(n_16)
);

NAND2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_188),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_161),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_20),
.B(n_161),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_107),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_65),
.C(n_92),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_22),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.C(n_50),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_23),
.B(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_24),
.B(n_29),
.C(n_34),
.Y(n_125)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_27),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_34),
.B2(n_40),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_33),
.Y(n_251)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_38),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_41),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_198)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_43),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_43),
.B(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_43),
.A2(n_46),
.B1(n_157),
.B2(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_46),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_49),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_61),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_52),
.A2(n_61),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_52),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_55),
.Y(n_287)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_56),
.B(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_60),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_61),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_64),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_65),
.B(n_93),
.Y(n_163)
);

XOR2x1_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_76),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_66)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_70),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_75),
.C(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_73),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.C(n_87),
.Y(n_77)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_81),
.Y(n_214)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_83),
.A2(n_87),
.B1(n_88),
.B2(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_105),
.B2(n_106),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_94),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_97),
.C(n_101),
.Y(n_159)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_136),
.B2(n_160),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_126),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.C(n_125),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_118),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_116),
.C(n_118),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_118),
.B(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_119),
.A2(n_120),
.B1(n_125),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_120),
.A2(n_121),
.B(n_124),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_131),
.Y(n_134)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_132),
.Y(n_210)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_148),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_147),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_146),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_158),
.B2(n_159),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

AO22x1_ASAP7_75t_SL g295 ( 
.A1(n_151),
.A2(n_152),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_151),
.B(n_296),
.Y(n_309)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_183),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_184),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.C(n_171),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_170),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.C(n_179),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_173),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_174),
.B(n_179),
.Y(n_327)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_222),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_195),
.A2(n_199),
.B1(n_200),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_195),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_197),
.B(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.C(n_219),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_201),
.B(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_205),
.A2(n_219),
.B1(n_220),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_205),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.C(n_215),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_206),
.A2(n_207),
.B1(n_215),
.B2(n_216),
.Y(n_305)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_208),
.B(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_208),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_208),
.B(n_286),
.Y(n_285)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_211),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp33_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2x1p5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AOI21x1_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_330),
.B(n_335),
.Y(n_225)
);

OAI21x1_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_319),
.B(n_329),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_299),
.B(n_318),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_277),
.B(n_298),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_260),
.B(n_276),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_231),
.B(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_232),
.A2(n_233),
.B1(n_239),
.B2(n_240),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_232),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx4f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_253),
.C(n_255),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_248),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_246),
.B(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_269),
.B(n_275),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_268),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_268),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_279),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_291),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_292),
.C(n_295),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_288),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_285),
.C(n_288),
.Y(n_307)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_296),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_301),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_308),
.B1(n_316),
.B2(n_317),
.Y(n_301)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_307),
.C(n_316),
.Y(n_328)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_311),
.C(n_314),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_328),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_328),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_325),
.C(n_326),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_334),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_334),
.Y(n_335)
);


endmodule