module fake_jpeg_24454_n_233 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_29),
.B(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_15),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_33),
.B1(n_29),
.B2(n_31),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_46),
.B1(n_51),
.B2(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_25),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_50),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_17),
.B1(n_27),
.B2(n_22),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_21),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_53),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_31),
.A2(n_26),
.B1(n_16),
.B2(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_25),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_54),
.B(n_25),
.C(n_34),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_0),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_62),
.B(n_54),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_52),
.B1(n_29),
.B2(n_46),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_44),
.B1(n_23),
.B2(n_49),
.Y(n_92)
);

MAJx3_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_38),
.C(n_30),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_66),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_17),
.B1(n_22),
.B2(n_48),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_54),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_54),
.B1(n_51),
.B2(n_43),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_92),
.B1(n_100),
.B2(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_48),
.B1(n_44),
.B2(n_40),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_69),
.B1(n_75),
.B2(n_55),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_55),
.B1(n_49),
.B2(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_58),
.B(n_73),
.C(n_38),
.D(n_68),
.Y(n_104)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_94),
.Y(n_101)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_93),
.A2(n_49),
.B1(n_55),
.B2(n_41),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_47),
.B(n_24),
.C(n_20),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_23),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_64),
.C(n_70),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_71),
.B1(n_76),
.B2(n_58),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_91),
.B1(n_85),
.B2(n_80),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_79),
.C(n_92),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_114),
.B1(n_96),
.B2(n_82),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_110),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_60),
.B(n_44),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_25),
.B1(n_21),
.B2(n_20),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_97),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_24),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_77),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_19),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_106),
.B(n_111),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_81),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_124),
.B1(n_133),
.B2(n_134),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_91),
.B1(n_85),
.B2(n_113),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_141),
.B(n_104),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_112),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_137),
.C(n_103),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_96),
.B1(n_82),
.B2(n_88),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_94),
.B1(n_30),
.B2(n_34),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_117),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_38),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_34),
.B1(n_30),
.B2(n_60),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_138),
.A2(n_110),
.B1(n_116),
.B2(n_107),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_142),
.A2(n_106),
.B(n_19),
.Y(n_144)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_155),
.C(n_161),
.Y(n_166)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_101),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_101),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_152),
.B(n_156),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_141),
.B(n_123),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_0),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_19),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_157),
.A2(n_144),
.B1(n_127),
.B2(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_133),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_13),
.C(n_5),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_146),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_137),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_168),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_154),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_129),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_132),
.C(n_136),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_177),
.C(n_166),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_142),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_186),
.C(n_188),
.Y(n_194)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_182),
.B(n_184),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_143),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_157),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

AO221x1_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_163),
.B1(n_166),
.B2(n_161),
.C(n_170),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_172),
.A2(n_159),
.B1(n_151),
.B2(n_149),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_181),
.A2(n_174),
.B1(n_175),
.B2(n_169),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_198),
.B1(n_186),
.B2(n_180),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_194),
.Y(n_207)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_200),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_169),
.B(n_154),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_185),
.B(n_149),
.Y(n_202)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_196),
.C(n_8),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_205),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_6),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_148),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_201),
.A2(n_180),
.B1(n_171),
.B2(n_128),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_208),
.C(n_209),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_201),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_2),
.B(n_5),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_6),
.C(n_7),
.Y(n_209)
);

FAx1_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_200),
.CI(n_197),
.CON(n_211),
.SN(n_211)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_215),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_209),
.B1(n_203),
.B2(n_12),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_6),
.C(n_8),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_9),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_219),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_207),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_9),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_212),
.C(n_216),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_225),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_222),
.A2(n_211),
.B(n_214),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_222),
.B(n_12),
.Y(n_227)
);

OAI311xp33_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_224),
.A3(n_13),
.B1(n_11),
.C1(n_228),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_229),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_11),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_11),
.B(n_13),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_232),
.Y(n_233)
);


endmodule