module fake_jpeg_9100_n_285 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_285);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_6),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_18),
.B1(n_25),
.B2(n_27),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_23),
.B1(n_18),
.B2(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_51),
.Y(n_62)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_23),
.B1(n_18),
.B2(n_37),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_59),
.B1(n_61),
.B2(n_65),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_23),
.B1(n_18),
.B2(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_60),
.B(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_23),
.B1(n_29),
.B2(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_54),
.B1(n_39),
.B2(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_50),
.B1(n_21),
.B2(n_20),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_24),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_93),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_84),
.Y(n_102)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_54),
.B1(n_49),
.B2(n_26),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_94),
.B1(n_97),
.B2(n_21),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_49),
.C(n_30),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_26),
.B1(n_48),
.B2(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_60),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_73),
.B1(n_70),
.B2(n_72),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_61),
.B1(n_65),
.B2(n_63),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_108),
.B1(n_85),
.B2(n_80),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_73),
.B1(n_69),
.B2(n_63),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_106),
.B(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_103),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_111),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_71),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_68),
.B1(n_59),
.B2(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_13),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

AO22x1_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_14),
.B1(n_19),
.B2(n_15),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_0),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_30),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_15),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_13),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_88),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_119),
.B(n_88),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_120),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_131),
.B1(n_84),
.B2(n_78),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_134),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_143),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_107),
.B1(n_108),
.B2(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_77),
.B(n_27),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_139),
.B(n_27),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_77),
.B(n_22),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_148),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_147),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_142),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_116),
.C(n_106),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_155),
.C(n_168),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_152),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_157),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_106),
.C(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_166),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_163),
.B(n_167),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_128),
.B1(n_34),
.B2(n_32),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_120),
.A2(n_115),
.B(n_83),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_121),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_115),
.C(n_91),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_127),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_177),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_131),
.B1(n_138),
.B2(n_126),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_170),
.A2(n_173),
.B1(n_176),
.B2(n_186),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_171),
.B(n_163),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_138),
.B1(n_134),
.B2(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_122),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_174),
.B(n_183),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_124),
.B1(n_128),
.B2(n_92),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_155),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_161),
.A2(n_19),
.B1(n_14),
.B2(n_15),
.Y(n_182)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_146),
.A2(n_19),
.B1(n_15),
.B2(n_31),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_147),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_176),
.B1(n_181),
.B2(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_166),
.B(n_144),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_209),
.B(n_1),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_146),
.C(n_168),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_200),
.C(n_208),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_148),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_191),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_144),
.C(n_153),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_205),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_159),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_160),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_172),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_173),
.A2(n_158),
.B1(n_167),
.B2(n_19),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_182),
.B1(n_186),
.B2(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

NAND2x1_ASAP7_75t_SL g213 ( 
.A(n_195),
.B(n_189),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_220),
.B(n_192),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_191),
.C(n_169),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_223),
.C(n_227),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_189),
.B(n_10),
.Y(n_218)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_22),
.Y(n_219)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_198),
.B(n_203),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_224),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_34),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_34),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_32),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_196),
.C(n_32),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_206),
.B1(n_192),
.B2(n_204),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_239),
.B1(n_218),
.B2(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_16),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_196),
.C(n_31),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_241),
.C(n_215),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_7),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_246),
.C(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_238),
.C(n_211),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_252),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_223),
.C(n_228),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_226),
.B1(n_8),
.B2(n_11),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_254),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_22),
.C(n_3),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_232),
.B(n_242),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_16),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_236),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_7),
.B1(n_12),
.B2(n_6),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_243),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_234),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_264),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_265),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_263),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_240),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_251),
.B(n_233),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_237),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_257),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_241),
.B(n_16),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_271),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_256),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_2),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_266),
.C(n_270),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_273),
.B(n_5),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_4),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_277),
.C(n_5),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_4),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_R g283 ( 
.A(n_282),
.B(n_22),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_22),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_16),
.B1(n_79),
.B2(n_276),
.Y(n_285)
);


endmodule