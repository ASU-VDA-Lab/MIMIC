module fake_ariane_1129_n_168 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_168);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_168;

wire n_83;
wire n_56;
wire n_60;
wire n_160;
wire n_64;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_152;
wire n_120;
wire n_106;
wire n_53;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_144;
wire n_130;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_43;
wire n_87;
wire n_81;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_54;

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_2),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_3),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_5),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_7),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_8),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_9),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_11),
.C(n_13),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_15),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_53),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_17),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_68),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_62),
.B(n_63),
.C(n_54),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_75),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_54),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_59),
.B(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_67),
.B(n_19),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_18),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_72),
.B(n_89),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_96),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

AO21x2_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_83),
.B(n_81),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_85),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_86),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_84),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_84),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_90),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_100),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_86),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

AOI21x1_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_114),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_20),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

AOI21x1_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_117),
.B(n_114),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_114),
.B(n_116),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_116),
.B1(n_113),
.B2(n_107),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_113),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_119),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_116),
.C(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_108),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_108),
.B1(n_112),
.B2(n_30),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_123),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_124),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_129),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_140),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_143),
.C(n_141),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_130),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_155),
.Y(n_161)
);

OAI221xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_156),
.B1(n_142),
.B2(n_134),
.C(n_151),
.Y(n_162)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_156),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_161),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_163),
.B1(n_162),
.B2(n_127),
.C(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

OAI221xp5_ASAP7_75t_R g168 ( 
.A1(n_167),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.C(n_36),
.Y(n_168)
);


endmodule