module fake_aes_10943_n_31 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_31);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g10 ( .A(n_3), .B(n_8), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
INVxp67_ASAP7_75t_SL g17 ( .A(n_10), .Y(n_17) );
AOI221xp5_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_0), .B1(n_3), .B2(n_4), .C(n_5), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_13), .B(n_0), .Y(n_19) );
BUFx3_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AOI22x1_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_15), .B1(n_13), .B2(n_10), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_16), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI311xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_18), .A3(n_16), .B(n_12), .C(n_21), .Y(n_25) );
NOR2xp33_ASAP7_75t_L g26 ( .A(n_24), .B(n_18), .Y(n_26) );
NOR3xp33_ASAP7_75t_SL g27 ( .A(n_26), .B(n_15), .C(n_7), .Y(n_27) );
NOR3x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_6), .C(n_9), .Y(n_28) );
NAND2xp33_ASAP7_75t_SL g29 ( .A(n_28), .B(n_27), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
XNOR2xp5_ASAP7_75t_L g31 ( .A(n_30), .B(n_28), .Y(n_31) );
endmodule