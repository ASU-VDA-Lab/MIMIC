module fake_jpeg_1945_n_518 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_518);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_518;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_14),
.B(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_52),
.Y(n_140)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g133 ( 
.A(n_54),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_55),
.B(n_69),
.Y(n_129)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_58),
.Y(n_128)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_60),
.Y(n_162)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_68),
.B(n_71),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_45),
.Y(n_70)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_1),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_45),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_82),
.B(n_97),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_36),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_15),
.B(n_13),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_1),
.Y(n_113)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_36),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_1),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g155 ( 
.A(n_94),
.B(n_28),
.CON(n_155),
.SN(n_155)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_23),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_38),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_102),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_38),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_25),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_104),
.B(n_25),
.Y(n_110)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

BUFx16f_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_110),
.B(n_78),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_44),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_70),
.A2(n_24),
.B1(n_46),
.B2(n_41),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_117),
.A2(n_136),
.B1(n_103),
.B2(n_43),
.Y(n_175)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_124),
.B(n_150),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_51),
.A2(n_49),
.B1(n_48),
.B2(n_47),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_68),
.A2(n_26),
.B(n_32),
.Y(n_145)
);

OR2x2_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_155),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_71),
.A2(n_24),
.B1(n_26),
.B2(n_32),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_43),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_58),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_63),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_94),
.B(n_41),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_69),
.B(n_46),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_159),
.B(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_101),
.B(n_44),
.Y(n_163)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_173),
.B(n_174),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g237 ( 
.A1(n_175),
.A2(n_117),
.B1(n_157),
.B2(n_135),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_176),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_133),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_177),
.B(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_205),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_129),
.A2(n_82),
.B1(n_108),
.B2(n_152),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_185),
.A2(n_214),
.B1(n_112),
.B2(n_162),
.Y(n_228)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_187),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_116),
.B(n_39),
.Y(n_188)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_114),
.Y(n_189)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_190),
.Y(n_252)
);

CKINVDCx12_ASAP7_75t_R g192 ( 
.A(n_133),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_192),
.Y(n_247)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_39),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_211),
.Y(n_218)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_199),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_133),
.B(n_33),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_137),
.A2(n_33),
.B(n_49),
.C(n_48),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_212),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_111),
.B(n_30),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_203),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_132),
.B(n_30),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_204),
.Y(n_219)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_155),
.B(n_47),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_210),
.Y(n_243)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_105),
.B(n_19),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_109),
.B(n_85),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_215),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_127),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_162),
.B1(n_131),
.B2(n_128),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_220),
.A2(n_230),
.B1(n_212),
.B2(n_141),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_146),
.B1(n_131),
.B2(n_128),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_115),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_121),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_168),
.B(n_123),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_200),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_153),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_250),
.B(n_142),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_251),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_253),
.B(n_265),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_179),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_266),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_256),
.B(n_267),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_184),
.B1(n_180),
.B2(n_154),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_260),
.B1(n_226),
.B2(n_252),
.Y(n_289)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_258),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_168),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_259),
.A2(n_264),
.B(n_239),
.Y(n_302)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_261),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_218),
.A2(n_212),
.B1(n_167),
.B2(n_120),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_262),
.A2(n_273),
.B1(n_276),
.B2(n_239),
.Y(n_301)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_214),
.B(n_157),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_245),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_182),
.Y(n_266)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_183),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_277),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_218),
.A2(n_140),
.B1(n_164),
.B2(n_143),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_271),
.A2(n_274),
.B1(n_230),
.B2(n_219),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_186),
.B(n_189),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_229),
.B(n_244),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_216),
.B1(n_243),
.B2(n_233),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_240),
.A2(n_164),
.B1(n_65),
.B2(n_81),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_232),
.Y(n_275)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_240),
.A2(n_197),
.B1(n_171),
.B2(n_169),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_190),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_241),
.Y(n_278)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_226),
.B(n_215),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_205),
.Y(n_312)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_285),
.Y(n_315)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_266),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_263),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_237),
.B1(n_225),
.B2(n_252),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_291),
.A2(n_268),
.B1(n_160),
.B2(n_135),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_223),
.C(n_237),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_293),
.C(n_294),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_237),
.C(n_221),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_267),
.C(n_272),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_295),
.A2(n_302),
.B(n_304),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_273),
.A2(n_236),
.B1(n_181),
.B2(n_170),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_297),
.A2(n_260),
.B1(n_280),
.B2(n_258),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_229),
.C(n_246),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_298),
.B(n_301),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_256),
.A2(n_244),
.B(n_232),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_227),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_274),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_264),
.A2(n_222),
.B(n_227),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_276),
.B(n_282),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_312),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_262),
.B(n_242),
.C(n_127),
.Y(n_313)
);

A2O1A1O1Ixp25_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_253),
.B(n_254),
.C(n_279),
.D(n_278),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_270),
.B(n_265),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_269),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_303),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_322),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_320),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_303),
.Y(n_321)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_321),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_271),
.Y(n_324)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_269),
.Y(n_325)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_328),
.Y(n_371)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_308),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_312),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_331),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_330),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_283),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_258),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_335),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_333),
.A2(n_339),
.B1(n_305),
.B2(n_288),
.Y(n_376)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_275),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_337),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_275),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_291),
.A2(n_268),
.B1(n_224),
.B2(n_248),
.Y(n_339)
);

OA21x2_ASAP7_75t_L g340 ( 
.A1(n_302),
.A2(n_242),
.B(n_261),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_340),
.A2(n_342),
.B1(n_304),
.B2(n_301),
.Y(n_351)
);

INVx13_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_341),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_284),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_344),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_284),
.B(n_217),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_217),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_345),
.B(n_300),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_338),
.A2(n_309),
.B(n_292),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_348),
.A2(n_353),
.B(n_356),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_294),
.C(n_293),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_364),
.C(n_327),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_351),
.A2(n_372),
.B1(n_376),
.B2(n_333),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_315),
.A2(n_285),
.B1(n_296),
.B2(n_307),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_352),
.A2(n_329),
.B1(n_330),
.B2(n_324),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_338),
.A2(n_316),
.B(n_341),
.Y(n_353)
);

NAND2x1_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_299),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_307),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_360),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_319),
.A2(n_343),
.B(n_317),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_359),
.A2(n_320),
.B(n_326),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_306),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_325),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_366),
.Y(n_387)
);

XOR2x2_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_297),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_367),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_313),
.C(n_311),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_322),
.B(n_331),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_365),
.B(n_305),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_336),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_315),
.B(n_313),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_332),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_321),
.A2(n_311),
.B1(n_288),
.B2(n_287),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_377),
.A2(n_393),
.B1(n_394),
.B2(n_399),
.Y(n_412)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g382 ( 
.A(n_358),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_382),
.B(n_391),
.Y(n_406)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_375),
.Y(n_383)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_384),
.A2(n_371),
.B(n_373),
.Y(n_415)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_385),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_392),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_388),
.A2(n_355),
.B1(n_373),
.B2(n_368),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_390),
.Y(n_418)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_340),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_352),
.A2(n_340),
.B1(n_339),
.B2(n_330),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_361),
.A2(n_342),
.B1(n_323),
.B2(n_344),
.Y(n_394)
);

A2O1A1O1Ixp25_ASAP7_75t_L g395 ( 
.A1(n_361),
.A2(n_340),
.B(n_323),
.C(n_335),
.D(n_328),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_395),
.A2(n_401),
.B(n_403),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_345),
.C(n_287),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_398),
.C(n_402),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_400),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_300),
.C(n_261),
.Y(n_398)
);

NAND3xp33_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_300),
.C(n_186),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_353),
.A2(n_204),
.B(n_195),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_348),
.B(n_367),
.C(n_347),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_359),
.A2(n_15),
.B(n_16),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_176),
.C(n_210),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_380),
.C(n_392),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_381),
.A2(n_356),
.B(n_357),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_403),
.B(n_389),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_393),
.A2(n_355),
.B1(n_351),
.B2(n_370),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_413),
.A2(n_397),
.B1(n_385),
.B2(n_172),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_414),
.A2(n_416),
.B1(n_425),
.B2(n_421),
.Y(n_447)
);

XOR2x2_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_158),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_387),
.A2(n_346),
.B1(n_374),
.B2(n_363),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_389),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_377),
.A2(n_374),
.B1(n_372),
.B2(n_365),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_420),
.A2(n_424),
.B1(n_427),
.B2(n_191),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_356),
.Y(n_422)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_422),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_73),
.C(n_86),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_404),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_394),
.A2(n_19),
.B1(n_16),
.B2(n_141),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_384),
.A2(n_154),
.B1(n_76),
.B2(n_52),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_381),
.A2(n_191),
.B1(n_80),
.B2(n_67),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_415),
.Y(n_428)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_422),
.Y(n_430)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_396),
.C(n_380),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_433),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_441),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_398),
.C(n_402),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_434),
.B(n_435),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_436),
.A2(n_442),
.B1(n_445),
.B2(n_122),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_414),
.A2(n_194),
.B1(n_158),
.B2(n_114),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_437),
.A2(n_447),
.B1(n_427),
.B2(n_425),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_209),
.C(n_114),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_443),
.Y(n_463)
);

XNOR2x1_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_107),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_444),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_412),
.A2(n_158),
.B1(n_90),
.B2(n_72),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_413),
.A2(n_417),
.B1(n_407),
.B2(n_421),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_418),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_411),
.A2(n_417),
.B(n_410),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_2),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_446),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_405),
.B(n_209),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_448),
.B(n_408),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_429),
.Y(n_450)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_450),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_423),
.C(n_416),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_451),
.B(n_454),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_452),
.B(n_444),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_453),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_405),
.C(n_407),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_434),
.B(n_426),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_455),
.B(n_457),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_428),
.B(n_426),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_408),
.C(n_209),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_458),
.B(n_437),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_SL g471 ( 
.A(n_464),
.B(n_439),
.Y(n_471)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_442),
.B1(n_430),
.B2(n_436),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_468),
.B(n_469),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_454),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_471),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_456),
.A2(n_441),
.B1(n_448),
.B2(n_209),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_472),
.B(n_473),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_28),
.C(n_22),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_22),
.C(n_3),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_474),
.B(n_476),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_22),
.C(n_4),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_465),
.B(n_2),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_478),
.B(n_461),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_4),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_479),
.B(n_481),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_4),
.Y(n_481)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_484),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_462),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_488),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_463),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_452),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_493),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_480),
.B(n_459),
.Y(n_493)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_482),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_489),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_470),
.A2(n_460),
.B(n_459),
.Y(n_495)
);

MAJx2_ASAP7_75t_L g504 ( 
.A(n_495),
.B(n_6),
.C(n_10),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_490),
.A2(n_460),
.B(n_474),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_496),
.A2(n_503),
.B(n_11),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_473),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_497),
.A2(n_499),
.B(n_501),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_6),
.Y(n_506)
);

NAND3xp33_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_476),
.C(n_479),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_502),
.A2(n_487),
.B(n_491),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_SL g503 ( 
.A1(n_486),
.A2(n_481),
.B1(n_7),
.B2(n_8),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_504),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_505),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_506),
.B(n_507),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_509),
.A2(n_498),
.B(n_502),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_511),
.A2(n_508),
.B(n_11),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_513),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_510),
.B(n_11),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_514),
.B(n_512),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_12),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_517),
.A2(n_12),
.B(n_505),
.Y(n_518)
);


endmodule