module fake_jpeg_22355_n_255 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_1),
.Y(n_71)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_21),
.B1(n_16),
.B2(n_18),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_61),
.B1(n_21),
.B2(n_22),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_33),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_20),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_28),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_78),
.Y(n_88)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_73),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_77),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_15),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_61),
.B1(n_30),
.B2(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_15),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_50),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_97),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_55),
.B1(n_63),
.B2(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_93),
.B1(n_80),
.B2(n_65),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_55),
.B1(n_43),
.B2(n_63),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_35),
.B(n_34),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_65),
.B(n_24),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_102),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_101),
.Y(n_129)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_80),
.B1(n_79),
.B2(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_58),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_35),
.B1(n_28),
.B2(n_20),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_109),
.Y(n_125)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_107),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_75),
.C(n_32),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_94),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_130),
.B(n_114),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_93),
.Y(n_132)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_126),
.B1(n_131),
.B2(n_108),
.Y(n_147)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_86),
.B1(n_72),
.B2(n_69),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_38),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_104),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_86),
.B1(n_102),
.B2(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_70),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_148),
.B1(n_150),
.B2(n_23),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_146),
.C(n_115),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_103),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_139),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_138),
.B(n_31),
.Y(n_168)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_104),
.A3(n_91),
.B1(n_103),
.B2(n_87),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_140),
.A2(n_145),
.B(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_122),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_154),
.B1(n_153),
.B2(n_140),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_130),
.B(n_131),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_151),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_89),
.B1(n_100),
.B2(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_100),
.B1(n_52),
.B2(n_68),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_88),
.B(n_100),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_88),
.B1(n_113),
.B2(n_123),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_155),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_161),
.C(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_26),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_48),
.C(n_47),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_31),
.C(n_26),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_145),
.B1(n_149),
.B2(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_170),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_31),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_171),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_169),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_31),
.C(n_19),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_22),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_172),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_31),
.C(n_2),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_146),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_154),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_187),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_185),
.A2(n_161),
.B(n_162),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_158),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_149),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_188)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_193),
.B(n_134),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_192),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_159),
.B1(n_173),
.B2(n_171),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_156),
.C(n_163),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_191),
.C(n_189),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_204),
.B(n_205),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_5),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_184),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_220),
.C(n_201),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_212),
.B(n_211),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_182),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_179),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_217),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_199),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_178),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_223),
.C(n_224),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_196),
.C(n_198),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_199),
.C(n_203),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_195),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_225),
.B(n_230),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_227),
.Y(n_233)
);

OAI221xp5_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_200),
.B1(n_183),
.B2(n_179),
.C(n_213),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_229),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_207),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_206),
.B(n_8),
.Y(n_230)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_231),
.Y(n_241)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_216),
.B(n_220),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_235),
.A2(n_11),
.B(n_12),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_10),
.Y(n_243)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_7),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_9),
.B(n_10),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_233),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_240),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_231),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_242),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_243),
.A2(n_238),
.B(n_14),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_244),
.A2(n_232),
.B(n_11),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_246),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_245),
.B(n_248),
.Y(n_251)
);

INVxp33_ASAP7_75t_SL g252 ( 
.A(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_252),
.B(n_250),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_243),
.C(n_11),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_14),
.B(n_246),
.Y(n_255)
);


endmodule