module fake_jpeg_562_n_525 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_59),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_21),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_90),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_15),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_64),
.A2(n_66),
.B(n_72),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_71),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_21),
.B(n_13),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_75),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_76),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_23),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_89),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_78),
.Y(n_199)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_82),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_83),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_27),
.Y(n_84)
);

HAxp5_ASAP7_75t_SL g193 ( 
.A(n_84),
.B(n_87),
.CON(n_193),
.SN(n_193)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_14),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_85),
.B(n_105),
.Y(n_189)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_27),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_14),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_20),
.B(n_41),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_93),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_98),
.Y(n_173)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_29),
.B(n_14),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_107),
.Y(n_141)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_104),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_20),
.B(n_1),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_24),
.B(n_1),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

BUFx24_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_24),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_110),
.B(n_2),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_31),
.B(n_2),
.C(n_4),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_52),
.Y(n_132)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_22),
.Y(n_113)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_30),
.Y(n_114)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_22),
.Y(n_116)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_48),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_37),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_22),
.Y(n_121)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_66),
.B1(n_120),
.B2(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_129),
.A2(n_135),
.B1(n_137),
.B2(n_142),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_84),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_131),
.B(n_153),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_132),
.A2(n_177),
.B(n_7),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_37),
.B1(n_50),
.B2(n_55),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_136),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_52),
.B1(n_55),
.B2(n_35),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_72),
.B(n_33),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_139),
.B(n_130),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_52),
.B1(n_35),
.B2(n_50),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_85),
.A2(n_31),
.B1(n_55),
.B2(n_35),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_145),
.A2(n_151),
.B1(n_168),
.B2(n_192),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_109),
.A2(n_37),
.B1(n_50),
.B2(n_53),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_87),
.B(n_54),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_57),
.B(n_54),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_160),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_60),
.B(n_51),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_61),
.B(n_51),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_165),
.B(n_171),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_121),
.A2(n_42),
.B1(n_40),
.B2(n_53),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_169),
.A2(n_193),
.B1(n_182),
.B2(n_138),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_62),
.A2(n_45),
.B1(n_39),
.B2(n_33),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_170),
.A2(n_135),
.B1(n_151),
.B2(n_164),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_65),
.B(n_39),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_78),
.A2(n_32),
.B1(n_30),
.B2(n_18),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_157),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_71),
.B(n_32),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_188),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_76),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_82),
.B(n_2),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_196),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_83),
.A2(n_18),
.B1(n_49),
.B2(n_7),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_108),
.B(n_5),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_136),
.B(n_106),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_203),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_137),
.A2(n_97),
.B1(n_94),
.B2(n_91),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_204),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_129),
.A2(n_49),
.B(n_80),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_123),
.B(n_98),
.C(n_18),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_206),
.B(n_262),
.C(n_265),
.Y(n_271)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_142),
.A2(n_49),
.B(n_18),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_209),
.Y(n_300)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_210),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_124),
.B(n_5),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_211),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_164),
.B(n_6),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_212),
.B(n_205),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_213),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_122),
.B(n_6),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_214),
.B(n_218),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_148),
.A2(n_49),
.B1(n_7),
.B2(n_8),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_216),
.Y(n_310)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_6),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_228),
.Y(n_276)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_223),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_49),
.B1(n_10),
.B2(n_11),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_224),
.A2(n_249),
.B1(n_255),
.B2(n_257),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_225),
.B(n_234),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_226),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_230),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_139),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_240),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_127),
.Y(n_233)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_233),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_125),
.B(n_166),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_237),
.A2(n_252),
.B1(n_144),
.B2(n_180),
.Y(n_273)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_141),
.B(n_189),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_241),
.B(n_248),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_172),
.B(n_183),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_253),
.Y(n_284)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_147),
.Y(n_244)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_244),
.Y(n_301)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_127),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_251),
.Y(n_287)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_246),
.B(n_260),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_247),
.B(n_250),
.Y(n_305)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_152),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_163),
.A2(n_185),
.B1(n_183),
.B2(n_126),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_128),
.B(n_146),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_170),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_150),
.A2(n_175),
.B1(n_179),
.B2(n_174),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_149),
.B(n_174),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_154),
.Y(n_254)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_149),
.A2(n_179),
.B1(n_158),
.B2(n_199),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_199),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_256),
.B(n_266),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_155),
.A2(n_176),
.B1(n_156),
.B2(n_184),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_201),
.B(n_158),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_259),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_201),
.B(n_186),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_154),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_181),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_263),
.Y(n_293)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_128),
.B(n_156),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_134),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_134),
.B(n_180),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_252),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_128),
.B(n_140),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_140),
.B(n_184),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_268),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_140),
.B(n_184),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_214),
.B(n_143),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_269),
.B(n_291),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_273),
.A2(n_303),
.B1(n_308),
.B2(n_315),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_251),
.A2(n_144),
.B1(n_186),
.B2(n_176),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_285),
.A2(n_294),
.B1(n_309),
.B2(n_311),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_SL g291 ( 
.A(n_231),
.B(n_218),
.C(n_239),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_243),
.A2(n_156),
.B1(n_176),
.B2(n_209),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_L g349 ( 
.A(n_296),
.B(n_315),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_207),
.A2(n_221),
.B1(n_237),
.B2(n_238),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_202),
.B(n_247),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_304),
.B(n_270),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_210),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_240),
.B(n_238),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_230),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_242),
.A2(n_206),
.B1(n_258),
.B2(n_253),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_235),
.A2(n_225),
.B1(n_264),
.B2(n_259),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_236),
.A2(n_203),
.B1(n_215),
.B2(n_211),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_203),
.A2(n_211),
.B1(n_234),
.B2(n_266),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_256),
.A2(n_220),
.B1(n_223),
.B2(n_244),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_263),
.B1(n_217),
.B2(n_222),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_L g320 ( 
.A1(n_270),
.A2(n_234),
.B(n_265),
.C(n_262),
.D(n_208),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_320),
.A2(n_337),
.B(n_340),
.Y(n_378)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_324),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_325),
.B(n_329),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_295),
.Y(n_327)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_327),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_228),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_328),
.B(n_334),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_262),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_265),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g367 ( 
.A1(n_330),
.A2(n_314),
.B(n_293),
.Y(n_367)
);

OR2x4_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_299),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_SL g374 ( 
.A1(n_331),
.A2(n_347),
.B(n_282),
.C(n_318),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_346),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_289),
.Y(n_333)
);

CKINVDCx11_ASAP7_75t_R g387 ( 
.A(n_333),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_229),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_303),
.A2(n_284),
.B1(n_292),
.B2(n_300),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_335),
.A2(n_339),
.B1(n_355),
.B2(n_358),
.Y(n_364)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_290),
.Y(n_336)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_299),
.A2(n_261),
.B(n_213),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_317),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_292),
.A2(n_246),
.B1(n_233),
.B2(n_245),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_278),
.A2(n_260),
.B1(n_254),
.B2(n_248),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_286),
.B(n_227),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_353),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_300),
.A2(n_298),
.B(n_276),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_342),
.A2(n_349),
.B(n_274),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_302),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_343),
.B(n_350),
.Y(n_384)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_313),
.Y(n_346)
);

O2A1O1Ixp33_ASAP7_75t_SL g347 ( 
.A1(n_287),
.A2(n_292),
.B(n_298),
.C(n_294),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_313),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_SL g375 ( 
.A(n_348),
.B(n_295),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_307),
.B(n_269),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_351),
.B(n_352),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_308),
.B(n_309),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_356),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_286),
.A2(n_273),
.B1(n_306),
.B2(n_278),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_288),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_281),
.B(n_317),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_297),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_314),
.A2(n_272),
.B1(n_312),
.B2(n_271),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_321),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_341),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_373),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_337),
.A2(n_314),
.B(n_310),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_375),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_370),
.B(n_381),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_345),
.A2(n_271),
.B1(n_310),
.B2(n_285),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_372),
.A2(n_326),
.B1(n_322),
.B2(n_357),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_319),
.Y(n_373)
);

A2O1A1O1Ixp25_ASAP7_75t_L g398 ( 
.A1(n_374),
.A2(n_330),
.B(n_342),
.C(n_347),
.D(n_329),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_344),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_354),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_331),
.A2(n_297),
.B(n_318),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_379),
.B(n_382),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_335),
.A2(n_277),
.B1(n_318),
.B2(n_301),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_383),
.A2(n_353),
.B1(n_325),
.B2(n_336),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_326),
.A2(n_301),
.B1(n_280),
.B2(n_274),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_385),
.A2(n_363),
.B1(n_389),
.B2(n_366),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_275),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_390),
.Y(n_396)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_347),
.B(n_280),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_391),
.B(n_402),
.Y(n_440)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_395),
.Y(n_434)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_397),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_398),
.Y(n_442)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_389),
.Y(n_399)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_322),
.C(n_338),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_410),
.C(n_382),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_362),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_360),
.B(n_348),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_403),
.B(n_409),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_362),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_405),
.Y(n_424)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_386),
.Y(n_406)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_406),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_377),
.Y(n_408)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_330),
.C(n_324),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_411),
.Y(n_430)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_387),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_364),
.A2(n_355),
.B1(n_339),
.B2(n_323),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_413),
.A2(n_383),
.B1(n_369),
.B2(n_385),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_414),
.B(n_364),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_360),
.B(n_346),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_415),
.B(n_417),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_361),
.B(n_333),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_416),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_384),
.B(n_283),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_420),
.Y(n_448)
);

NOR4xp25_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_379),
.C(n_359),
.D(n_374),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_419),
.A2(n_374),
.B1(n_392),
.B2(n_390),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_407),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_429),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_359),
.C(n_372),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_416),
.C(n_400),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_365),
.Y(n_429)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_374),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_378),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_435),
.A2(n_413),
.B1(n_400),
.B2(n_412),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_380),
.Y(n_436)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_436),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_283),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_411),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_443),
.A2(n_421),
.B1(n_439),
.B2(n_424),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_449),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_402),
.C(n_405),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_456),
.C(n_460),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_422),
.A2(n_396),
.B1(n_391),
.B2(n_408),
.Y(n_447)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_393),
.Y(n_449)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_450),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_440),
.A2(n_393),
.B(n_398),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_451),
.A2(n_452),
.B(n_419),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_441),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_453),
.B(n_439),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_459),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_374),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_461),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_387),
.C(n_406),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_432),
.A2(n_399),
.B1(n_394),
.B2(n_397),
.Y(n_457)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_457),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_433),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_378),
.C(n_395),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_435),
.A2(n_388),
.B1(n_371),
.B2(n_376),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_432),
.A2(n_371),
.B1(n_320),
.B2(n_332),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_463),
.B(n_458),
.Y(n_470)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_470),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_446),
.A2(n_424),
.B(n_440),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_471),
.A2(n_459),
.B(n_445),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_472),
.B(n_474),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_421),
.C(n_425),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_425),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_476),
.B(n_479),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_430),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_477),
.B(n_438),
.Y(n_486)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_478),
.A2(n_465),
.B(n_474),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_430),
.Y(n_479)
);

A2O1A1Ixp33_ASAP7_75t_SL g480 ( 
.A1(n_478),
.A2(n_451),
.B(n_461),
.C(n_460),
.Y(n_480)
);

AOI22x1_ASAP7_75t_L g494 ( 
.A1(n_480),
.A2(n_475),
.B1(n_454),
.B2(n_455),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g481 ( 
.A(n_464),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_483),
.Y(n_498)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_472),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_486),
.B(n_487),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_445),
.C(n_448),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_468),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_438),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_491),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_469),
.C(n_473),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_499),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_494),
.Y(n_508)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_496),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_473),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_466),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_482),
.A2(n_475),
.B1(n_476),
.B2(n_479),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_489),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_SL g505 ( 
.A(n_500),
.B(n_480),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_484),
.A2(n_423),
.B1(n_428),
.B2(n_434),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_501),
.B(n_423),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_505),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_428),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_507),
.Y(n_514)
);

FAx1_ASAP7_75t_SL g507 ( 
.A(n_493),
.B(n_480),
.CI(n_449),
.CON(n_507),
.SN(n_507)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_509),
.B(n_466),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_493),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_510),
.Y(n_512)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_511),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_498),
.Y(n_515)
);

AOI21xp33_ASAP7_75t_L g520 ( 
.A1(n_515),
.A2(n_434),
.B(n_371),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_494),
.C(n_496),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_516),
.A2(n_504),
.B(n_508),
.Y(n_519)
);

AO21x1_ASAP7_75t_SL g518 ( 
.A1(n_513),
.A2(n_507),
.B(n_508),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_519),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_520),
.A2(n_514),
.B(n_512),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_517),
.C(n_516),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_522),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_375),
.Y(n_525)
);


endmodule