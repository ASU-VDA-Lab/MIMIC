module fake_jpeg_564_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_43;
wire n_37;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_17),
.A2(n_18),
.B1(n_25),
.B2(n_22),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_14),
.B1(n_13),
.B2(n_10),
.Y(n_18)
);

CKINVDCx12_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_27),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_14),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_24)
);

OA21x2_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_17),
.B(n_26),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_13),
.A2(n_3),
.B1(n_9),
.B2(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_15),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_32),
.B(n_36),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_34),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_33),
.B1(n_32),
.B2(n_36),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_15),
.B(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_41),
.Y(n_43)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AO221x1_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_39),
.B1(n_38),
.B2(n_33),
.C(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_45),
.B(n_37),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_37),
.B(n_29),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_46),
.Y(n_49)
);


endmodule