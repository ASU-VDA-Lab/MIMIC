module fake_jpeg_22328_n_133 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_33),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_40),
.B1(n_25),
.B2(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_22),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_56),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_20),
.B(n_28),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_13),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_1),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_63),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_42),
.B1(n_23),
.B2(n_29),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_68),
.B1(n_73),
.B2(n_79),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_23),
.B1(n_21),
.B2(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_5),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_21),
.B1(n_5),
.B2(n_8),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_48),
.B1(n_43),
.B2(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_12),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_13),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_60),
.B1(n_61),
.B2(n_52),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_60),
.B1(n_49),
.B2(n_59),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_89),
.B1(n_91),
.B2(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_52),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_94),
.C(n_64),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_76),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_99),
.Y(n_109)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_98),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_83),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_80),
.C(n_78),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_80),
.B1(n_64),
.B2(n_77),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_85),
.B1(n_90),
.B2(n_86),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_107),
.C(n_101),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_66),
.B1(n_68),
.B2(n_82),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_99),
.B1(n_106),
.B2(n_104),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_82),
.B1(n_86),
.B2(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_109),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_114),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_112),
.B(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_124),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g129 ( 
.A(n_125),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_108),
.C(n_118),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_125),
.B(n_88),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

OAI31xp33_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_120),
.A3(n_85),
.B(n_126),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_129),
.B(n_93),
.Y(n_133)
);


endmodule