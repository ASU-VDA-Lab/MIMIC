module real_jpeg_25560_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_4),
.A2(n_39),
.B1(n_51),
.B2(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_4),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_4),
.A2(n_55),
.B1(n_56),
.B2(n_84),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_4),
.A2(n_26),
.B1(n_30),
.B2(n_84),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_26),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_6),
.B(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_6),
.B(n_56),
.C(n_58),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_39),
.B1(n_43),
.B2(n_51),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_6),
.B(n_82),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_6),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_6),
.B(n_26),
.C(n_90),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_6),
.A2(n_25),
.B(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_7),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_9),
.A2(n_26),
.B1(n_30),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_74),
.Y(n_87)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_11),
.A2(n_39),
.B1(n_51),
.B2(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_62),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_11),
.A2(n_26),
.B1(n_30),
.B2(n_62),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_13),
.A2(n_39),
.B1(n_51),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_13),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_65),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_65),
.B1(n_98),
.B2(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_13),
.A2(n_26),
.B1(n_30),
.B2(n_65),
.Y(n_123)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_14),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_126),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_104),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_18),
.B(n_104),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_77),
.B2(n_78),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_52),
.B1(n_75),
.B2(n_76),
.Y(n_20)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_36),
.B2(n_37),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_24),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_163)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_25),
.A2(n_29),
.B1(n_33),
.B2(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_25),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_26),
.A2(n_30),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_27),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_30),
.B(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_33),
.A2(n_165),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B(n_42),
.C(n_46),
.Y(n_37)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_39),
.B1(n_47),
.B2(n_51),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_38),
.A2(n_44),
.B1(n_47),
.B2(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_39),
.B(n_117),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_42),
.A2(n_43),
.B(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_43),
.B(n_88),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_43),
.B(n_178),
.Y(n_177)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_48),
.C(n_51),
.Y(n_46)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_69),
.C(n_72),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_60),
.B(n_63),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_56),
.B1(n_89),
.B2(n_90),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_56),
.B(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_66),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_64),
.B(n_82),
.Y(n_136)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_67),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_95),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B(n_91),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_88),
.A2(n_91),
.B(n_132),
.Y(n_148)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_112),
.B1(n_114),
.B2(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B(n_101),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_115),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_106),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_115),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B(n_113),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_110),
.A2(n_113),
.B(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_118),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_122),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_140),
.B(n_190),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_137),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_128),
.B(n_137),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.C(n_133),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_184),
.B(n_189),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_161),
.B(n_183),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_155),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_155),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_148),
.C(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_159),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_170),
.B(n_182),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_168),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_175),
.B(n_181),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_173),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_188),
.Y(n_189)
);


endmodule