module fake_netlist_6_2516_n_1906 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1906);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1906;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_72),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_135),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_183),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_90),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_102),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_45),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_53),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_3),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_14),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_15),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_137),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_19),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_23),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_41),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_120),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_40),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_153),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_136),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_177),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_57),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_11),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_154),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_58),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_81),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_94),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_116),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_53),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_82),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_39),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_93),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_147),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_0),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_71),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_79),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_43),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_152),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_70),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_155),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_144),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_176),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_25),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_184),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_68),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_57),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_130),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_67),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_104),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_97),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_62),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_178),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_54),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_141),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_9),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_107),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_126),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_1),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_33),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_142),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_31),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_55),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_108),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_100),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_54),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_12),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_115),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_132),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_25),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_98),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_60),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_163),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_44),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_148),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_145),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_111),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_16),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_37),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_95),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_73),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_59),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_170),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_45),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_138),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_166),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_55),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_143),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_88),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_36),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_118),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_117),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_175),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_114),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_63),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_22),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_14),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_23),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_87),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_48),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_113),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_15),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_164),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_8),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_80),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_179),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_26),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_134),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_38),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_106),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_123),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_31),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_162),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_1),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_34),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_36),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_182),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_51),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_8),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_29),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_172),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_39),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_41),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_35),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_156),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_110),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_10),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_74),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_150),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_26),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_186),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_10),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_17),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_12),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_83),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_13),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_50),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_58),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_128),
.Y(n_338)
);

INVx4_ASAP7_75t_R g339 ( 
.A(n_181),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_35),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_78),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_50),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_49),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_140),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_151),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_52),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_149),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_99),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_171),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_92),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_103),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_42),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_185),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_34),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_69),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_125),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_44),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_65),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_91),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_66),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_16),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_3),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_49),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_101),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_167),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_89),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_121),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_64),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_112),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_29),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_75),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_51),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_86),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_11),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_19),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_13),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_32),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_76),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_180),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_40),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_129),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_77),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_33),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_30),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_281),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_250),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_228),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_234),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_286),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_286),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_229),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_245),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_251),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_281),
.Y(n_394)
);

INVxp33_ASAP7_75t_SL g395 ( 
.A(n_196),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_281),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_281),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_281),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_204),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_212),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_276),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_267),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_206),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_253),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_212),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_259),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_283),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_283),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_289),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_267),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_235),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_236),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_289),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_199),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_255),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_261),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_262),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_241),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_196),
.Y(n_419)
);

BUFx2_ASAP7_75t_SL g420 ( 
.A(n_246),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_329),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_258),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_266),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_271),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_269),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_273),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_296),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_277),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_278),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_295),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_299),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_259),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_308),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_297),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_301),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_317),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_326),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_331),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_254),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_238),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_240),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_243),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_333),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_303),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_313),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_259),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_244),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_315),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_306),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_248),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_197),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_197),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_254),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_300),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_300),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_306),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_332),
.Y(n_462)
);

BUFx2_ASAP7_75t_SL g463 ( 
.A(n_246),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_318),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_358),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_358),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_194),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_205),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_207),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_210),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_220),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_257),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_222),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_224),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_227),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_260),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_282),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_343),
.Y(n_478)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_201),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_343),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_346),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_230),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_346),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_357),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_232),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_419),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_385),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_387),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_477),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_477),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_414),
.A2(n_337),
.B1(n_336),
.B2(n_370),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_382),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_385),
.B(n_382),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_477),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_391),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_200),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_477),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_402),
.A2(n_242),
.B(n_200),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_411),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_453),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_459),
.B(n_242),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_458),
.B(n_467),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_468),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_460),
.B(n_292),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_394),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_396),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_412),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_397),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_398),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_458),
.B(n_189),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_410),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_441),
.Y(n_516)
);

OA21x2_ASAP7_75t_L g517 ( 
.A1(n_410),
.A2(n_363),
.B(n_357),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_408),
.A2(n_413),
.B(n_409),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_408),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_413),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_478),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_478),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g524 ( 
.A(n_458),
.B(n_282),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_393),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_469),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_480),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_480),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_481),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_442),
.Y(n_530)
);

BUFx8_ASAP7_75t_L g531 ( 
.A(n_465),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_470),
.B(n_292),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_481),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_483),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_483),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_457),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_484),
.Y(n_537)
);

NOR2x1_ASAP7_75t_L g538 ( 
.A(n_420),
.B(n_345),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_484),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_466),
.B(n_345),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_388),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_471),
.B(n_473),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_475),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_388),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_485),
.B(n_189),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_399),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_403),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_389),
.A2(n_237),
.B(n_233),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_418),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_422),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_425),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_427),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_400),
.B(n_363),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_431),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_433),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_390),
.A2(n_247),
.B(n_239),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_440),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_437),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_438),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_439),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_444),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_440),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_447),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_454),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_455),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_563),
.B(n_386),
.Y(n_567)
);

AND3x2_ASAP7_75t_L g568 ( 
.A(n_541),
.B(n_314),
.C(n_448),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_563),
.B(n_420),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_515),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_487),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_497),
.B(n_282),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_513),
.B(n_401),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_487),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_557),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_492),
.B(n_463),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_546),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_495),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_495),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_495),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_546),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_517),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_492),
.B(n_463),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_541),
.B(n_456),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_497),
.B(n_282),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_547),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_501),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_517),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_513),
.B(n_395),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_497),
.B(n_282),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_557),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_492),
.B(n_405),
.Y(n_596)
);

NOR2x1p5_ASAP7_75t_L g597 ( 
.A(n_509),
.B(n_392),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_517),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_517),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_550),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_515),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_550),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_519),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_552),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_495),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_519),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_519),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_557),
.B(n_392),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_557),
.B(n_395),
.Y(n_609)
);

INVx8_ASAP7_75t_L g610 ( 
.A(n_524),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_552),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_538),
.B(n_347),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_557),
.B(n_404),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_554),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_L g615 ( 
.A(n_545),
.B(n_415),
.C(n_404),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_519),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_554),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_486),
.B(n_421),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_520),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_488),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_555),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_555),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

BUFx8_ASAP7_75t_SL g624 ( 
.A(n_488),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_520),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_559),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_553),
.B(n_432),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_559),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_520),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_524),
.B(n_347),
.Y(n_630)
);

AND3x1_ASAP7_75t_L g631 ( 
.A(n_491),
.B(n_479),
.C(n_252),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_495),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_SL g633 ( 
.A1(n_541),
.A2(n_451),
.B1(n_406),
.B2(n_461),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_520),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_521),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_560),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_560),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_SL g638 ( 
.A(n_486),
.B(n_201),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_521),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_521),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_561),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_553),
.B(n_347),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_564),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_524),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_521),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_564),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_516),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_553),
.B(n_416),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_502),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_558),
.B(n_347),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_522),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_524),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_505),
.B(n_416),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_505),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_L g655 ( 
.A1(n_491),
.A2(n_265),
.B1(n_198),
.B2(n_311),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_515),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_502),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_522),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_536),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_495),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_505),
.B(n_417),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_544),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_515),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_505),
.B(n_417),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_526),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_526),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_545),
.B(n_424),
.C(n_423),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_536),
.B(n_424),
.C(n_423),
.Y(n_668)
);

BUFx4f_ASAP7_75t_L g669 ( 
.A(n_544),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_558),
.B(n_347),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_526),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_526),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_515),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_543),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_494),
.B(n_426),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_544),
.B(n_462),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_496),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_543),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_522),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_494),
.B(n_426),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_522),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_558),
.B(n_371),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_530),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_523),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_496),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_523),
.Y(n_686)
);

BUFx4f_ASAP7_75t_L g687 ( 
.A(n_558),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_515),
.Y(n_688)
);

BUFx10_ASAP7_75t_L g689 ( 
.A(n_532),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_523),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_525),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_504),
.B(n_479),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_543),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_543),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_523),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_494),
.B(n_428),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_504),
.B(n_443),
.Y(n_697)
);

INVx8_ASAP7_75t_L g698 ( 
.A(n_524),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_558),
.B(n_371),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_494),
.Y(n_700)
);

AND2x6_ASAP7_75t_L g701 ( 
.A(n_494),
.B(n_371),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_543),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_527),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_542),
.A2(n_231),
.B1(n_209),
.B2(n_322),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_558),
.B(n_371),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_527),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_527),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_503),
.B(n_429),
.Y(n_708)
);

AND2x6_ASAP7_75t_L g709 ( 
.A(n_503),
.B(n_249),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_507),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_558),
.B(n_429),
.Y(n_711)
);

NOR3xp33_ASAP7_75t_L g712 ( 
.A(n_668),
.B(n_434),
.C(n_430),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_571),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_577),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_692),
.B(n_449),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_571),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_593),
.B(n_576),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_574),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_582),
.B(n_589),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_700),
.B(n_531),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_647),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_700),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_627),
.B(n_430),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_574),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_708),
.B(n_452),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_697),
.A2(n_476),
.B1(n_472),
.B2(n_506),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_586),
.B(n_506),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_578),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_578),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_596),
.B(n_506),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_689),
.B(n_531),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_648),
.B(n_649),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_600),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_618),
.B(n_434),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_573),
.B(n_531),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_675),
.A2(n_540),
.B1(n_310),
.B2(n_445),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_583),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_709),
.B(n_267),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_654),
.B(n_540),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_665),
.B(n_540),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_666),
.B(n_515),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_602),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_671),
.B(n_515),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_672),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_615),
.B(n_435),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_583),
.B(n_566),
.Y(n_746)
);

NOR2x1p5_ASAP7_75t_L g747 ( 
.A(n_676),
.B(n_445),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_604),
.B(n_562),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_611),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_689),
.B(n_531),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_595),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_585),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_585),
.B(n_565),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_614),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_592),
.B(n_565),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_592),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_657),
.B(n_659),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_598),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_617),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_689),
.B(n_531),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_621),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_598),
.A2(n_500),
.B1(n_518),
.B2(n_556),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_599),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_599),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_622),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_657),
.B(n_446),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_667),
.B(n_446),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_680),
.A2(n_211),
.B1(n_192),
.B2(n_312),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_595),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_609),
.B(n_566),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_626),
.B(n_566),
.Y(n_771)
);

NOR2x1p5_ASAP7_75t_L g772 ( 
.A(n_696),
.B(n_450),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_628),
.B(n_566),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_636),
.B(n_566),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_637),
.B(n_566),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_653),
.B(n_450),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_603),
.Y(n_777)
);

OR2x2_ASAP7_75t_L g778 ( 
.A(n_659),
.B(n_464),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_647),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_606),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_606),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_674),
.A2(n_500),
.B(n_548),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_641),
.B(n_565),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_643),
.B(n_565),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_646),
.B(n_565),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_L g786 ( 
.A(n_567),
.B(n_464),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_678),
.B(n_267),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_572),
.B(n_565),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_662),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_L g790 ( 
.A(n_709),
.B(n_267),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_572),
.B(n_565),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_661),
.B(n_325),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_607),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_710),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_588),
.B(n_499),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_623),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_693),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_709),
.B(n_267),
.Y(n_798)
);

OAI22xp33_ASAP7_75t_L g799 ( 
.A1(n_587),
.A2(n_542),
.B1(n_327),
.B2(n_328),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_669),
.B(n_587),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_711),
.A2(n_532),
.B1(n_264),
.B2(n_263),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_677),
.B(n_203),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_587),
.A2(n_288),
.B1(n_256),
.B2(n_268),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_588),
.B(n_642),
.Y(n_804)
);

AND2x6_ASAP7_75t_L g805 ( 
.A(n_694),
.B(n_274),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_702),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_607),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_669),
.B(n_562),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_616),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_616),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_619),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_642),
.B(n_499),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_579),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_619),
.Y(n_814)
);

O2A1O1Ixp5_ASAP7_75t_L g815 ( 
.A1(n_711),
.A2(n_670),
.B(n_682),
.C(n_650),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_594),
.B(n_499),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_591),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_587),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_625),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_683),
.B(n_562),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_R g821 ( 
.A(n_683),
.B(n_525),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_709),
.A2(n_500),
.B1(n_518),
.B2(n_556),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_664),
.B(n_267),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_624),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_644),
.B(n_267),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_579),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_594),
.B(n_608),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_594),
.B(n_499),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_594),
.B(n_499),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_610),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_625),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_569),
.B(n_512),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_613),
.B(n_190),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_709),
.B(n_270),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_594),
.B(n_532),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_594),
.B(n_532),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_673),
.B(n_532),
.Y(n_837)
);

NAND2xp33_ASAP7_75t_L g838 ( 
.A(n_709),
.B(n_272),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_673),
.B(n_688),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_673),
.B(n_518),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_638),
.B(n_321),
.C(n_319),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_688),
.B(n_518),
.Y(n_842)
);

BUFx6f_ASAP7_75t_SL g843 ( 
.A(n_591),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_688),
.B(n_518),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_575),
.B(n_518),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_707),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_633),
.B(n_190),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_575),
.B(n_508),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_612),
.A2(n_556),
.B1(n_548),
.B2(n_524),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_624),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_644),
.B(n_279),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_663),
.B(n_508),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_629),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_663),
.B(n_510),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_663),
.B(n_510),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_569),
.B(n_191),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_629),
.A2(n_548),
.B(n_287),
.C(n_369),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_569),
.A2(n_285),
.B1(n_275),
.B2(n_280),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_644),
.B(n_291),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_707),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_704),
.B(n_191),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_655),
.B(n_193),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_579),
.B(n_580),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_706),
.Y(n_864)
);

BUFx8_ASAP7_75t_L g865 ( 
.A(n_685),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_631),
.A2(n_349),
.B1(n_294),
.B2(n_293),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_638),
.B(n_193),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_644),
.B(n_195),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_634),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_634),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_568),
.B(n_195),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_713),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_717),
.B(n_792),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_746),
.A2(n_687),
.B(n_601),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_713),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_792),
.B(n_591),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_728),
.B(n_729),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_728),
.B(n_706),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_729),
.B(n_635),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_737),
.B(n_752),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_737),
.B(n_635),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_752),
.A2(n_216),
.B1(n_215),
.B2(n_203),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_732),
.B(n_644),
.Y(n_883)
);

NOR2x2_ASAP7_75t_L g884 ( 
.A(n_862),
.B(n_620),
.Y(n_884)
);

OR2x2_ASAP7_75t_SL g885 ( 
.A(n_841),
.B(n_734),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_821),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_757),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_716),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_776),
.B(n_808),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_716),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_718),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_776),
.A2(n_597),
.B1(n_612),
.B2(n_701),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_861),
.A2(n_612),
.B1(n_701),
.B2(n_341),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_718),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_756),
.B(n_639),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_724),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_724),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_SL g898 ( 
.A1(n_715),
.A2(n_620),
.B1(n_691),
.B2(n_375),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_830),
.B(n_652),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_789),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_748),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_722),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_756),
.B(n_639),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_766),
.B(n_723),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_777),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_748),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_714),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_758),
.B(n_640),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_758),
.B(n_640),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_725),
.A2(n_612),
.B1(n_701),
.B2(n_656),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_763),
.A2(n_383),
.B1(n_215),
.B2(n_216),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_715),
.B(n_570),
.Y(n_912)
);

AND2x6_ASAP7_75t_SL g913 ( 
.A(n_862),
.B(n_307),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_820),
.B(n_652),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_865),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_865),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_733),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_721),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_763),
.B(n_645),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_722),
.Y(n_920)
);

AND2x6_ASAP7_75t_SL g921 ( 
.A(n_861),
.B(n_309),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_778),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_821),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_742),
.Y(n_924)
);

NOR2x1p5_ASAP7_75t_L g925 ( 
.A(n_817),
.B(n_218),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_764),
.B(n_727),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_722),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_SL g928 ( 
.A1(n_779),
.A2(n_354),
.B1(n_361),
.B2(n_226),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_867),
.A2(n_612),
.B1(n_701),
.B2(n_320),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_725),
.A2(n_767),
.B1(n_745),
.B2(n_832),
.Y(n_930)
);

NOR3xp33_ASAP7_75t_SL g931 ( 
.A(n_866),
.B(n_223),
.C(n_218),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_726),
.B(n_549),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_722),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_751),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_749),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_761),
.B(n_512),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_780),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_786),
.B(n_549),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_751),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_802),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_764),
.B(n_730),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_754),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_840),
.B(n_645),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_751),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_772),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_800),
.B(n_761),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_842),
.B(n_651),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_759),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_751),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_867),
.A2(n_612),
.B1(n_701),
.B2(n_350),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_765),
.B(n_719),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_844),
.B(n_651),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_745),
.A2(n_701),
.B1(n_656),
.B2(n_601),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_767),
.A2(n_656),
.B1(n_570),
.B2(n_601),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_744),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_739),
.B(n_658),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_781),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_740),
.B(n_797),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_856),
.B(n_799),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_817),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_824),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_794),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_850),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_806),
.B(n_658),
.Y(n_964)
);

INVx6_ASAP7_75t_L g965 ( 
.A(n_747),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_744),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_719),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_793),
.Y(n_968)
);

INVx5_ASAP7_75t_L g969 ( 
.A(n_830),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_804),
.A2(n_359),
.B1(n_364),
.B2(n_368),
.Y(n_970)
);

INVx8_ASAP7_75t_L g971 ( 
.A(n_843),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_769),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_856),
.B(n_202),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_770),
.B(n_679),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_765),
.B(n_652),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_793),
.Y(n_976)
);

INVx3_ASAP7_75t_SL g977 ( 
.A(n_847),
.Y(n_977)
);

AND2x6_ASAP7_75t_L g978 ( 
.A(n_830),
.B(n_827),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_818),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_830),
.B(n_858),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_736),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_796),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_813),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_796),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_753),
.B(n_679),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_871),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_755),
.B(n_681),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_807),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_807),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_796),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_768),
.B(n_652),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_810),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_796),
.B(n_514),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_810),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_871),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_803),
.B(n_202),
.Y(n_996)
);

INVx5_ASAP7_75t_L g997 ( 
.A(n_805),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_831),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_848),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_845),
.A2(n_687),
.B(n_610),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_831),
.B(n_846),
.Y(n_1001)
);

OR2x6_ASAP7_75t_L g1002 ( 
.A(n_720),
.B(n_610),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_846),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_813),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_SL g1005 ( 
.A(n_833),
.B(n_226),
.C(n_223),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_SL g1006 ( 
.A1(n_857),
.A2(n_705),
.B(n_682),
.C(n_699),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_712),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_860),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_769),
.B(n_580),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_801),
.B(n_208),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_860),
.B(n_681),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_869),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_735),
.A2(n_356),
.B1(n_367),
.B2(n_581),
.Y(n_1013)
);

INVxp67_ASAP7_75t_SL g1014 ( 
.A(n_826),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_823),
.B(n_514),
.Y(n_1015)
);

NOR3xp33_ASAP7_75t_SL g1016 ( 
.A(n_823),
.B(n_361),
.C(n_375),
.Y(n_1016)
);

CKINVDCx11_ASAP7_75t_R g1017 ( 
.A(n_843),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_869),
.B(n_684),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_809),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_731),
.B(n_213),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_826),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_762),
.A2(n_383),
.B1(n_377),
.B2(n_374),
.Y(n_1022)
);

BUFx5_ASAP7_75t_L g1023 ( 
.A(n_811),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_814),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_771),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_819),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_870),
.B(n_684),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_853),
.B(n_686),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_805),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_731),
.B(n_213),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_864),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_762),
.B(n_837),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_805),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_863),
.B(n_214),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_750),
.B(n_214),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_805),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_795),
.B(n_533),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_805),
.A2(n_610),
.B1(n_698),
.B2(n_690),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_773),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_750),
.B(n_217),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_787),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_852),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_839),
.Y(n_1043)
);

NOR2x2_ASAP7_75t_L g1044 ( 
.A(n_760),
.B(n_549),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_854),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_760),
.B(n_217),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_774),
.B(n_219),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_835),
.B(n_219),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_787),
.B(n_533),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_934),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_959),
.A2(n_834),
.B1(n_838),
.B2(n_836),
.Y(n_1051)
);

BUFx8_ASAP7_75t_SL g1052 ( 
.A(n_886),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_904),
.B(n_534),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_874),
.A2(n_782),
.B(n_743),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_963),
.B(n_738),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_941),
.A2(n_687),
.B(n_698),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_941),
.A2(n_698),
.B(n_822),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_873),
.B(n_812),
.Y(n_1058)
);

AND2x6_ASAP7_75t_L g1059 ( 
.A(n_980),
.B(n_788),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_900),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_SL g1061 ( 
.A(n_969),
.B(n_221),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_918),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_971),
.B(n_698),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_907),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_926),
.A2(n_822),
.B(n_849),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_926),
.A2(n_849),
.B(n_791),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_985),
.A2(n_741),
.B(n_815),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_930),
.B(n_775),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_912),
.B(n_855),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_889),
.B(n_999),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_934),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_969),
.A2(n_798),
.B(n_790),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_973),
.A2(n_868),
.B1(n_783),
.B2(n_784),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_960),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_905),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_971),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_981),
.B(n_785),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1041),
.A2(n_958),
.B(n_932),
.C(n_924),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_958),
.B(n_581),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_R g1080 ( 
.A(n_923),
.B(n_816),
.Y(n_1080)
);

NOR2x1_ASAP7_75t_SL g1081 ( 
.A(n_969),
.B(n_851),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_946),
.A2(n_829),
.B1(n_828),
.B2(n_859),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_SL g1083 ( 
.A(n_1036),
.B(n_221),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_1017),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_971),
.B(n_851),
.Y(n_1085)
);

AOI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1022),
.A2(n_362),
.B1(n_372),
.B2(n_374),
.C(n_377),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_969),
.A2(n_660),
.B(n_632),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_955),
.B(n_225),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_940),
.B(n_534),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_987),
.A2(n_605),
.B(n_825),
.Y(n_1090)
);

OR2x6_ASAP7_75t_SL g1091 ( 
.A(n_1022),
.B(n_335),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_922),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_934),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1042),
.B(n_605),
.Y(n_1094)
);

OAI21xp33_ASAP7_75t_L g1095 ( 
.A1(n_887),
.A2(n_340),
.B(n_352),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_939),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_917),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_902),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_877),
.A2(n_880),
.B1(n_1032),
.B2(n_893),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_955),
.B(n_225),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_935),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_R g1102 ( 
.A(n_1016),
.B(n_284),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_877),
.A2(n_859),
.B1(n_551),
.B2(n_549),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1010),
.A2(n_551),
.B1(n_353),
.B2(n_355),
.Y(n_1104)
);

CKINVDCx16_ASAP7_75t_R g1105 ( 
.A(n_898),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_SL g1106 ( 
.A1(n_1007),
.A2(n_373),
.B1(n_366),
.B2(n_365),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_SL g1107 ( 
.A1(n_977),
.A2(n_373),
.B1(n_366),
.B2(n_365),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_986),
.B(n_284),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_942),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_979),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_995),
.Y(n_1111)
);

NOR3xp33_ASAP7_75t_L g1112 ( 
.A(n_876),
.B(n_379),
.C(n_353),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_948),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_951),
.B(n_355),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_902),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_880),
.A2(n_551),
.B1(n_379),
.B2(n_378),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_974),
.A2(n_660),
.B(n_590),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_936),
.B(n_967),
.Y(n_1118)
);

NOR2xp67_ASAP7_75t_SL g1119 ( 
.A(n_997),
.B(n_360),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_SL g1120 ( 
.A1(n_936),
.A2(n_381),
.B1(n_378),
.B2(n_360),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_974),
.A2(n_584),
.B(n_590),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_962),
.A2(n_825),
.B(n_699),
.C(n_605),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_937),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_872),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_966),
.B(n_381),
.Y(n_1125)
);

NOR2x1_ASAP7_75t_L g1126 ( 
.A(n_927),
.B(n_511),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1045),
.B(n_686),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_R g1128 ( 
.A(n_961),
.B(n_290),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_965),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_885),
.B(n_298),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_902),
.B(n_302),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_920),
.Y(n_1132)
);

BUFx8_ASAP7_75t_L g1133 ( 
.A(n_915),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_956),
.B(n_1025),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1039),
.B(n_938),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_R g1136 ( 
.A(n_927),
.B(n_304),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_901),
.B(n_539),
.Y(n_1137)
);

OAI22x1_ASAP7_75t_L g1138 ( 
.A1(n_925),
.A2(n_305),
.B1(n_316),
.B2(n_324),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1032),
.A2(n_539),
.B1(n_695),
.B2(n_690),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_943),
.A2(n_584),
.B(n_590),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1034),
.B(n_695),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_996),
.A2(n_703),
.B(n_630),
.C(n_529),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_929),
.A2(n_703),
.B1(n_660),
.B2(n_632),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_875),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_945),
.B(n_528),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_943),
.A2(n_660),
.B(n_632),
.Y(n_1146)
);

INVx6_ASAP7_75t_L g1147 ( 
.A(n_965),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_906),
.B(n_528),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_939),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_993),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_888),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_950),
.A2(n_632),
.B1(n_590),
.B2(n_584),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_890),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1043),
.B(n_528),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_920),
.B(n_330),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_920),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_933),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_933),
.B(n_529),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_933),
.Y(n_1159)
);

AOI22x1_ASAP7_75t_L g1160 ( 
.A1(n_1015),
.A2(n_334),
.B1(n_338),
.B2(n_344),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_928),
.B(n_348),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_891),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_947),
.A2(n_952),
.B(n_1000),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1044),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_957),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_952),
.A2(n_524),
.B(n_493),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1043),
.B(n_1049),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_931),
.B(n_351),
.Y(n_1168)
);

BUFx5_ASAP7_75t_L g1169 ( 
.A(n_978),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_882),
.B(n_911),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1036),
.B(n_339),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_894),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_987),
.A2(n_498),
.B(n_489),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_882),
.B(n_0),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1043),
.B(n_537),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_896),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1009),
.A2(n_498),
.B(n_489),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_989),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_897),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_916),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_968),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_994),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_911),
.B(n_2),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_921),
.B(n_2),
.Y(n_1184)
);

OAI22x1_ASAP7_75t_L g1185 ( 
.A1(n_913),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_1185)
);

OR2x6_ASAP7_75t_SL g1186 ( 
.A(n_884),
.B(n_4),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_892),
.A2(n_498),
.B(n_489),
.C(n_493),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_972),
.A2(n_493),
.B(n_490),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_SL g1189 ( 
.A(n_997),
.B(n_524),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_878),
.A2(n_490),
.B(n_535),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1049),
.B(n_1037),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1013),
.A2(n_490),
.B(n_537),
.C(n_535),
.Y(n_1192)
);

OR2x6_ASAP7_75t_SL g1193 ( 
.A(n_1031),
.B(n_5),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_1005),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1064),
.Y(n_1195)
);

CKINVDCx8_ASAP7_75t_R g1196 ( 
.A(n_1060),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1191),
.A2(n_980),
.B1(n_1002),
.B2(n_1014),
.Y(n_1197)
);

AOI211x1_ASAP7_75t_L g1198 ( 
.A1(n_1070),
.A2(n_1030),
.B(n_1046),
.C(n_1040),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1078),
.A2(n_910),
.B(n_1047),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1062),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1134),
.B(n_1019),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1134),
.B(n_1077),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_SL g1203 ( 
.A(n_1102),
.B(n_1035),
.C(n_1020),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_SL g1204 ( 
.A1(n_1187),
.A2(n_883),
.B(n_1048),
.C(n_991),
.Y(n_1204)
);

O2A1O1Ixp5_ASAP7_75t_L g1205 ( 
.A1(n_1069),
.A2(n_975),
.B(n_964),
.C(n_984),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1163),
.A2(n_997),
.B(n_1002),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1170),
.B(n_1024),
.Y(n_1207)
);

NAND3xp33_ASAP7_75t_SL g1208 ( 
.A(n_1161),
.B(n_970),
.C(n_1033),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1171),
.A2(n_997),
.B(n_1002),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1091),
.B(n_1026),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_1098),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1122),
.A2(n_964),
.A3(n_1027),
.B(n_1028),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1090),
.A2(n_1018),
.B(n_1011),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1150),
.B(n_984),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1171),
.A2(n_1038),
.B(n_954),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1054),
.A2(n_1028),
.B(n_1027),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1067),
.A2(n_1011),
.B(n_1018),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1092),
.B(n_939),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1191),
.B(n_1135),
.Y(n_1219)
);

AND3x4_ASAP7_75t_L g1220 ( 
.A(n_1129),
.B(n_1021),
.C(n_1012),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1167),
.A2(n_953),
.B1(n_983),
.B2(n_1004),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1053),
.B(n_976),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1140),
.A2(n_903),
.B(n_908),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1068),
.A2(n_1001),
.B(n_903),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1130),
.A2(n_1114),
.B1(n_1108),
.B2(n_1194),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1099),
.A2(n_1001),
.B(n_878),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_1111),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1174),
.A2(n_1006),
.B(n_988),
.C(n_1008),
.Y(n_1228)
);

NOR2xp67_ASAP7_75t_L g1229 ( 
.A(n_1110),
.B(n_983),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1099),
.A2(n_992),
.A3(n_998),
.B(n_1003),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1057),
.A2(n_879),
.B(n_881),
.Y(n_1231)
);

AOI221x1_ASAP7_75t_L g1232 ( 
.A1(n_1183),
.A2(n_909),
.B1(n_881),
.B2(n_895),
.C(n_908),
.Y(n_1232)
);

BUFx5_ASAP7_75t_L g1233 ( 
.A(n_1059),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1158),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1072),
.A2(n_899),
.B(n_879),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1066),
.A2(n_899),
.B(n_895),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1056),
.A2(n_1141),
.B(n_1051),
.Y(n_1237)
);

NAND3x1_ASAP7_75t_L g1238 ( 
.A(n_1184),
.B(n_6),
.C(n_7),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1192),
.A2(n_1029),
.A3(n_919),
.B(n_1023),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1164),
.B(n_944),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1097),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1101),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1146),
.A2(n_914),
.B(n_1023),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1167),
.B(n_1023),
.Y(n_1244)
);

NOR2x1_ASAP7_75t_SL g1245 ( 
.A(n_1063),
.B(n_949),
.Y(n_1245)
);

AOI211x1_ASAP7_75t_L g1246 ( 
.A1(n_1109),
.A2(n_7),
.B(n_9),
.C(n_17),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1190),
.A2(n_1023),
.B(n_978),
.Y(n_1247)
);

NOR3xp33_ASAP7_75t_L g1248 ( 
.A(n_1168),
.B(n_490),
.C(n_978),
.Y(n_1248)
);

AOI31xp67_ASAP7_75t_L g1249 ( 
.A1(n_1073),
.A2(n_990),
.A3(n_982),
.B(n_949),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1089),
.B(n_982),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1113),
.B(n_537),
.Y(n_1251)
);

O2A1O1Ixp5_ASAP7_75t_SL g1252 ( 
.A1(n_1116),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1117),
.A2(n_85),
.B(n_188),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_SL g1254 ( 
.A1(n_1081),
.A2(n_84),
.B(n_187),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1121),
.A2(n_1173),
.B(n_1177),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1058),
.B(n_537),
.Y(n_1256)
);

INVx6_ASAP7_75t_SL g1257 ( 
.A(n_1085),
.Y(n_1257)
);

OAI22x1_ASAP7_75t_L g1258 ( 
.A1(n_1118),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1137),
.B(n_535),
.Y(n_1259)
);

AOI211x1_ASAP7_75t_L g1260 ( 
.A1(n_1095),
.A2(n_22),
.B(n_24),
.C(n_27),
.Y(n_1260)
);

O2A1O1Ixp5_ASAP7_75t_L g1261 ( 
.A1(n_1061),
.A2(n_24),
.B(n_28),
.C(n_30),
.Y(n_1261)
);

AOI221xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1086),
.A2(n_535),
.B1(n_32),
.B2(n_37),
.C(n_38),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1112),
.A2(n_535),
.B(n_42),
.C(n_43),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_SL g1264 ( 
.A(n_1052),
.B(n_535),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1079),
.B(n_28),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1125),
.B(n_46),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1166),
.A2(n_96),
.B(n_133),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1106),
.B(n_46),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1124),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1088),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1120),
.B(n_56),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1154),
.A2(n_105),
.B(n_61),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1098),
.Y(n_1273)
);

INVx5_ASAP7_75t_L g1274 ( 
.A(n_1063),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1082),
.A2(n_109),
.B(n_119),
.Y(n_1275)
);

NOR4xp25_ASAP7_75t_L g1276 ( 
.A(n_1104),
.B(n_60),
.C(n_122),
.D(n_124),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1142),
.A2(n_1083),
.B(n_1100),
.C(n_1162),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1175),
.A2(n_1139),
.B(n_1188),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1103),
.A2(n_1143),
.A3(n_1152),
.B(n_1116),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1147),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1147),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1083),
.A2(n_1152),
.B(n_1127),
.Y(n_1282)
);

AO22x2_ASAP7_75t_L g1283 ( 
.A1(n_1144),
.A2(n_1181),
.B1(n_1151),
.B2(n_1172),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1153),
.A2(n_1176),
.B1(n_1179),
.B2(n_1063),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1127),
.A2(n_1094),
.B(n_1166),
.Y(n_1285)
);

AOI221x1_ASAP7_75t_L g1286 ( 
.A1(n_1185),
.A2(n_1138),
.B1(n_1103),
.B2(n_1107),
.C(n_1143),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1087),
.A2(n_1094),
.B(n_1126),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1148),
.B(n_1145),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1075),
.A2(n_1123),
.B(n_1165),
.Y(n_1289)
);

NAND3xp33_ASAP7_75t_L g1290 ( 
.A(n_1160),
.B(n_1145),
.C(n_1155),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1178),
.A2(n_1182),
.A3(n_1156),
.B(n_1059),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1059),
.B(n_1055),
.Y(n_1292)
);

NOR2xp67_ASAP7_75t_SL g1293 ( 
.A(n_1105),
.B(n_1084),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1131),
.A2(n_1119),
.B(n_1158),
.C(n_1071),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1050),
.A2(n_1149),
.B(n_1071),
.C(n_1096),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1076),
.B(n_1180),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1074),
.B(n_1186),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1059),
.A2(n_1159),
.B(n_1157),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1085),
.A2(n_1169),
.B1(n_1050),
.B2(n_1093),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1156),
.A2(n_1169),
.A3(n_1189),
.B(n_1193),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1080),
.B(n_1128),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_L g1302 ( 
.A(n_1085),
.B(n_1133),
.C(n_1132),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1189),
.A2(n_1093),
.B(n_1096),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1149),
.A2(n_1098),
.B(n_1115),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1136),
.B(n_1169),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1169),
.B(n_1115),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1169),
.A2(n_1132),
.B(n_1133),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1090),
.A2(n_1054),
.B(n_1163),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1170),
.A2(n_715),
.B(n_959),
.C(n_873),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1069),
.A2(n_1163),
.B(n_969),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_R g1311 ( 
.A(n_1060),
.B(n_721),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1170),
.A2(n_715),
.B1(n_959),
.B2(n_725),
.Y(n_1312)
);

AOI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1068),
.A2(n_1163),
.B(n_1065),
.Y(n_1313)
);

AOI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1170),
.A2(n_655),
.B1(n_715),
.B2(n_862),
.C(n_959),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1060),
.B(n_1062),
.Y(n_1315)
);

AND2x6_ASAP7_75t_L g1316 ( 
.A(n_1167),
.B(n_980),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1090),
.A2(n_1054),
.B(n_1163),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1064),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1134),
.B(n_717),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1060),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1170),
.A2(n_959),
.B(n_930),
.C(n_715),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1134),
.B(n_717),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1053),
.B(n_732),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1134),
.B(n_717),
.Y(n_1324)
);

O2A1O1Ixp5_ASAP7_75t_SL g1325 ( 
.A1(n_1068),
.A2(n_1030),
.B(n_1035),
.C(n_1020),
.Y(n_1325)
);

CKINVDCx8_ASAP7_75t_R g1326 ( 
.A(n_1060),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1069),
.A2(n_1163),
.B(n_969),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1060),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1134),
.B(n_717),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1163),
.A2(n_1187),
.A3(n_1122),
.B(n_1099),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1063),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1158),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1150),
.B(n_1074),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1163),
.A2(n_1187),
.A3(n_1122),
.B(n_1099),
.Y(n_1334)
);

NAND2x1_ASAP7_75t_L g1335 ( 
.A(n_1156),
.B(n_984),
.Y(n_1335)
);

INVx4_ASAP7_75t_L g1336 ( 
.A(n_1098),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1069),
.A2(n_1163),
.B(n_969),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1134),
.B(n_717),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1090),
.A2(n_1054),
.B(n_1163),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1069),
.A2(n_1163),
.B(n_969),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1090),
.A2(n_1054),
.B(n_1163),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1134),
.B(n_717),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1069),
.A2(n_1163),
.B(n_969),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1323),
.B(n_1250),
.Y(n_1344)
);

OR2x6_ASAP7_75t_L g1345 ( 
.A(n_1209),
.B(n_1307),
.Y(n_1345)
);

AO32x2_ASAP7_75t_L g1346 ( 
.A1(n_1284),
.A2(n_1197),
.A3(n_1221),
.B1(n_1249),
.B2(n_1252),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1202),
.B(n_1268),
.Y(n_1347)
);

NAND3xp33_ASAP7_75t_L g1348 ( 
.A(n_1312),
.B(n_1314),
.C(n_1321),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1225),
.A2(n_1220),
.B1(n_1329),
.B2(n_1322),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1266),
.A2(n_1271),
.B1(n_1208),
.B2(n_1258),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1309),
.A2(n_1325),
.B(n_1275),
.Y(n_1351)
);

BUFx12f_ASAP7_75t_L g1352 ( 
.A(n_1281),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1341),
.A2(n_1223),
.B(n_1247),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1311),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1278),
.A2(n_1255),
.B(n_1231),
.Y(n_1355)
);

AOI22x1_ASAP7_75t_L g1356 ( 
.A1(n_1283),
.A2(n_1343),
.B1(n_1340),
.B2(n_1337),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1319),
.B(n_1324),
.Y(n_1357)
);

BUFx12f_ASAP7_75t_L g1358 ( 
.A(n_1315),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1313),
.A2(n_1226),
.B(n_1327),
.Y(n_1359)
);

OAI22x1_ASAP7_75t_L g1360 ( 
.A1(n_1299),
.A2(n_1210),
.B1(n_1270),
.B2(n_1302),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1277),
.A2(n_1342),
.B(n_1338),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1274),
.Y(n_1362)
);

OR2x6_ASAP7_75t_L g1363 ( 
.A(n_1298),
.B(n_1305),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1196),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1195),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1235),
.A2(n_1243),
.B(n_1236),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1213),
.A2(n_1253),
.B(n_1287),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1241),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1280),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1282),
.A2(n_1285),
.A3(n_1215),
.B(n_1286),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1242),
.Y(n_1371)
);

NAND2x1p5_ASAP7_75t_L g1372 ( 
.A(n_1274),
.B(n_1331),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1207),
.A2(n_1222),
.B1(n_1201),
.B2(n_1316),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1248),
.A2(n_1224),
.B(n_1204),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1205),
.A2(n_1261),
.B(n_1262),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1272),
.A2(n_1228),
.B(n_1216),
.Y(n_1376)
);

OR2x6_ASAP7_75t_L g1377 ( 
.A(n_1292),
.B(n_1198),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1256),
.A2(n_1265),
.B(n_1251),
.Y(n_1378)
);

A2O1A1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1263),
.A2(n_1203),
.B(n_1290),
.C(n_1269),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1216),
.A2(n_1244),
.B(n_1217),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_1283),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1217),
.A2(n_1267),
.B(n_1259),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1276),
.A2(n_1295),
.B(n_1294),
.Y(n_1383)
);

OR3x4_ASAP7_75t_SL g1384 ( 
.A(n_1238),
.B(n_1257),
.C(n_1301),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_SL g1385 ( 
.A(n_1326),
.B(n_1293),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1227),
.A2(n_1288),
.B1(n_1240),
.B2(n_1328),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1318),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1229),
.B(n_1332),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1289),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1230),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1257),
.A2(n_1320),
.B1(n_1200),
.B2(n_1218),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1316),
.B(n_1230),
.Y(n_1392)
);

INVx8_ASAP7_75t_L g1393 ( 
.A(n_1274),
.Y(n_1393)
);

INVx8_ASAP7_75t_L g1394 ( 
.A(n_1331),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1234),
.B(n_1332),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1303),
.A2(n_1306),
.B(n_1304),
.Y(n_1396)
);

OAI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1264),
.A2(n_1234),
.B1(n_1331),
.B2(n_1297),
.Y(n_1397)
);

OR3x4_ASAP7_75t_SL g1398 ( 
.A(n_1246),
.B(n_1260),
.C(n_1300),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1335),
.A2(n_1233),
.B(n_1291),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1279),
.A2(n_1214),
.B(n_1333),
.C(n_1330),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1316),
.A2(n_1214),
.B(n_1333),
.Y(n_1401)
);

BUFx12f_ASAP7_75t_L g1402 ( 
.A(n_1296),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1233),
.A2(n_1291),
.B(n_1212),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1233),
.A2(n_1291),
.B(n_1212),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1233),
.A2(n_1212),
.B(n_1239),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1300),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1273),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1300),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1273),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1273),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1233),
.A2(n_1239),
.B(n_1330),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1245),
.A2(n_1330),
.B(n_1334),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1211),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_L g1414 ( 
.A(n_1336),
.B(n_1312),
.C(n_1314),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1279),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1310),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1323),
.B(n_904),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1195),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1321),
.B(n_1319),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1323),
.B(n_904),
.Y(n_1421)
);

NOR2xp67_ASAP7_75t_L g1422 ( 
.A(n_1281),
.B(n_721),
.Y(n_1422)
);

AND2x6_ASAP7_75t_SL g1423 ( 
.A(n_1297),
.B(n_1184),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1311),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1195),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1291),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1312),
.A2(n_715),
.B1(n_1321),
.B2(n_1225),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1195),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1312),
.A2(n_715),
.B1(n_1321),
.B2(n_1225),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1250),
.B(n_1302),
.Y(n_1432)
);

OAI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1312),
.A2(n_1314),
.B1(n_1091),
.B2(n_1225),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1280),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1250),
.B(n_1302),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1321),
.B(n_1319),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1206),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1312),
.A2(n_715),
.B1(n_1314),
.B2(n_391),
.Y(n_1439)
);

AO21x2_ASAP7_75t_L g1440 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1206),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1311),
.Y(n_1441)
);

OR2x6_ASAP7_75t_L g1442 ( 
.A(n_1209),
.B(n_1307),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1323),
.B(n_904),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1312),
.A2(n_715),
.B1(n_1321),
.B2(n_1225),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1323),
.B(n_904),
.Y(n_1445)
);

AO21x2_ASAP7_75t_L g1446 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1206),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1202),
.B(n_1219),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_SL g1448 ( 
.A1(n_1245),
.A2(n_1254),
.B(n_1275),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1312),
.A2(n_1321),
.B(n_1309),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1291),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1195),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1195),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1312),
.A2(n_1321),
.B(n_1309),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1237),
.A2(n_1232),
.B(n_1308),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1273),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1280),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1312),
.A2(n_1314),
.B(n_715),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1458)
);

AO21x2_ASAP7_75t_L g1459 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1206),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1312),
.A2(n_715),
.B1(n_1321),
.B2(n_1225),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1237),
.A2(n_1232),
.B(n_1308),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1237),
.A2(n_1232),
.B(n_1308),
.Y(n_1463)
);

BUFx10_ASAP7_75t_L g1464 ( 
.A(n_1297),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1312),
.A2(n_715),
.B1(n_1321),
.B2(n_1225),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1311),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1311),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1311),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1312),
.A2(n_715),
.B1(n_1321),
.B2(n_1225),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1321),
.A2(n_1309),
.B(n_1314),
.C(n_1266),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1237),
.A2(n_1232),
.B(n_1308),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1312),
.B(n_1309),
.Y(n_1476)
);

NOR2xp67_ASAP7_75t_L g1477 ( 
.A(n_1281),
.B(n_721),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1237),
.A2(n_1199),
.B(n_1206),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1274),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1237),
.A2(n_1232),
.B(n_1308),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1308),
.A2(n_1339),
.B(n_1317),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1457),
.A2(n_1460),
.B(n_1428),
.C(n_1466),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1401),
.B(n_1432),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1357),
.B(n_1420),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1430),
.A2(n_1472),
.B(n_1444),
.Y(n_1486)
);

AOI21x1_ASAP7_75t_SL g1487 ( 
.A1(n_1392),
.A2(n_1437),
.B(n_1420),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1344),
.B(n_1347),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1376),
.A2(n_1351),
.B(n_1382),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1357),
.B(n_1437),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1417),
.B(n_1421),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1439),
.A2(n_1433),
.B1(n_1348),
.B2(n_1350),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1443),
.B(n_1445),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1447),
.B(n_1432),
.Y(n_1494)
);

AOI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1433),
.A2(n_1473),
.B1(n_1449),
.B2(n_1453),
.C(n_1476),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1361),
.B(n_1476),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1473),
.B(n_1373),
.Y(n_1497)
);

NOR2xp67_ASAP7_75t_L g1498 ( 
.A(n_1422),
.B(n_1477),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1373),
.B(n_1349),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1381),
.B(n_1400),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1434),
.Y(n_1501)
);

AOI221x1_ASAP7_75t_SL g1502 ( 
.A1(n_1414),
.A2(n_1386),
.B1(n_1397),
.B2(n_1391),
.C(n_1387),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1379),
.A2(n_1350),
.B(n_1400),
.C(n_1397),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1381),
.B(n_1389),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1365),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1441),
.Y(n_1506)
);

INVx3_ASAP7_75t_SL g1507 ( 
.A(n_1364),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1382),
.A2(n_1380),
.B(n_1416),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1363),
.B(n_1415),
.Y(n_1509)
);

CKINVDCx16_ASAP7_75t_R g1510 ( 
.A(n_1441),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1435),
.B(n_1377),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_R g1512 ( 
.A(n_1364),
.B(n_1385),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1435),
.B(n_1377),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1368),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1354),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1363),
.B(n_1415),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1379),
.A2(n_1377),
.B1(n_1469),
.B2(n_1424),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1438),
.A2(n_1440),
.B(n_1459),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1434),
.Y(n_1519)
);

NOR2xp67_ASAP7_75t_L g1520 ( 
.A(n_1352),
.B(n_1402),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1363),
.B(n_1419),
.Y(n_1521)
);

INVx3_ASAP7_75t_SL g1522 ( 
.A(n_1467),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1378),
.B(n_1370),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1395),
.B(n_1388),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1425),
.B(n_1429),
.Y(n_1525)
);

BUFx4_ASAP7_75t_SL g1526 ( 
.A(n_1369),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1378),
.B(n_1370),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1451),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1468),
.A2(n_1402),
.B1(n_1358),
.B2(n_1452),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1362),
.B(n_1480),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1358),
.A2(n_1413),
.B1(n_1369),
.B2(n_1407),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1409),
.B(n_1410),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1378),
.B(n_1370),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1440),
.A2(n_1459),
.B(n_1479),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1360),
.B(n_1407),
.Y(n_1535)
);

OA22x2_ASAP7_75t_L g1536 ( 
.A1(n_1448),
.A2(n_1406),
.B1(n_1408),
.B2(n_1384),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1370),
.B(n_1383),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1390),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1372),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1423),
.A2(n_1352),
.B1(n_1372),
.B2(n_1456),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1396),
.B(n_1399),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1455),
.B(n_1464),
.Y(n_1542)
);

AOI21x1_ASAP7_75t_SL g1543 ( 
.A1(n_1427),
.A2(n_1450),
.B(n_1398),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1345),
.A2(n_1442),
.B(n_1446),
.Y(n_1544)
);

AOI21x1_ASAP7_75t_SL g1545 ( 
.A1(n_1398),
.A2(n_1383),
.B(n_1346),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1380),
.A2(n_1405),
.B(n_1411),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1345),
.A2(n_1442),
.B1(n_1394),
.B2(n_1393),
.Y(n_1547)
);

O2A1O1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1375),
.A2(n_1374),
.B(n_1345),
.C(n_1442),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1393),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1455),
.B(n_1412),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1394),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1412),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1403),
.B(n_1404),
.Y(n_1553)
);

OA21x2_ASAP7_75t_L g1554 ( 
.A1(n_1366),
.A2(n_1353),
.B(n_1367),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1346),
.B(n_1359),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1454),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_SL g1557 ( 
.A1(n_1355),
.A2(n_1462),
.B(n_1481),
.Y(n_1557)
);

AOI221x1_ASAP7_75t_SL g1558 ( 
.A1(n_1346),
.A2(n_1356),
.B1(n_1481),
.B2(n_1462),
.C(n_1474),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1463),
.B(n_1474),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1463),
.A2(n_1418),
.B1(n_1426),
.B2(n_1431),
.Y(n_1560)
);

O2A1O1Ixp5_ASAP7_75t_L g1561 ( 
.A1(n_1436),
.A2(n_1458),
.B(n_1461),
.C(n_1465),
.Y(n_1561)
);

O2A1O1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1470),
.A2(n_1471),
.B(n_1475),
.C(n_1478),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1482),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1376),
.A2(n_1351),
.B(n_1382),
.Y(n_1564)
);

BUFx4_ASAP7_75t_R g1565 ( 
.A(n_1464),
.Y(n_1565)
);

NOR2xp67_ASAP7_75t_L g1566 ( 
.A(n_1422),
.B(n_922),
.Y(n_1566)
);

AOI21x1_ASAP7_75t_SL g1567 ( 
.A1(n_1420),
.A2(n_1437),
.B(n_1266),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1439),
.A2(n_1312),
.B1(n_1225),
.B2(n_1314),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1401),
.B(n_1432),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1357),
.B(n_1420),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1344),
.B(n_1347),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1344),
.B(n_1347),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1344),
.B(n_1347),
.Y(n_1573)
);

AOI21x1_ASAP7_75t_SL g1574 ( 
.A1(n_1392),
.A2(n_1266),
.B(n_1305),
.Y(n_1574)
);

BUFx2_ASAP7_75t_R g1575 ( 
.A(n_1364),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1357),
.B(n_1420),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1371),
.Y(n_1577)
);

NOR2xp67_ASAP7_75t_L g1578 ( 
.A(n_1422),
.B(n_922),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1357),
.B(n_1420),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_1441),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1357),
.B(n_1420),
.Y(n_1581)
);

INVx5_ASAP7_75t_L g1582 ( 
.A(n_1393),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1439),
.A2(n_1312),
.B1(n_1225),
.B2(n_1314),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1538),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1521),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_R g1586 ( 
.A(n_1506),
.B(n_1582),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1509),
.B(n_1516),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1553),
.B(n_1550),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1494),
.B(n_1537),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1505),
.B(n_1514),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1528),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1518),
.A2(n_1534),
.B(n_1557),
.Y(n_1592)
);

AOI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1496),
.A2(n_1492),
.B(n_1563),
.Y(n_1593)
);

AOI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1568),
.A2(n_1583),
.B1(n_1495),
.B2(n_1483),
.C(n_1486),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1553),
.Y(n_1595)
);

OR2x6_ASAP7_75t_L g1596 ( 
.A(n_1544),
.B(n_1548),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1485),
.B(n_1490),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1582),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1559),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1526),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1509),
.B(n_1516),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1503),
.B(n_1547),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1500),
.B(n_1511),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1500),
.B(n_1513),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1508),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1484),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1504),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1504),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1484),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1523),
.B(n_1527),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1555),
.B(n_1489),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_SL g1612 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1533),
.B(n_1489),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1485),
.B(n_1490),
.Y(n_1614)
);

A2O1A1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1483),
.A2(n_1495),
.B(n_1503),
.C(n_1502),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1497),
.A2(n_1499),
.B(n_1517),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1561),
.A2(n_1562),
.B(n_1541),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1546),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1525),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1569),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1564),
.B(n_1577),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1554),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1552),
.Y(n_1623)
);

AO21x2_ASAP7_75t_L g1624 ( 
.A1(n_1558),
.A2(n_1576),
.B(n_1581),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1556),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1570),
.A2(n_1576),
.B1(n_1579),
.B2(n_1581),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1570),
.B(n_1579),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1535),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1539),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1545),
.A2(n_1560),
.B(n_1543),
.Y(n_1630)
);

INVxp67_ASAP7_75t_L g1631 ( 
.A(n_1536),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1567),
.A2(n_1569),
.B(n_1536),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1530),
.Y(n_1633)
);

OR2x6_ASAP7_75t_L g1634 ( 
.A(n_1549),
.B(n_1551),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1595),
.B(n_1549),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1613),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1611),
.B(n_1572),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1584),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1611),
.B(n_1599),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1622),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1624),
.B(n_1571),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1622),
.Y(n_1642)
);

INVxp67_ASAP7_75t_SL g1643 ( 
.A(n_1613),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1584),
.Y(n_1644)
);

OAI33xp33_ASAP7_75t_L g1645 ( 
.A1(n_1591),
.A2(n_1540),
.A3(n_1529),
.B1(n_1531),
.B2(n_1545),
.B3(n_1515),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1624),
.B(n_1573),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1600),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1595),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1624),
.B(n_1488),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_1625),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1621),
.B(n_1491),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1624),
.B(n_1532),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1616),
.A2(n_1512),
.B1(n_1510),
.B2(n_1524),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1587),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1608),
.B(n_1532),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1621),
.B(n_1493),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1618),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1618),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1594),
.B(n_1498),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1605),
.A2(n_1487),
.B(n_1574),
.Y(n_1660)
);

OAI211xp5_ASAP7_75t_L g1661 ( 
.A1(n_1594),
.A2(n_1566),
.B(n_1578),
.C(n_1520),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_SL g1662 ( 
.A(n_1615),
.B(n_1575),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1610),
.B(n_1542),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1601),
.B(n_1501),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1623),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1645),
.B(n_1627),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1638),
.Y(n_1667)
);

OA222x2_ASAP7_75t_L g1668 ( 
.A1(n_1641),
.A2(n_1596),
.B1(n_1602),
.B2(n_1631),
.C1(n_1606),
.C2(n_1598),
.Y(n_1668)
);

OAI211xp5_ASAP7_75t_L g1669 ( 
.A1(n_1659),
.A2(n_1616),
.B(n_1626),
.C(n_1631),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1640),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1659),
.A2(n_1602),
.B1(n_1626),
.B2(n_1630),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1635),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1654),
.Y(n_1673)
);

AOI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1645),
.A2(n_1614),
.B1(n_1597),
.B2(n_1608),
.C(n_1591),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1662),
.A2(n_1602),
.B1(n_1632),
.B2(n_1596),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1638),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1663),
.B(n_1587),
.Y(n_1677)
);

OAI211xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1661),
.A2(n_1614),
.B(n_1597),
.C(n_1627),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1662),
.A2(n_1602),
.B1(n_1632),
.B2(n_1596),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_SL g1680 ( 
.A1(n_1661),
.A2(n_1612),
.B1(n_1602),
.B2(n_1630),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1648),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1653),
.A2(n_1641),
.B1(n_1646),
.B2(n_1649),
.C(n_1652),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1663),
.B(n_1637),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1646),
.A2(n_1619),
.B1(n_1603),
.B2(n_1604),
.C(n_1628),
.Y(n_1684)
);

AO21x2_ASAP7_75t_L g1685 ( 
.A1(n_1652),
.A2(n_1592),
.B(n_1617),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1638),
.Y(n_1686)
);

AOI221xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1649),
.A2(n_1619),
.B1(n_1585),
.B2(n_1603),
.C(n_1607),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1651),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1644),
.Y(n_1689)
);

AOI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1655),
.A2(n_1586),
.B(n_1585),
.C(n_1522),
.Y(n_1690)
);

OAI31xp33_ASAP7_75t_L g1691 ( 
.A1(n_1664),
.A2(n_1609),
.A3(n_1620),
.B(n_1606),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1648),
.B(n_1588),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_1647),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1650),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1636),
.A2(n_1629),
.B1(n_1589),
.B2(n_1633),
.C(n_1590),
.Y(n_1695)
);

OR2x6_ASAP7_75t_L g1696 ( 
.A(n_1635),
.B(n_1634),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1647),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1665),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1642),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_R g1700 ( 
.A(n_1664),
.B(n_1580),
.Y(n_1700)
);

OAI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1636),
.A2(n_1620),
.B1(n_1633),
.B2(n_1519),
.C(n_1593),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1665),
.Y(n_1702)
);

INVx4_ASAP7_75t_L g1703 ( 
.A(n_1693),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1670),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1667),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1666),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1687),
.B(n_1643),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1668),
.B(n_1639),
.Y(n_1708)
);

INVx5_ASAP7_75t_L g1709 ( 
.A(n_1696),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1700),
.B(n_1635),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1700),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1696),
.Y(n_1712)
);

INVx4_ASAP7_75t_SL g1713 ( 
.A(n_1692),
.Y(n_1713)
);

AO21x1_ASAP7_75t_L g1714 ( 
.A1(n_1666),
.A2(n_1643),
.B(n_1593),
.Y(n_1714)
);

AOI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1699),
.A2(n_1658),
.B(n_1657),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1673),
.Y(n_1716)
);

INVx4_ASAP7_75t_SL g1717 ( 
.A(n_1692),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1676),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1686),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1689),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1693),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1698),
.Y(n_1722)
);

INVxp67_ASAP7_75t_SL g1723 ( 
.A(n_1694),
.Y(n_1723)
);

INVx4_ASAP7_75t_SL g1724 ( 
.A(n_1692),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1707),
.B(n_1683),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1715),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1713),
.B(n_1672),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1715),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1706),
.B(n_1702),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1713),
.B(n_1688),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1713),
.B(n_1681),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1705),
.Y(n_1732)
);

NAND2x1p5_ASAP7_75t_L g1733 ( 
.A(n_1709),
.B(n_1660),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1705),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_L g1735 ( 
.A(n_1706),
.B(n_1669),
.C(n_1671),
.D(n_1680),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1722),
.B(n_1684),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1713),
.B(n_1681),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1721),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1713),
.B(n_1637),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1722),
.B(n_1674),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1705),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1713),
.B(n_1717),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1718),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1716),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1718),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1718),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1704),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1713),
.B(n_1637),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1717),
.B(n_1651),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1717),
.B(n_1656),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1719),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1719),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1719),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1717),
.B(n_1656),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1707),
.B(n_1677),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1720),
.Y(n_1756)
);

NOR3xp33_ASAP7_75t_L g1757 ( 
.A(n_1703),
.B(n_1679),
.C(n_1675),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1709),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1716),
.B(n_1682),
.Y(n_1759)
);

AND2x4_ASAP7_75t_SL g1760 ( 
.A(n_1703),
.B(n_1671),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1717),
.B(n_1691),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1704),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1703),
.B(n_1695),
.Y(n_1763)
);

NOR3xp33_ASAP7_75t_L g1764 ( 
.A(n_1703),
.B(n_1678),
.C(n_1701),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1717),
.B(n_1685),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1764),
.B(n_1703),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1738),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1742),
.B(n_1724),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1744),
.Y(n_1770)
);

NOR2xp67_ASAP7_75t_L g1771 ( 
.A(n_1758),
.B(n_1709),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1738),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1732),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1725),
.B(n_1723),
.Y(n_1774)
);

NAND2x1_ASAP7_75t_L g1775 ( 
.A(n_1758),
.B(n_1708),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1732),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1734),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1725),
.B(n_1714),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1761),
.B(n_1724),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1734),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1755),
.B(n_1714),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1741),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1761),
.B(n_1724),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1758),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1739),
.B(n_1724),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1741),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1743),
.Y(n_1787)
);

OR2x6_ASAP7_75t_L g1788 ( 
.A(n_1758),
.B(n_1703),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1739),
.B(n_1724),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1743),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1748),
.B(n_1724),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1748),
.B(n_1724),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1745),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1745),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1746),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1733),
.Y(n_1796)
);

AOI211xp5_ASAP7_75t_L g1797 ( 
.A1(n_1735),
.A2(n_1714),
.B(n_1711),
.C(n_1710),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1746),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1751),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1735),
.A2(n_1710),
.B(n_1711),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1740),
.B(n_1721),
.Y(n_1801)
);

NOR2x1_ASAP7_75t_R g1802 ( 
.A(n_1740),
.B(n_1721),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1766),
.B(n_1749),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1766),
.B(n_1749),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1773),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1769),
.B(n_1750),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1784),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1769),
.B(n_1750),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1773),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1779),
.B(n_1754),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1800),
.B(n_1759),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1779),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1784),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1776),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1770),
.B(n_1759),
.Y(n_1815)
);

NOR2x1_ASAP7_75t_L g1816 ( 
.A(n_1767),
.B(n_1721),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1783),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_L g1818 ( 
.A(n_1797),
.B(n_1757),
.C(n_1763),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1776),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1774),
.B(n_1755),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1780),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1774),
.B(n_1729),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1783),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1801),
.B(n_1736),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1778),
.B(n_1729),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1780),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1778),
.B(n_1736),
.Y(n_1827)
);

INVxp67_ASAP7_75t_L g1828 ( 
.A(n_1802),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1782),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1785),
.B(n_1754),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1828),
.B(n_1811),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1818),
.A2(n_1775),
.B1(n_1781),
.B2(n_1708),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1827),
.A2(n_1775),
.B1(n_1781),
.B2(n_1708),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1809),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1809),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1814),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1820),
.B(n_1768),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1812),
.B(n_1768),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1824),
.A2(n_1760),
.B(n_1771),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1820),
.B(n_1772),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1810),
.A2(n_1760),
.B1(n_1709),
.B2(n_1712),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_SL g1842 ( 
.A(n_1817),
.B(n_1690),
.C(n_1772),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1815),
.A2(n_1760),
.B1(n_1798),
.B2(n_1799),
.C(n_1795),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1814),
.Y(n_1844)
);

INVx1_ASAP7_75t_SL g1845 ( 
.A(n_1823),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1826),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1826),
.Y(n_1847)
);

AOI21xp33_ASAP7_75t_SL g1848 ( 
.A1(n_1827),
.A2(n_1507),
.B(n_1788),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1803),
.B(n_1708),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1829),
.Y(n_1850)
);

INVx2_ASAP7_75t_SL g1851 ( 
.A(n_1837),
.Y(n_1851)
);

INVx4_ASAP7_75t_L g1852 ( 
.A(n_1840),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1831),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1832),
.A2(n_1825),
.B1(n_1822),
.B2(n_1805),
.C(n_1819),
.Y(n_1854)
);

NOR2x1_ASAP7_75t_L g1855 ( 
.A(n_1845),
.B(n_1816),
.Y(n_1855)
);

CKINVDCx20_ASAP7_75t_R g1856 ( 
.A(n_1845),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1838),
.B(n_1810),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1834),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1843),
.B(n_1803),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1848),
.B(n_1806),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1849),
.B(n_1804),
.Y(n_1861)
);

NAND3xp33_ASAP7_75t_L g1862 ( 
.A(n_1855),
.B(n_1833),
.C(n_1841),
.Y(n_1862)
);

AOI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1854),
.A2(n_1842),
.B1(n_1847),
.B2(n_1846),
.C(n_1844),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1857),
.B(n_1806),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1859),
.A2(n_1839),
.B(n_1825),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1852),
.B(n_1804),
.Y(n_1866)
);

NAND4xp25_ASAP7_75t_L g1867 ( 
.A(n_1860),
.B(n_1850),
.C(n_1836),
.D(n_1835),
.Y(n_1867)
);

A2O1A1Ixp33_ASAP7_75t_L g1868 ( 
.A1(n_1853),
.A2(n_1856),
.B(n_1851),
.C(n_1861),
.Y(n_1868)
);

NAND4xp25_ASAP7_75t_L g1869 ( 
.A(n_1852),
.B(n_1822),
.C(n_1808),
.D(n_1830),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1858),
.A2(n_1788),
.B(n_1807),
.Y(n_1870)
);

AOI21xp33_ASAP7_75t_SL g1871 ( 
.A1(n_1851),
.A2(n_1813),
.B(n_1807),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1862),
.A2(n_1813),
.B(n_1808),
.Y(n_1872)
);

INVxp67_ASAP7_75t_SL g1873 ( 
.A(n_1866),
.Y(n_1873)
);

OAI321xp33_ASAP7_75t_L g1874 ( 
.A1(n_1869),
.A2(n_1788),
.A3(n_1830),
.B1(n_1829),
.B2(n_1821),
.C(n_1785),
.Y(n_1874)
);

AND3x1_ASAP7_75t_L g1875 ( 
.A(n_1868),
.B(n_1791),
.C(n_1789),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1864),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1871),
.B(n_1789),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1876),
.B(n_1867),
.Y(n_1878)
);

OAI32xp33_ASAP7_75t_L g1879 ( 
.A1(n_1872),
.A2(n_1863),
.A3(n_1796),
.B1(n_1733),
.B2(n_1782),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1873),
.B(n_1865),
.Y(n_1880)
);

AOI21xp33_ASAP7_75t_SL g1881 ( 
.A1(n_1877),
.A2(n_1788),
.B(n_1870),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1877),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1875),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1874),
.Y(n_1884)
);

AOI322xp5_ASAP7_75t_L g1885 ( 
.A1(n_1884),
.A2(n_1796),
.A3(n_1794),
.B1(n_1786),
.B2(n_1777),
.C1(n_1793),
.C2(n_1790),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_R g1886 ( 
.A(n_1880),
.B(n_1697),
.Y(n_1886)
);

AOI211xp5_ASAP7_75t_L g1887 ( 
.A1(n_1881),
.A2(n_1792),
.B(n_1791),
.C(n_1787),
.Y(n_1887)
);

INVx2_ASAP7_75t_SL g1888 ( 
.A(n_1878),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1883),
.B(n_1792),
.Y(n_1889)
);

AND4x1_ASAP7_75t_L g1890 ( 
.A(n_1889),
.B(n_1882),
.C(n_1879),
.D(n_1575),
.Y(n_1890)
);

AOI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1888),
.A2(n_1765),
.B1(n_1727),
.B2(n_1730),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1886),
.B(n_1697),
.Y(n_1892)
);

INVx2_ASAP7_75t_SL g1893 ( 
.A(n_1892),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1893),
.B(n_1891),
.Y(n_1894)
);

BUFx2_ASAP7_75t_L g1895 ( 
.A(n_1894),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1894),
.B(n_1887),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1895),
.B(n_1890),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1896),
.B(n_1885),
.Y(n_1898)
);

AOI22x1_ASAP7_75t_L g1899 ( 
.A1(n_1898),
.A2(n_1765),
.B1(n_1565),
.B2(n_1726),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1897),
.A2(n_1765),
.B1(n_1733),
.B2(n_1712),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1765),
.B1(n_1731),
.B2(n_1737),
.Y(n_1901)
);

OAI22x1_ASAP7_75t_L g1902 ( 
.A1(n_1901),
.A2(n_1899),
.B1(n_1762),
.B2(n_1747),
.Y(n_1902)
);

AOI21xp33_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1728),
.B(n_1726),
.Y(n_1903)
);

AO21x2_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1762),
.B(n_1747),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1904),
.A2(n_1762),
.B1(n_1747),
.B2(n_1753),
.Y(n_1905)
);

AOI211xp5_ASAP7_75t_L g1906 ( 
.A1(n_1905),
.A2(n_1751),
.B(n_1752),
.C(n_1756),
.Y(n_1906)
);


endmodule