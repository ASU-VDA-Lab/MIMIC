module fake_jpeg_8230_n_110 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_20),
.B1(n_12),
.B2(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_11),
.B(n_21),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_35),
.B(n_42),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_20),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.C(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_15),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_12),
.B1(n_19),
.B2(n_16),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_14),
.B(n_18),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_14),
.B(n_18),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_40),
.B1(n_33),
.B2(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_66),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_40),
.B1(n_29),
.B2(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_65),
.Y(n_69)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_72),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_44),
.C(n_51),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_61),
.C(n_58),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_48),
.B(n_50),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_57),
.B(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_65),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_57),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_82),
.C(n_76),
.Y(n_88)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_13),
.B(n_23),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_13),
.B1(n_15),
.B2(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_82),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_88),
.C(n_13),
.Y(n_96)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_91),
.B1(n_23),
.B2(n_2),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_68),
.B1(n_71),
.B2(n_41),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_13),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_90),
.B(n_92),
.Y(n_98)
);

OAI322xp33_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_83),
.A3(n_79),
.B1(n_13),
.B2(n_23),
.C1(n_0),
.C2(n_2),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_1),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_99),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_91),
.B(n_23),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_95),
.B1(n_4),
.B2(n_5),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_104),
.B(n_8),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_106),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_103),
.C(n_8),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_107),
.Y(n_110)
);


endmodule