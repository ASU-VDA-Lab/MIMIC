module fake_aes_4436_n_757 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_757);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_757;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_627;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g95 ( .A(n_53), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_52), .Y(n_97) );
XNOR2xp5_ASAP7_75t_L g98 ( .A(n_14), .B(n_84), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_32), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_44), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_0), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_0), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_48), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_70), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_83), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_56), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_4), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_68), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_93), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_86), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_74), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_16), .Y(n_112) );
NOR2xp67_ASAP7_75t_L g113 ( .A(n_47), .B(n_59), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_90), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_6), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_25), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_20), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_78), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_10), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_11), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_33), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_18), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_60), .Y(n_124) );
INVxp67_ASAP7_75t_L g125 ( .A(n_22), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_51), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_82), .Y(n_127) );
INVxp67_ASAP7_75t_SL g128 ( .A(n_16), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_31), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_11), .B(n_41), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_118), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_99), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_99), .Y(n_133) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_111), .B(n_21), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_108), .B(n_1), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_108), .Y(n_136) );
INVx6_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_117), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_118), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_118), .Y(n_140) );
OAI22xp33_ASAP7_75t_L g141 ( .A1(n_117), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_122), .B(n_5), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_95), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_111), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g145 ( .A1(n_122), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_102), .B(n_7), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_109), .B(n_8), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_101), .B(n_96), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_102), .B(n_9), .Y(n_149) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_109), .A2(n_49), .B(n_92), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_112), .B(n_9), .Y(n_151) );
INVx6_ASAP7_75t_L g152 ( .A(n_118), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_132), .B(n_116), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_137), .Y(n_154) );
INVx2_ASAP7_75t_SL g155 ( .A(n_144), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_148), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_137), .Y(n_157) );
OR2x6_ASAP7_75t_L g158 ( .A(n_142), .B(n_112), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_137), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_132), .B(n_107), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_133), .B(n_116), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_133), .B(n_125), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
INVxp67_ASAP7_75t_L g165 ( .A(n_148), .Y(n_165) );
NOR2xp33_ASAP7_75t_SL g166 ( .A(n_134), .B(n_106), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_134), .A2(n_120), .B1(n_115), .B2(n_119), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_134), .B(n_136), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_139), .Y(n_171) );
OR2x6_ASAP7_75t_L g172 ( .A(n_142), .B(n_115), .Y(n_172) );
AND2x6_ASAP7_75t_L g173 ( .A(n_151), .B(n_110), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_142), .Y(n_174) );
OR2x6_ASAP7_75t_L g175 ( .A(n_145), .B(n_146), .Y(n_175) );
OAI22xp33_ASAP7_75t_L g176 ( .A1(n_138), .A2(n_119), .B1(n_120), .B2(n_128), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
AO22x2_ASAP7_75t_L g179 ( .A1(n_145), .A2(n_129), .B1(n_127), .B2(n_126), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_143), .B(n_123), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g183 ( .A1(n_138), .A2(n_98), .B1(n_130), .B2(n_127), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_143), .B(n_123), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_149), .Y(n_185) );
AND2x6_ASAP7_75t_L g186 ( .A(n_149), .B(n_110), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_152), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_135), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_180), .B(n_100), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_185), .B(n_147), .Y(n_190) );
AOI22x1_ASAP7_75t_L g191 ( .A1(n_154), .A2(n_131), .B1(n_140), .B2(n_139), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_161), .B(n_103), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_165), .A2(n_141), .B(n_124), .C(n_126), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_166), .B(n_150), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_181), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_173), .B(n_104), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_186), .B(n_124), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_170), .A2(n_141), .B1(n_98), .B2(n_129), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_173), .B(n_105), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_173), .A2(n_150), .B1(n_121), .B2(n_97), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_173), .B(n_114), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_173), .B(n_150), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_159), .B(n_113), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_181), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_186), .B(n_150), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_169), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_168), .A2(n_150), .B1(n_140), .B2(n_131), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_175), .A2(n_118), .B1(n_140), .B2(n_131), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_184), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_184), .Y(n_213) );
NOR2xp67_ASAP7_75t_L g214 ( .A(n_164), .B(n_54), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_175), .A2(n_152), .B1(n_139), .B2(n_13), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_188), .B(n_152), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_163), .B(n_152), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_177), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_163), .B(n_152), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_153), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_175), .A2(n_139), .B1(n_12), .B2(n_13), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_153), .A2(n_139), .B(n_50), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_162), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_155), .B(n_139), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_165), .B(n_46), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_186), .B(n_55), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_186), .B(n_10), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_203), .A2(n_162), .B(n_158), .Y(n_229) );
AO32x1_ASAP7_75t_L g230 ( .A1(n_208), .A2(n_182), .A3(n_187), .B1(n_183), .B2(n_156), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_197), .B(n_174), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_190), .B(n_172), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_189), .B(n_172), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_206), .A2(n_172), .B(n_158), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_194), .A2(n_158), .B1(n_179), .B2(n_176), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_194), .B(n_182), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_221), .A2(n_179), .B1(n_176), .B2(n_186), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_206), .A2(n_171), .B(n_167), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_192), .B(n_12), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_216), .A2(n_171), .B(n_167), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_208), .A2(n_171), .B(n_167), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_196), .B(n_179), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_227), .Y(n_243) );
OR2x6_ASAP7_75t_SL g244 ( .A(n_199), .B(n_14), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_199), .B(n_15), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_196), .A2(n_171), .B(n_58), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_200), .B(n_15), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_205), .A2(n_61), .B(n_91), .Y(n_248) );
AO32x1_ASAP7_75t_L g249 ( .A1(n_205), .A2(n_213), .A3(n_212), .B1(n_195), .B2(n_209), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_212), .A2(n_17), .B(n_18), .C(n_19), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_202), .B(n_17), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_209), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_214), .B(n_19), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_209), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_213), .B(n_20), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_198), .A2(n_23), .B1(n_24), .B2(n_26), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_201), .A2(n_27), .B(n_28), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_204), .B(n_94), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_220), .A2(n_29), .B(n_30), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_210), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_236), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_249), .A2(n_195), .B(n_219), .Y(n_262) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_238), .A2(n_222), .B(n_214), .Y(n_263) );
AND2x6_ASAP7_75t_L g264 ( .A(n_258), .B(n_223), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_249), .A2(n_195), .B(n_217), .Y(n_266) );
AO31x2_ASAP7_75t_L g267 ( .A1(n_241), .A2(n_198), .A3(n_226), .B(n_218), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_240), .A2(n_222), .B(n_226), .Y(n_268) );
AOI21x1_ASAP7_75t_L g269 ( .A1(n_253), .A2(n_225), .B(n_218), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_249), .A2(n_223), .B(n_220), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_246), .A2(n_218), .B(n_210), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_233), .B(n_193), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_230), .A2(n_224), .B(n_211), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_239), .A2(n_215), .B(n_210), .C(n_207), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_258), .Y(n_275) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_257), .A2(n_228), .B(n_191), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_234), .B(n_207), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_248), .A2(n_228), .B(n_207), .Y(n_278) );
AO31x2_ASAP7_75t_L g279 ( .A1(n_250), .A2(n_228), .A3(n_191), .B(n_207), .Y(n_279) );
AOI221x1_ASAP7_75t_L g280 ( .A1(n_237), .A2(n_34), .B1(n_35), .B2(n_36), .C(n_37), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_229), .A2(n_38), .B(n_39), .C(n_40), .Y(n_281) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_259), .A2(n_42), .B(n_43), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_278), .A2(n_255), .B(n_256), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_272), .B(n_235), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_265), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_265), .B(n_245), .Y(n_286) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_270), .A2(n_242), .B(n_247), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_275), .B(n_231), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_275), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_264), .B(n_244), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_274), .A2(n_256), .B1(n_243), .B2(n_270), .Y(n_291) );
OR2x6_ASAP7_75t_L g292 ( .A(n_261), .B(n_251), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_262), .A2(n_230), .B(n_254), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_261), .B(n_260), .Y(n_294) );
AO31x2_ASAP7_75t_L g295 ( .A1(n_262), .A2(n_230), .A3(n_252), .B(n_62), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_264), .B(n_45), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_263), .A2(n_57), .B(n_63), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g299 ( .A1(n_266), .A2(n_64), .B(n_65), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_267), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_264), .B(n_89), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_264), .A2(n_66), .B1(n_67), .B2(n_69), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_271), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_267), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_282), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_300), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_293), .A2(n_266), .B(n_273), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_300), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_301), .B(n_267), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_305), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_305), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_285), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_289), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_304), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_287), .B(n_279), .Y(n_318) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_291), .A2(n_273), .B(n_268), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_304), .Y(n_320) );
NOR2x1_ASAP7_75t_SL g321 ( .A(n_292), .B(n_269), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_284), .B(n_279), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_304), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_296), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_287), .B(n_279), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_291), .A2(n_281), .B(n_280), .Y(n_326) );
AO21x2_ASAP7_75t_L g327 ( .A1(n_299), .A2(n_276), .B(n_72), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_306), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_295), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_295), .B(n_276), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_295), .B(n_71), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_286), .B(n_73), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_295), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_294), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_298), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_306), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_306), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_298), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_299), .Y(n_341) );
AO21x2_ASAP7_75t_L g342 ( .A1(n_283), .A2(n_75), .B(n_77), .Y(n_342) );
OA21x2_ASAP7_75t_L g343 ( .A1(n_283), .A2(n_79), .B(n_80), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_290), .A2(n_81), .B1(n_85), .B2(n_87), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_303), .A2(n_88), .B1(n_292), .B2(n_288), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_307), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_311), .B(n_294), .Y(n_347) );
INVxp67_ASAP7_75t_SL g348 ( .A(n_314), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_307), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_322), .B(n_309), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_314), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
INVx3_ASAP7_75t_L g353 ( .A(n_323), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_309), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_323), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_311), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_312), .Y(n_358) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_317), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_312), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_312), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_312), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_322), .B(n_292), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_318), .B(n_325), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_323), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_323), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_316), .Y(n_368) );
AND2x4_ASAP7_75t_SL g369 ( .A(n_335), .B(n_292), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_318), .B(n_325), .Y(n_370) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_342), .B(n_297), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_324), .B(n_292), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_318), .B(n_306), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_324), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_317), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_313), .B(n_306), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_325), .B(n_302), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_313), .B(n_315), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_320), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_315), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_310), .B(n_330), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_320), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_310), .Y(n_385) );
NAND2x1_ASAP7_75t_L g386 ( .A(n_310), .B(n_320), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_323), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_310), .B(n_330), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_310), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_320), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_308), .B(n_336), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_336), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_329), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_332), .B(n_334), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_338), .Y(n_395) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_323), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_338), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_338), .Y(n_398) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_323), .Y(n_399) );
AO21x2_ASAP7_75t_L g400 ( .A1(n_337), .A2(n_340), .B(n_326), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_329), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_308), .B(n_334), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_338), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_329), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_332), .B(n_329), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_332), .B(n_334), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_334), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_308), .B(n_331), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_308), .B(n_331), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_337), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_308), .B(n_331), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_323), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_341), .B(n_333), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_365), .B(n_319), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_346), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_352), .Y(n_416) );
AND2x4_ASAP7_75t_SL g417 ( .A(n_347), .B(n_344), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_376), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_346), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_365), .B(n_319), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_370), .B(n_319), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_351), .B(n_333), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g423 ( .A(n_351), .B(n_345), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_348), .B(n_341), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_349), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_347), .B(n_319), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_349), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_376), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_370), .B(n_319), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_383), .B(n_339), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_383), .B(n_339), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_382), .B(n_345), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_388), .B(n_339), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_388), .B(n_339), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_354), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_382), .B(n_326), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_352), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_408), .B(n_328), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_354), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_408), .B(n_328), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_409), .B(n_328), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_363), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_363), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_352), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_385), .B(n_321), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_368), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_368), .Y(n_447) );
INVx5_ASAP7_75t_L g448 ( .A(n_387), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_379), .B(n_326), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_409), .B(n_340), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_360), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_350), .B(n_342), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_385), .B(n_321), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_379), .B(n_326), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_386), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_375), .B(n_326), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_411), .B(n_342), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_375), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_411), .B(n_342), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_378), .B(n_342), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_378), .B(n_327), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_394), .B(n_327), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_355), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_389), .B(n_327), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_394), .B(n_327), .Y(n_465) );
AOI21xp33_ASAP7_75t_SL g466 ( .A1(n_374), .A2(n_344), .B(n_343), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_360), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_405), .B(n_327), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_405), .B(n_343), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_350), .B(n_343), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_380), .B(n_343), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_406), .B(n_343), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_355), .B(n_343), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_357), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_360), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_357), .B(n_361), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_406), .B(n_373), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_358), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_358), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_373), .B(n_389), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_359), .B(n_369), .Y(n_481) );
NAND2x1p5_ASAP7_75t_SL g482 ( .A(n_371), .B(n_398), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_361), .B(n_362), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_362), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_393), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_364), .B(n_372), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_392), .B(n_384), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_410), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_390), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_410), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_372), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_393), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_401), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_401), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_364), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_392), .B(n_384), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_404), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_386), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_369), .A2(n_413), .B1(n_391), .B2(n_371), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_404), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_407), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_391), .B(n_402), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_384), .B(n_407), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_395), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_395), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_377), .Y(n_506) );
BUFx3_ASAP7_75t_L g507 ( .A(n_369), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_377), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_489), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_477), .B(n_402), .Y(n_510) );
AND3x2_ASAP7_75t_L g511 ( .A(n_423), .B(n_381), .C(n_399), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_477), .B(n_400), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_480), .B(n_353), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_485), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_415), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_502), .B(n_397), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_480), .B(n_353), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_502), .B(n_397), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_485), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_414), .B(n_400), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_450), .B(n_413), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_450), .B(n_400), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_428), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_495), .B(n_491), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_415), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_414), .B(n_400), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_419), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_424), .B(n_403), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_419), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_420), .B(n_403), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_420), .B(n_403), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_492), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_425), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_438), .B(n_395), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_421), .B(n_398), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_438), .B(n_398), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_421), .B(n_397), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_486), .B(n_353), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_425), .B(n_353), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_440), .B(n_399), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_440), .B(n_356), .Y(n_541) );
OAI21xp33_ASAP7_75t_L g542 ( .A1(n_429), .A2(n_396), .B(n_412), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_427), .B(n_356), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_445), .B(n_412), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_430), .B(n_356), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_427), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_435), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_430), .B(n_356), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_431), .B(n_366), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_431), .B(n_366), .Y(n_550) );
NAND2x2_ASAP7_75t_L g551 ( .A(n_507), .B(n_412), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_432), .B(n_366), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_435), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_439), .B(n_366), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_439), .B(n_367), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_442), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_441), .B(n_367), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_441), .B(n_367), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_442), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_418), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_433), .B(n_367), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_492), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_443), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_433), .B(n_387), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_443), .B(n_387), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_434), .B(n_387), .Y(n_566) );
INVx3_ASAP7_75t_L g567 ( .A(n_455), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_434), .B(n_387), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_418), .Y(n_569) );
INVx3_ASAP7_75t_SL g570 ( .A(n_481), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_446), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_483), .B(n_387), .Y(n_572) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_500), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_446), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_507), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_500), .Y(n_576) );
OR2x6_ASAP7_75t_L g577 ( .A(n_498), .B(n_455), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_483), .B(n_487), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_503), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_503), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_476), .B(n_426), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_447), .B(n_458), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_504), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_447), .Y(n_584) );
OAI211xp5_ASAP7_75t_L g585 ( .A1(n_499), .A2(n_498), .B(n_466), .C(n_459), .Y(n_585) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_455), .B(n_422), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_458), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_449), .B(n_454), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_457), .B(n_459), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_488), .Y(n_590) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_448), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_457), .B(n_460), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_487), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_488), .Y(n_594) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_504), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_490), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_460), .B(n_461), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_496), .B(n_508), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_496), .B(n_508), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_471), .A2(n_473), .B(n_470), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_506), .B(n_490), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_506), .B(n_493), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_505), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_588), .B(n_436), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_570), .A2(n_452), .B1(n_497), .B2(n_494), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_509), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_588), .B(n_456), .Y(n_607) );
AOI21xp33_ASAP7_75t_L g608 ( .A1(n_585), .A2(n_452), .B(n_445), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_509), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_570), .B(n_448), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_551), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_512), .B(n_461), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_560), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_602), .Y(n_614) );
OAI32xp33_ASAP7_75t_L g615 ( .A1(n_551), .A2(n_493), .A3(n_501), .B1(n_497), .B2(n_494), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_601), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_598), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_552), .A2(n_417), .B1(n_445), .B2(n_453), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_512), .B(n_501), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_599), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_583), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_576), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_586), .A2(n_474), .B1(n_479), .B2(n_478), .C(n_463), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_582), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_580), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_589), .B(n_474), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_580), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_515), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_510), .B(n_453), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_560), .B(n_463), .C(n_479), .Y(n_630) );
NOR2x1p5_ASAP7_75t_L g631 ( .A(n_567), .B(n_453), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_525), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_510), .B(n_478), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_589), .B(n_484), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_578), .B(n_465), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_576), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_573), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_569), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_521), .B(n_465), .Y(n_639) );
BUFx2_ASAP7_75t_SL g640 ( .A(n_575), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_527), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_523), .B(n_468), .Y(n_642) );
NOR2xp67_ASAP7_75t_L g643 ( .A(n_569), .B(n_448), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_529), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_522), .B(n_505), .C(n_464), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_552), .A2(n_417), .B1(n_468), .B2(n_462), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_513), .B(n_462), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_533), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_546), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_544), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_542), .A2(n_472), .B(n_469), .C(n_464), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_579), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_592), .B(n_469), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_592), .B(n_472), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_538), .A2(n_464), .B1(n_437), .B2(n_444), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_593), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_583), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_603), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_517), .B(n_535), .Y(n_659) );
NAND3xp33_ASAP7_75t_SL g660 ( .A(n_524), .B(n_416), .C(n_437), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_535), .B(n_416), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_537), .B(n_444), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_537), .B(n_451), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_581), .B(n_451), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_541), .B(n_467), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_603), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_530), .B(n_531), .Y(n_667) );
INVx4_ASAP7_75t_L g668 ( .A(n_511), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_516), .B(n_467), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_541), .B(n_475), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_604), .B(n_526), .Y(n_671) );
OAI322xp33_ASAP7_75t_SL g672 ( .A1(n_653), .A2(n_556), .A3(n_559), .B1(n_563), .B2(n_553), .C1(n_571), .C2(n_574), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_668), .B(n_567), .Y(n_673) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_607), .A2(n_526), .B1(n_520), .B2(n_597), .C1(n_540), .C2(n_547), .Y(n_674) );
AOI321xp33_ASAP7_75t_L g675 ( .A1(n_651), .A2(n_520), .A3(n_597), .B1(n_600), .B2(n_540), .C(n_558), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_616), .B(n_528), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_L g677 ( .A1(n_643), .A2(n_544), .B(n_591), .C(n_567), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_637), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_650), .B(n_557), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_606), .B(n_518), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_637), .Y(n_681) );
OAI22xp33_ASAP7_75t_SL g682 ( .A1(n_610), .A2(n_668), .B1(n_577), .B2(n_613), .Y(n_682) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_622), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_609), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_624), .B(n_596), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_640), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_610), .A2(n_577), .B1(n_544), .B2(n_536), .Y(n_687) );
INVx1_ASAP7_75t_SL g688 ( .A(n_652), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_618), .A2(n_577), .B1(n_534), .B2(n_595), .Y(n_689) );
INVxp67_ASAP7_75t_L g690 ( .A(n_609), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_656), .Y(n_691) );
INVx1_ASAP7_75t_SL g692 ( .A(n_633), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_622), .Y(n_693) );
OAI21xp5_ASAP7_75t_SL g694 ( .A1(n_611), .A2(n_511), .B(n_572), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_608), .A2(n_594), .B1(n_590), .B2(n_587), .C(n_584), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_617), .B(n_543), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_645), .A2(n_558), .B1(n_557), .B2(n_568), .Y(n_697) );
INVx2_ASAP7_75t_SL g698 ( .A(n_629), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_628), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_632), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_650), .B(n_561), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_641), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_644), .Y(n_703) );
OAI222xp33_ASAP7_75t_L g704 ( .A1(n_623), .A2(n_561), .B1(n_549), .B2(n_550), .C1(n_548), .C2(n_545), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_648), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_646), .A2(n_568), .B1(n_566), .B2(n_564), .Y(n_706) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_615), .A2(n_566), .B1(n_564), .B2(n_448), .Y(n_707) );
INVx2_ASAP7_75t_SL g708 ( .A(n_669), .Y(n_708) );
OAI22xp33_ASAP7_75t_SL g709 ( .A1(n_686), .A2(n_613), .B1(n_638), .B2(n_611), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_678), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_672), .A2(n_605), .B1(n_620), .B2(n_614), .C(n_638), .Y(n_711) );
AOI21xp33_ASAP7_75t_L g712 ( .A1(n_682), .A2(n_605), .B(n_630), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_697), .B(n_635), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_704), .A2(n_625), .B1(n_627), .B2(n_660), .C(n_645), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_675), .B(n_636), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_674), .A2(n_660), .B1(n_642), .B2(n_639), .Y(n_716) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_683), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_699), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_694), .A2(n_631), .B(n_636), .C(n_626), .Y(n_719) );
OAI221xp5_ASAP7_75t_SL g720 ( .A1(n_697), .A2(n_655), .B1(n_612), .B2(n_634), .C(n_619), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_696), .B(n_647), .Y(n_721) );
AOI21xp33_ASAP7_75t_SL g722 ( .A1(n_687), .A2(n_482), .B(n_654), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_700), .Y(n_723) );
AOI322xp5_ASAP7_75t_L g724 ( .A1(n_692), .A2(n_659), .A3(n_663), .B1(n_662), .B2(n_661), .C1(n_665), .C2(n_670), .Y(n_724) );
AOI32xp33_ASAP7_75t_L g725 ( .A1(n_688), .A2(n_649), .A3(n_664), .B1(n_667), .B2(n_658), .Y(n_725) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_707), .A2(n_448), .B1(n_666), .B2(n_658), .Y(n_726) );
BUFx3_ASAP7_75t_L g727 ( .A(n_691), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_685), .B(n_666), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_702), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_696), .B(n_657), .Y(n_730) );
NAND5xp2_ASAP7_75t_L g731 ( .A(n_677), .B(n_554), .C(n_555), .D(n_539), .E(n_565), .Y(n_731) );
NAND3xp33_ASAP7_75t_L g732 ( .A(n_695), .B(n_657), .C(n_621), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_689), .A2(n_621), .B1(n_514), .B2(n_519), .C(n_532), .Y(n_733) );
NOR4xp25_ASAP7_75t_L g734 ( .A(n_690), .B(n_514), .C(n_519), .D(n_532), .Y(n_734) );
OAI221xp5_ASAP7_75t_SL g735 ( .A1(n_706), .A2(n_475), .B1(n_482), .B2(n_562), .C(n_677), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_681), .B(n_562), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_676), .A2(n_671), .B1(n_685), .B2(n_708), .Y(n_737) );
OAI211xp5_ASAP7_75t_SL g738 ( .A1(n_673), .A2(n_684), .B(n_683), .C(n_703), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_714), .A2(n_715), .B1(n_722), .B2(n_712), .C(n_720), .Y(n_739) );
AOI211xp5_ASAP7_75t_L g740 ( .A1(n_709), .A2(n_735), .B(n_726), .C(n_719), .Y(n_740) );
NAND4xp25_ASAP7_75t_SL g741 ( .A(n_716), .B(n_725), .C(n_724), .D(n_711), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g742 ( .A1(n_716), .A2(n_738), .B1(n_734), .B2(n_733), .C(n_717), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_673), .A2(n_717), .B(n_727), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_743), .B(n_718), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_741), .Y(n_745) );
INVxp67_ASAP7_75t_L g746 ( .A(n_739), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_745), .B(n_746), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_744), .A2(n_742), .B1(n_740), .B2(n_713), .Y(n_748) );
NOR3x1_ASAP7_75t_L g749 ( .A(n_747), .B(n_744), .C(n_732), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_748), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_749), .Y(n_751) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_750), .A2(n_737), .B1(n_729), .B2(n_723), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_751), .A2(n_710), .B1(n_721), .B2(n_730), .Y(n_753) );
AO21x1_ASAP7_75t_L g754 ( .A1(n_753), .A2(n_752), .B(n_728), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_754), .A2(n_728), .B(n_693), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_755), .A2(n_676), .B1(n_698), .B2(n_701), .Y(n_756) );
AOI222xp33_ASAP7_75t_L g757 ( .A1(n_756), .A2(n_736), .B1(n_705), .B2(n_680), .C1(n_679), .C2(n_731), .Y(n_757) );
endmodule