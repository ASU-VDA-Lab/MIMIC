module real_aes_16003_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_735;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_0), .Y(n_511) );
AND2x4_ASAP7_75t_L g868 ( .A(n_1), .B(n_869), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_2), .A2(n_4), .B1(n_180), .B2(n_181), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_3), .A2(n_20), .B1(n_131), .B2(n_133), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_5), .A2(n_52), .B1(n_198), .B2(n_199), .Y(n_197) );
BUFx3_ASAP7_75t_L g541 ( .A(n_6), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_7), .A2(n_13), .B1(n_138), .B2(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g869 ( .A(n_8), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_9), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_10), .B(n_178), .Y(n_547) );
OR2x2_ASAP7_75t_L g818 ( .A(n_11), .B(n_32), .Y(n_818) );
BUFx2_ASAP7_75t_L g874 ( .A(n_11), .Y(n_874) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_12), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_14), .B(n_195), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_15), .B(n_216), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_16), .A2(n_86), .B1(n_131), .B2(n_195), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_17), .A2(n_29), .B1(n_844), .B2(n_845), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_17), .Y(n_845) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_18), .A2(n_48), .B(n_147), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_19), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_21), .B(n_133), .Y(n_561) );
INVx4_ASAP7_75t_R g224 ( .A(n_22), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_23), .B(n_136), .Y(n_161) );
OAI22x1_ASAP7_75t_SL g109 ( .A1(n_24), .A2(n_110), .B1(n_111), .B2(n_115), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_24), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_25), .A2(n_88), .B1(n_113), .B2(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_25), .Y(n_113) );
AO32x1_ASAP7_75t_L g515 ( .A1(n_26), .A2(n_144), .A3(n_145), .B1(n_516), .B2(n_519), .Y(n_515) );
AO32x2_ASAP7_75t_L g612 ( .A1(n_26), .A2(n_144), .A3(n_145), .B1(n_516), .B2(n_519), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_27), .B(n_133), .Y(n_170) );
INVx1_ASAP7_75t_L g188 ( .A(n_28), .Y(n_188) );
INVx1_ASAP7_75t_L g844 ( .A(n_29), .Y(n_844) );
A2O1A1Ixp33_ASAP7_75t_SL g266 ( .A1(n_30), .A2(n_135), .B(n_138), .C(n_267), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g137 ( .A1(n_31), .A2(n_45), .B1(n_138), .B2(n_139), .Y(n_137) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_32), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_33), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_34), .A2(n_51), .B1(n_133), .B2(n_225), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_35), .A2(n_93), .B1(n_131), .B2(n_139), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_36), .B(n_549), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_37), .B(n_570), .Y(n_590) );
INVx1_ASAP7_75t_L g167 ( .A(n_38), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_39), .B(n_138), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_40), .A2(n_68), .B1(n_139), .B2(n_524), .Y(n_523) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_41), .Y(n_247) );
INVx2_ASAP7_75t_L g813 ( .A(n_42), .Y(n_813) );
BUFx3_ASAP7_75t_L g816 ( .A(n_43), .Y(n_816) );
INVx1_ASAP7_75t_L g830 ( .A(n_43), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_44), .B(n_592), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_46), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_47), .A2(n_85), .B1(n_138), .B2(n_139), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_49), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_50), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_53), .A2(n_78), .B1(n_163), .B2(n_570), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_54), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_55), .A2(n_82), .B1(n_131), .B2(n_195), .Y(n_537) );
INVx1_ASAP7_75t_L g147 ( .A(n_56), .Y(n_147) );
AND2x4_ASAP7_75t_L g149 ( .A(n_57), .B(n_150), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_58), .A2(n_92), .B1(n_139), .B2(n_177), .Y(n_176) );
AO22x1_ASAP7_75t_L g193 ( .A1(n_59), .A2(n_73), .B1(n_162), .B2(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_60), .B(n_131), .Y(n_546) );
INVx1_ASAP7_75t_L g150 ( .A(n_61), .Y(n_150) );
AND2x2_ASAP7_75t_L g269 ( .A(n_62), .B(n_144), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_63), .B(n_144), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_64), .A2(n_105), .B1(n_863), .B2(n_875), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_65), .A2(n_837), .B(n_848), .Y(n_847) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_66), .A2(n_141), .B(n_198), .C(n_510), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_67), .B(n_131), .C(n_551), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_69), .B(n_198), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_70), .Y(n_262) );
AND2x2_ASAP7_75t_L g512 ( .A(n_71), .B(n_229), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_72), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_74), .B(n_133), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_75), .A2(n_99), .B1(n_163), .B2(n_195), .Y(n_572) );
INVx2_ASAP7_75t_L g136 ( .A(n_76), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_77), .B(n_249), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_79), .B(n_144), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_80), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_81), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_83), .B(n_154), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_84), .A2(n_108), .B1(n_109), .B2(n_116), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_84), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_87), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g114 ( .A(n_88), .Y(n_114) );
INVx1_ASAP7_75t_L g833 ( .A(n_89), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_89), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_90), .A2(n_103), .B1(n_139), .B2(n_225), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_91), .B(n_570), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_94), .B(n_144), .Y(n_244) );
INVx1_ASAP7_75t_L g489 ( .A(n_95), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_95), .B(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_96), .B(n_216), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g840 ( .A(n_97), .Y(n_840) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_98), .A2(n_184), .B(n_198), .C(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g228 ( .A(n_100), .B(n_229), .Y(n_228) );
NAND2xp33_ASAP7_75t_L g252 ( .A(n_101), .B(n_178), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_102), .Y(n_560) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_809), .B(n_819), .Y(n_105) );
XOR2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_117), .Y(n_106) );
INVx1_ASAP7_75t_L g116 ( .A(n_109), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_111), .Y(n_115) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_485), .B(n_490), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
XNOR2xp5_ASAP7_75t_L g842 ( .A(n_120), .B(n_843), .Y(n_842) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_362), .Y(n_120) );
NOR2x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_310), .Y(n_121) );
OAI211xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_189), .B(n_230), .C(n_295), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_125), .A2(n_231), .B(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_155), .Y(n_125) );
INVx2_ASAP7_75t_L g291 ( .A(n_126), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_126), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g402 ( .A(n_127), .B(n_157), .Y(n_402) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_SL g270 ( .A(n_128), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_128), .B(n_173), .Y(n_307) );
AND2x2_ASAP7_75t_L g340 ( .A(n_128), .B(n_257), .Y(n_340) );
OR2x2_ASAP7_75t_L g345 ( .A(n_128), .B(n_173), .Y(n_345) );
AO31x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_143), .A3(n_148), .B(n_151), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_134), .B1(n_137), .B2(n_140), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_131), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_SL g570 ( .A(n_131), .Y(n_570) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_132), .Y(n_133) );
INVx3_ASAP7_75t_L g138 ( .A(n_132), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_132), .Y(n_139) );
INVx1_ASAP7_75t_L g163 ( .A(n_132), .Y(n_163) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
INVx1_ASAP7_75t_L g182 ( .A(n_132), .Y(n_182) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
INVx1_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
INVx1_ASAP7_75t_L g200 ( .A(n_132), .Y(n_200) );
INVx1_ASAP7_75t_L g225 ( .A(n_132), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_133), .B(n_262), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_133), .A2(n_225), .B1(n_506), .B2(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g524 ( .A(n_133), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_134), .A2(n_176), .B1(n_179), .B2(n_183), .Y(n_175) );
OAI22x1_ASAP7_75t_L g205 ( .A1(n_134), .A2(n_183), .B1(n_206), .B2(n_208), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_134), .A2(n_140), .B1(n_523), .B2(n_525), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_134), .A2(n_135), .B1(n_537), .B2(n_538), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_134), .A2(n_569), .B1(n_571), .B2(n_572), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_134), .A2(n_590), .B(n_591), .Y(n_589) );
INVx6_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_135), .A2(n_193), .B(n_196), .C(n_202), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_135), .A2(n_252), .B(n_253), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_135), .B(n_193), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_135), .A2(n_265), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_135), .A2(n_546), .B(n_547), .Y(n_545) );
BUFx8_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
INVx1_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
INVx4_ASAP7_75t_L g207 ( .A(n_138), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_139), .B(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g180 ( .A(n_139), .Y(n_180) );
INVx2_ASAP7_75t_L g549 ( .A(n_139), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_140), .A2(n_169), .B(n_170), .Y(n_168) );
OAI21x1_ASAP7_75t_L g196 ( .A1(n_140), .A2(n_197), .B(n_201), .Y(n_196) );
AOI21x1_ASAP7_75t_L g586 ( .A1(n_140), .A2(n_587), .B(n_588), .Y(n_586) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g250 ( .A(n_142), .Y(n_250) );
AOI31xp67_ASAP7_75t_L g535 ( .A1(n_143), .A2(n_148), .A3(n_536), .B(n_539), .Y(n_535) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2x1_ASAP7_75t_L g254 ( .A(n_144), .B(n_255), .Y(n_254) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g171 ( .A(n_145), .B(n_148), .Y(n_171) );
BUFx3_ASAP7_75t_L g521 ( .A(n_145), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_145), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_145), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g557 ( .A(n_145), .Y(n_557) );
INVx2_ASAP7_75t_SL g584 ( .A(n_145), .Y(n_584) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
INVx1_ASAP7_75t_L g255 ( .A(n_148), .Y(n_255) );
OAI21x1_ASAP7_75t_L g544 ( .A1(n_148), .A2(n_545), .B(n_548), .Y(n_544) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_148), .A2(n_559), .B(n_562), .Y(n_558) );
BUFx10_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
INVx1_ASAP7_75t_L g203 ( .A(n_149), .Y(n_203) );
BUFx10_ASAP7_75t_L g210 ( .A(n_149), .Y(n_210) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_149), .A2(n_521), .A3(n_522), .B(n_526), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx2_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_153), .B(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_153), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g229 ( .A(n_153), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_153), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI21xp33_ASAP7_75t_L g202 ( .A1(n_154), .A2(n_201), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g209 ( .A(n_154), .Y(n_209) );
INVx2_ASAP7_75t_L g217 ( .A(n_154), .Y(n_217) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g484 ( .A(n_156), .Y(n_484) );
OR2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_172), .Y(n_156) );
AND2x2_ASAP7_75t_L g285 ( .A(n_157), .B(n_173), .Y(n_285) );
INVx3_ASAP7_75t_L g293 ( .A(n_157), .Y(n_293) );
NAND2x1p5_ASAP7_75t_SL g325 ( .A(n_157), .B(n_309), .Y(n_325) );
INVx1_ASAP7_75t_L g343 ( .A(n_157), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_157), .B(n_288), .Y(n_368) );
BUFx2_ASAP7_75t_L g454 ( .A(n_157), .Y(n_454) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_168), .B(n_171), .Y(n_159) );
OAI21xp33_ASAP7_75t_SL g160 ( .A1(n_161), .A2(n_162), .B(n_164), .Y(n_160) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_163), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
BUFx4f_ASAP7_75t_L g265 ( .A(n_166), .Y(n_265) );
INVx1_ASAP7_75t_L g551 ( .A(n_166), .Y(n_551) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g238 ( .A(n_173), .Y(n_238) );
INVx1_ASAP7_75t_L g294 ( .A(n_173), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_173), .B(n_270), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_173), .B(n_257), .Y(n_403) );
AO31x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .A3(n_185), .B(n_187), .Y(n_173) );
AOI21x1_ASAP7_75t_L g258 ( .A1(n_174), .A2(n_259), .B(n_269), .Y(n_258) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
OAI22xp33_ASAP7_75t_L g223 ( .A1(n_178), .A2(n_224), .B1(n_225), .B2(n_226), .Y(n_223) );
O2A1O1Ixp5_ASAP7_75t_L g559 ( .A1(n_181), .A2(n_265), .B(n_560), .C(n_561), .Y(n_559) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_182), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_183), .B(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g508 ( .A(n_184), .Y(n_508) );
INVx1_ASAP7_75t_SL g571 ( .A(n_184), .Y(n_571) );
AO31x2_ASAP7_75t_L g567 ( .A1(n_185), .A2(n_521), .A3(n_568), .B(n_573), .Y(n_567) );
INVx2_ASAP7_75t_SL g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_SL g519 ( .A(n_186), .Y(n_519) );
OR2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_213), .Y(n_189) );
INVx1_ASAP7_75t_L g461 ( .A(n_190), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_204), .Y(n_190) );
OR2x2_ASAP7_75t_L g233 ( .A(n_191), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g298 ( .A(n_191), .Y(n_298) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVxp67_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g592 ( .A(n_195), .Y(n_592) );
INVx1_ASAP7_75t_L g277 ( .A(n_196), .Y(n_277) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_200), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g279 ( .A(n_202), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_203), .A2(n_260), .B(n_266), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_203), .A2(n_504), .B(n_509), .Y(n_503) );
INVx2_ASAP7_75t_L g234 ( .A(n_204), .Y(n_234) );
OR2x2_ASAP7_75t_L g299 ( .A(n_204), .B(n_214), .Y(n_299) );
AND2x2_ASAP7_75t_L g304 ( .A(n_204), .B(n_214), .Y(n_304) );
INVx2_ASAP7_75t_L g349 ( .A(n_204), .Y(n_349) );
AND2x2_ASAP7_75t_L g390 ( .A(n_204), .B(n_243), .Y(n_390) );
AND2x2_ASAP7_75t_L g424 ( .A(n_204), .B(n_321), .Y(n_424) );
AO31x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_209), .A3(n_210), .B(n_211), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_207), .A2(n_247), .B(n_248), .C(n_249), .Y(n_246) );
INVx2_ASAP7_75t_L g543 ( .A(n_209), .Y(n_543) );
INVx2_ASAP7_75t_L g227 ( .A(n_210), .Y(n_227) );
INVx1_ASAP7_75t_L g235 ( .A(n_213), .Y(n_235) );
INVx1_ASAP7_75t_L g354 ( .A(n_213), .Y(n_354) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g274 ( .A(n_214), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g315 ( .A(n_214), .B(n_276), .Y(n_315) );
INVx2_ASAP7_75t_L g321 ( .A(n_214), .Y(n_321) );
AND2x2_ASAP7_75t_L g376 ( .A(n_214), .B(n_243), .Y(n_376) );
AND2x2_ASAP7_75t_L g433 ( .A(n_214), .B(n_242), .Y(n_433) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_218), .B(n_228), .Y(n_214) );
AOI21x1_ASAP7_75t_L g502 ( .A1(n_215), .A2(n_503), .B(n_512), .Y(n_502) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_222), .B(n_227), .Y(n_218) );
INVx1_ASAP7_75t_L g564 ( .A(n_225), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_236), .B1(n_271), .B2(n_282), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
NAND3xp33_ASAP7_75t_SL g411 ( .A(n_233), .B(n_412), .C(n_414), .Y(n_411) );
INVx1_ASAP7_75t_L g330 ( .A(n_234), .Y(n_330) );
AND2x2_ASAP7_75t_L g380 ( .A(n_234), .B(n_242), .Y(n_380) );
INVx1_ASAP7_75t_L g480 ( .A(n_235), .Y(n_480) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_237), .B(n_435), .Y(n_471) );
BUFx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g326 ( .A(n_238), .Y(n_326) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_256), .Y(n_240) );
INVx1_ASAP7_75t_L g314 ( .A(n_241), .Y(n_314) );
BUFx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g394 ( .A(n_242), .B(n_275), .Y(n_394) );
AND2x2_ASAP7_75t_L g413 ( .A(n_242), .B(n_320), .Y(n_413) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g281 ( .A(n_243), .Y(n_281) );
BUFx3_ASAP7_75t_L g319 ( .A(n_243), .Y(n_319) );
AND2x2_ASAP7_75t_L g348 ( .A(n_243), .B(n_349), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_251), .B(n_254), .Y(n_245) );
INVx2_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_250), .A2(n_563), .B1(n_564), .B2(n_565), .Y(n_562) );
INVx2_ASAP7_75t_L g441 ( .A(n_256), .Y(n_441) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_270), .Y(n_256) );
INVx2_ASAP7_75t_L g309 ( .A(n_257), .Y(n_309) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g288 ( .A(n_258), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B(n_265), .Y(n_260) );
INVx1_ASAP7_75t_L g289 ( .A(n_270), .Y(n_289) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x6_ASAP7_75t_L g272 ( .A(n_273), .B(n_280), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g328 ( .A(n_274), .B(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g458 ( .A(n_274), .Y(n_458) );
INVx1_ASAP7_75t_L g303 ( .A(n_275), .Y(n_303) );
AND2x2_ASAP7_75t_L g383 ( .A(n_275), .B(n_321), .Y(n_383) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g320 ( .A(n_276), .B(n_321), .Y(n_320) );
AOI21x1_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2x1_ASAP7_75t_L g332 ( .A(n_281), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g416 ( .A(n_281), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_290), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_283), .A2(n_324), .B1(n_327), .B2(n_331), .Y(n_323) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_284), .A2(n_304), .B1(n_336), .B2(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
BUFx2_ASAP7_75t_SL g322 ( .A(n_285), .Y(n_322) );
AND2x4_ASAP7_75t_L g440 ( .A(n_285), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g449 ( .A(n_285), .Y(n_449) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g361 ( .A(n_287), .Y(n_361) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_288), .B(n_293), .Y(n_419) );
INVxp67_ASAP7_75t_L g448 ( .A(n_288), .Y(n_448) );
AND2x2_ASAP7_75t_L g453 ( .A(n_288), .B(n_319), .Y(n_453) );
OR2x2_ASAP7_75t_L g435 ( .A(n_289), .B(n_309), .Y(n_435) );
INVx1_ASAP7_75t_L g316 ( .A(n_290), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_291), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g355 ( .A(n_292), .B(n_340), .Y(n_355) );
AND2x4_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_293), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g339 ( .A(n_293), .Y(n_339) );
OR2x2_ASAP7_75t_L g434 ( .A(n_293), .B(n_435), .Y(n_434) );
OAI21xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .B(n_305), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g358 ( .A(n_297), .Y(n_358) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g352 ( .A(n_298), .B(n_349), .Y(n_352) );
INVx2_ASAP7_75t_L g476 ( .A(n_298), .Y(n_476) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
AND2x2_ASAP7_75t_L g405 ( .A(n_302), .B(n_348), .Y(n_405) );
AND2x2_ASAP7_75t_L g430 ( .A(n_302), .B(n_376), .Y(n_430) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g333 ( .A(n_303), .Y(n_333) );
AND2x2_ASAP7_75t_L g360 ( .A(n_304), .B(n_314), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_304), .B(n_359), .Y(n_372) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g457 ( .A(n_307), .Y(n_457) );
OR2x2_ASAP7_75t_L g473 ( .A(n_307), .B(n_368), .Y(n_473) );
INVx1_ASAP7_75t_L g397 ( .A(n_309), .Y(n_397) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_334), .C(n_356), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_316), .B1(n_317), .B2(n_322), .C(n_323), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AND2x2_ASAP7_75t_L g336 ( .A(n_315), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_315), .B(n_380), .Y(n_464) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx3_ASAP7_75t_L g359 ( .A(n_319), .Y(n_359) );
AND3x1_ASAP7_75t_L g455 ( .A(n_319), .B(n_456), .C(n_457), .Y(n_455) );
AND2x2_ASAP7_75t_L g442 ( .A(n_320), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g452 ( .A(n_320), .Y(n_452) );
INVxp67_ASAP7_75t_L g466 ( .A(n_322), .Y(n_466) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
OR2x2_ASAP7_75t_L g421 ( .A(n_325), .B(n_345), .Y(n_421) );
INVx2_ASAP7_75t_L g456 ( .A(n_325), .Y(n_456) );
INVx1_ASAP7_75t_L g374 ( .A(n_326), .Y(n_374) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_328), .A2(n_376), .B(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_329), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g337 ( .A(n_330), .Y(n_337) );
OR2x2_ASAP7_75t_L g431 ( .A(n_330), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g391 ( .A(n_333), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_333), .B(n_390), .Y(n_470) );
AND3x1_ASAP7_75t_L g334 ( .A(n_335), .B(n_341), .C(n_346), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
AND2x2_ASAP7_75t_L g385 ( .A(n_337), .B(n_376), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_338), .A2(n_405), .B1(n_406), .B2(n_408), .Y(n_404) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
OAI321xp33_ASAP7_75t_L g427 ( .A1(n_339), .A2(n_428), .A3(n_429), .B1(n_431), .B2(n_434), .C(n_436), .Y(n_427) );
AND2x2_ASAP7_75t_L g479 ( .A(n_339), .B(n_344), .Y(n_479) );
AND2x2_ASAP7_75t_L g377 ( .A(n_340), .B(n_343), .Y(n_377) );
INVx2_ASAP7_75t_L g386 ( .A(n_342), .Y(n_386) );
AND2x2_ASAP7_75t_L g395 ( .A(n_342), .B(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g407 ( .A(n_345), .B(n_397), .Y(n_407) );
INVx2_ASAP7_75t_L g439 ( .A(n_345), .Y(n_439) );
OAI21xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_350), .B(n_355), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g443 ( .A(n_349), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_352), .B(n_359), .Y(n_369) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_361), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_359), .B(n_383), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_359), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g460 ( .A(n_359), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g428 ( .A(n_361), .Y(n_428) );
NOR2xp67_ASAP7_75t_L g362 ( .A(n_363), .B(n_425), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_387), .C(n_410), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_378), .Y(n_364) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_369), .B1(n_370), .B2(n_373), .C(n_375), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
OR2x2_ASAP7_75t_L g418 ( .A(n_367), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI21xp33_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_384), .B(n_386), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g415 ( .A(n_383), .B(n_416), .Y(n_415) );
OAI21xp33_ASAP7_75t_SL g398 ( .A1(n_384), .A2(n_399), .B(n_404), .Y(n_398) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_392), .B(n_395), .C(n_398), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_389), .B(n_464), .Y(n_463) );
NAND2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_397), .B(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_400), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_417), .B1(n_420), .B2(n_422), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_419), .Y(n_482) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_462), .C(n_477), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_444), .Y(n_426) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_440), .B(n_442), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_450), .C(n_459), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
AOI32xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .A3(n_454), .B1(n_455), .B2(n_458), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g478 ( .A(n_453), .B(n_479), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_465), .B(n_467), .Y(n_462) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI22x1_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B1(n_472), .B2(n_474), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_470), .A2(n_482), .B(n_483), .Y(n_481) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_480), .B(n_481), .Y(n_477) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx8_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx12f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_488), .Y(n_487) );
BUFx8_ASAP7_75t_SL g493 ( .A(n_488), .Y(n_493) );
AND2x2_ASAP7_75t_L g853 ( .A(n_488), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g870 ( .A(n_489), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_494), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
NAND4xp75_ASAP7_75t_L g494 ( .A(n_495), .B(n_683), .C(n_737), .D(n_781), .Y(n_494) );
NOR2x1_ASAP7_75t_L g495 ( .A(n_496), .B(n_636), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_602), .Y(n_496) );
O2A1O1Ixp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_528), .B(n_532), .C(n_575), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_513), .Y(n_498) );
AND2x2_ASAP7_75t_L g653 ( .A(n_499), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g642 ( .A(n_500), .B(n_578), .Y(n_642) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_501), .Y(n_608) );
AND2x2_ASAP7_75t_L g657 ( .A(n_501), .B(n_520), .Y(n_657) );
INVx1_ASAP7_75t_L g669 ( .A(n_501), .Y(n_669) );
INVx1_ASAP7_75t_L g767 ( .A(n_501), .Y(n_767) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g530 ( .A(n_502), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_505), .B(n_508), .Y(n_504) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g595 ( .A(n_514), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_520), .Y(n_514) );
AND2x2_ASAP7_75t_L g531 ( .A(n_515), .B(n_520), .Y(n_531) );
INVx1_ASAP7_75t_L g635 ( .A(n_515), .Y(n_635) );
INVx1_ASAP7_75t_L g746 ( .A(n_515), .Y(n_746) );
OAI21x1_ASAP7_75t_L g585 ( .A1(n_519), .A2(n_586), .B(n_589), .Y(n_585) );
INVx3_ASAP7_75t_L g578 ( .A(n_520), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_520), .B(n_582), .Y(n_633) );
AND2x2_ASAP7_75t_L g668 ( .A(n_520), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_L g708 ( .A(n_529), .Y(n_708) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g577 ( .A(n_530), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_530), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g610 ( .A(n_530), .Y(n_610) );
OR2x2_ASAP7_75t_L g674 ( .A(n_530), .B(n_582), .Y(n_674) );
OR2x2_ASAP7_75t_L g745 ( .A(n_530), .B(n_746), .Y(n_745) );
INVx2_ASAP7_75t_SL g682 ( .A(n_531), .Y(n_682) );
AND2x2_ASAP7_75t_L g734 ( .A(n_531), .B(n_597), .Y(n_734) );
AND2x2_ASAP7_75t_L g791 ( .A(n_531), .B(n_708), .Y(n_791) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_554), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_533), .B(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g800 ( .A(n_533), .B(n_801), .Y(n_800) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_542), .Y(n_533) );
INVx2_ASAP7_75t_L g601 ( .A(n_534), .Y(n_601) );
AND2x2_ASAP7_75t_L g626 ( .A(n_534), .B(n_605), .Y(n_626) );
AND2x2_ASAP7_75t_L g696 ( .A(n_534), .B(n_567), .Y(n_696) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g650 ( .A(n_535), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_540), .A2(n_541), .B1(n_832), .B2(n_834), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g604 ( .A(n_542), .B(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g665 ( .A(n_542), .B(n_556), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B(n_553), .Y(n_542) );
OAI21x1_ASAP7_75t_L g621 ( .A1(n_543), .A2(n_544), .B(n_553), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B(n_552), .Y(n_548) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g672 ( .A(n_555), .B(n_649), .Y(n_672) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_567), .Y(n_555) );
INVx2_ASAP7_75t_SL g594 ( .A(n_556), .Y(n_594) );
BUFx2_ASAP7_75t_L g647 ( .A(n_556), .Y(n_647) );
INVx1_ASAP7_75t_L g719 ( .A(n_556), .Y(n_719) );
AND2x2_ASAP7_75t_L g752 ( .A(n_556), .B(n_600), .Y(n_752) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_566), .Y(n_556) );
OA21x2_ASAP7_75t_L g605 ( .A1(n_557), .A2(n_558), .B(n_566), .Y(n_605) );
INVx2_ASAP7_75t_L g580 ( .A(n_567), .Y(n_580) );
INVx1_ASAP7_75t_L g600 ( .A(n_567), .Y(n_600) );
INVx1_ASAP7_75t_L g628 ( .A(n_567), .Y(n_628) );
AND2x2_ASAP7_75t_L g718 ( .A(n_567), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g759 ( .A(n_567), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g775 ( .A(n_567), .B(n_760), .Y(n_775) );
AND2x2_ASAP7_75t_L g801 ( .A(n_567), .B(n_605), .Y(n_801) );
OAI32xp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_579), .A3(n_594), .B1(n_595), .B2(n_598), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_577), .B(n_742), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_577), .B(n_780), .Y(n_779) );
AND2x4_ASAP7_75t_L g611 ( .A(n_578), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g713 ( .A(n_578), .Y(n_713) );
INVx1_ASAP7_75t_L g773 ( .A(n_578), .Y(n_773) );
INVx1_ASAP7_75t_L g711 ( .A(n_579), .Y(n_711) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx2_ASAP7_75t_SL g615 ( .A(n_580), .Y(n_615) );
AND2x2_ASAP7_75t_L g704 ( .A(n_580), .B(n_619), .Y(n_704) );
AND2x2_ASAP7_75t_L g772 ( .A(n_581), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx3_ASAP7_75t_L g597 ( .A(n_582), .Y(n_597) );
AND2x2_ASAP7_75t_L g607 ( .A(n_582), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g643 ( .A(n_582), .Y(n_643) );
AND2x2_ASAP7_75t_L g654 ( .A(n_582), .B(n_612), .Y(n_654) );
AND2x2_ASAP7_75t_L g678 ( .A(n_582), .B(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g688 ( .A(n_582), .B(n_679), .Y(n_688) );
INVxp67_ASAP7_75t_L g742 ( .A(n_582), .Y(n_742) );
BUFx2_ASAP7_75t_L g754 ( .A(n_582), .Y(n_754) );
INVx1_ASAP7_75t_L g758 ( .A(n_582), .Y(n_758) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_593), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_594), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g750 ( .A(n_594), .Y(n_750) );
AND2x2_ASAP7_75t_L g658 ( .A(n_597), .B(n_635), .Y(n_658) );
AND2x2_ASAP7_75t_L g787 ( .A(n_597), .B(n_611), .Y(n_787) );
OAI22xp5_ASAP7_75t_SL g675 ( .A1(n_598), .A2(n_676), .B1(n_680), .B2(n_681), .Y(n_675) );
O2A1O1Ixp5_ASAP7_75t_R g749 ( .A1(n_598), .A2(n_750), .B(n_751), .C(n_753), .Y(n_749) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g603 ( .A(n_599), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g617 ( .A(n_601), .Y(n_617) );
INVx1_ASAP7_75t_L g660 ( .A(n_601), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_601), .B(n_630), .Y(n_736) );
AND2x2_ASAP7_75t_L g748 ( .A(n_601), .B(n_619), .Y(n_748) );
AOI222xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_606), .B1(n_609), .B2(n_613), .C1(n_623), .C2(n_631), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_603), .A2(n_645), .B1(n_723), .B2(n_784), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_603), .A2(n_667), .B1(n_803), .B2(n_805), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_604), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_604), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g778 ( .A(n_604), .Y(n_778) );
INVx1_ASAP7_75t_L g808 ( .A(n_604), .Y(n_808) );
INVx1_ASAP7_75t_L g622 ( .A(n_605), .Y(n_622) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g677 ( .A(n_608), .Y(n_677) );
AOI321xp33_ASAP7_75t_L g755 ( .A1(n_609), .A2(n_653), .A3(n_756), .B1(n_761), .B2(n_762), .C(n_763), .Y(n_755) );
AND2x4_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
OR2x2_ASAP7_75t_L g687 ( .A(n_610), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g707 ( .A(n_611), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g679 ( .A(n_612), .Y(n_679) );
NAND2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
OR2x2_ASAP7_75t_L g680 ( .A(n_615), .B(n_649), .Y(n_680) );
AND2x2_ASAP7_75t_L g700 ( .A(n_615), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g790 ( .A(n_616), .Y(n_790) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx2_ASAP7_75t_L g721 ( .A(n_618), .Y(n_721) );
NAND2x1p5_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g630 ( .A(n_620), .Y(n_630) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g649 ( .A(n_621), .B(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_624), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVxp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_626), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g761 ( .A(n_630), .Y(n_761) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_632), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g694 ( .A(n_633), .Y(n_694) );
INVx1_ASAP7_75t_L g644 ( .A(n_634), .Y(n_644) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_635), .Y(n_692) );
INVx2_ASAP7_75t_L g726 ( .A(n_635), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_661), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_645), .B(n_651), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_640), .B(n_644), .Y(n_639) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g777 ( .A1(n_641), .A2(n_728), .B1(n_778), .B2(n_779), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx2_ASAP7_75t_L g743 ( .A(n_642), .Y(n_743) );
AND2x2_ASAP7_75t_L g667 ( .A(n_643), .B(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g681 ( .A(n_643), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g732 ( .A(n_643), .Y(n_732) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g712 ( .A(n_647), .B(n_648), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_647), .B(n_696), .Y(n_728) );
AND2x2_ASAP7_75t_L g774 ( .A(n_647), .B(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_648), .B(n_752), .Y(n_789) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g701 ( .A(n_649), .Y(n_701) );
INVx1_ASAP7_75t_L g760 ( .A(n_650), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_655), .B(n_659), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g722 ( .A(n_654), .B(n_677), .Y(n_722) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_657), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g731 ( .A(n_657), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_660), .B(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_675), .Y(n_661) );
OAI21xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B(n_670), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_663), .A2(n_730), .B1(n_733), .B2(n_735), .Y(n_729) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI311xp33_ASAP7_75t_L g763 ( .A1(n_665), .A2(n_764), .A3(n_765), .B(n_768), .C(n_769), .Y(n_763) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g691 ( .A(n_668), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_668), .B(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g762 ( .A(n_672), .Y(n_762) );
INVx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
INVx2_ASAP7_75t_L g768 ( .A(n_678), .Y(n_768) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_682), .Y(n_785) );
NOR2x1_ASAP7_75t_L g683 ( .A(n_684), .B(n_709), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_689), .C(n_697), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AO21x1_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_693), .B(n_695), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AO221x1_ASAP7_75t_L g770 ( .A1(n_691), .A2(n_771), .B1(n_774), .B2(n_776), .C(n_777), .Y(n_770) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g769 ( .A(n_696), .Y(n_769) );
OAI21xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_702), .B(n_705), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_713), .B(n_714), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g764 ( .A(n_713), .Y(n_764) );
AOI221x1_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_722), .B1(n_723), .B2(n_727), .C(n_729), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_720), .Y(n_715) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g747 ( .A(n_718), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AO22x1_ASAP7_75t_L g794 ( .A1(n_722), .A2(n_795), .B1(n_797), .B2(n_800), .Y(n_794) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g771 ( .A(n_725), .B(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_726), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVxp33_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_770), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_755), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_747), .B(n_749), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_744), .C(n_745), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g780 ( .A(n_742), .Y(n_780) );
AND2x2_ASAP7_75t_L g766 ( .A(n_746), .B(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g776 ( .A(n_752), .B(n_761), .Y(n_776) );
INVxp67_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NAND2x1p5_ASAP7_75t_L g804 ( .A(n_758), .B(n_766), .Y(n_804) );
INVx2_ASAP7_75t_L g796 ( .A(n_761), .Y(n_796) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g799 ( .A(n_767), .Y(n_799) );
AND2x2_ASAP7_75t_L g795 ( .A(n_775), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g807 ( .A(n_775), .Y(n_807) );
NOR2x1_ASAP7_75t_L g781 ( .A(n_782), .B(n_792), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_786), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_787), .A2(n_788), .B1(n_790), .B2(n_791), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_802), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OR2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx4_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AND2x6_ASAP7_75t_SL g811 ( .A(n_812), .B(n_814), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx3_ASAP7_75t_L g823 ( .A(n_813), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_813), .B(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_817), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NOR2x1_ASAP7_75t_L g854 ( .A(n_816), .B(n_818), .Y(n_854) );
NOR3x1_ASAP7_75t_L g866 ( .A(n_816), .B(n_867), .C(n_870), .Y(n_866) );
AND2x6_ASAP7_75t_SL g827 ( .A(n_817), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_855), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_841), .B(n_846), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .Y(n_821) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_822), .Y(n_862) );
BUFx3_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_831), .B(n_835), .Y(n_824) );
BUFx3_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx5_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx3_ASAP7_75t_L g839 ( .A(n_827), .Y(n_839) );
CKINVDCx8_ASAP7_75t_R g861 ( .A(n_827), .Y(n_861) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI21xp5_ASAP7_75t_SL g856 ( .A1(n_831), .A2(n_836), .B(n_857), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVxp67_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_840), .Y(n_837) );
BUFx2_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NAND3xp33_ASAP7_75t_L g855 ( .A(n_842), .B(n_856), .C(n_862), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_847), .Y(n_846) );
INVx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx6_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
BUFx10_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx6f_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx3_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx3_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx3_ASAP7_75t_SL g863 ( .A(n_864), .Y(n_863) );
INVx4_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
AND2x6_ASAP7_75t_L g865 ( .A(n_866), .B(n_871), .Y(n_865) );
AND2x6_ASAP7_75t_L g876 ( .A(n_866), .B(n_871), .Y(n_876) );
INVx2_ASAP7_75t_SL g867 ( .A(n_868), .Y(n_867) );
NOR2x1p5_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx3_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
endmodule