module fake_jpeg_6360_n_24 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_4),
.A2(n_2),
.B1(n_0),
.B2(n_6),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_2),
.B(n_0),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx12_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g14 ( 
.A(n_8),
.B(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_14),
.B(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_18),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_5),
.B1(n_13),
.B2(n_8),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_15),
.B1(n_12),
.B2(n_9),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_5),
.B(n_11),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_9),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_23),
.B1(n_9),
.B2(n_20),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_19),
.C(n_20),
.Y(n_23)
);


endmodule