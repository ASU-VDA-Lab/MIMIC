module fake_jpeg_3038_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_2),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

MAJIxp5_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_1),
.C(n_6),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_18),
.Y(n_26)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_0),
.B1(n_3),
.B2(n_14),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_15),
.B1(n_10),
.B2(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_0),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_17),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_15),
.B(n_13),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_20),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_23),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_38),
.Y(n_44)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_19),
.B(n_21),
.Y(n_37)
);

FAx1_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_41),
.CI(n_20),
.CON(n_42),
.SN(n_42)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_40),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_3),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_45),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_47),
.C(n_34),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_32),
.B(n_29),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_46),
.B(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_38),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_50),
.B(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_36),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_53),
.B(n_42),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_31),
.B(n_53),
.Y(n_55)
);


endmodule