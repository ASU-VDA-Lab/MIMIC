module fake_jpeg_3048_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_40),
.Y(n_67)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_53),
.B1(n_46),
.B2(n_48),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_68),
.B1(n_49),
.B2(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_60),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_41),
.B1(n_51),
.B2(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_57),
.Y(n_77)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_74),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_70),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_79),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_61),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_86),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_61),
.B1(n_45),
.B2(n_59),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_55),
.B(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_41),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_54),
.B1(n_42),
.B2(n_45),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_55),
.B1(n_50),
.B2(n_47),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_23),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_73),
.B1(n_72),
.B2(n_54),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_92),
.B1(n_101),
.B2(n_25),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_73),
.B1(n_45),
.B2(n_50),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_83),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_102),
.B1(n_105),
.B2(n_3),
.Y(n_113)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_83),
.B1(n_85),
.B2(n_5),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_77),
.B1(n_84),
.B2(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_47),
.B1(n_1),
.B2(n_2),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_112),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_30),
.C(n_28),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_120),
.C(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_4),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_6),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_118),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_102),
.B1(n_95),
.B2(n_105),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_121),
.B(n_123),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_24),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_122),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_21),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_134),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_106),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_129)
);

NOR4xp25_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_112),
.C(n_13),
.D(n_14),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_106),
.B(n_10),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_9),
.B(n_11),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_138),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_131),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_119),
.B1(n_124),
.B2(n_114),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_9),
.C(n_15),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_145),
.C(n_131),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_16),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_137),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_150),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_132),
.B1(n_125),
.B2(n_134),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_142),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_143),
.A2(n_135),
.B1(n_128),
.B2(n_133),
.Y(n_148)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_152),
.A2(n_153),
.B(n_146),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_151),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_150),
.B1(n_126),
.B2(n_152),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_127),
.CI(n_17),
.CON(n_157),
.SN(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_16),
.C(n_17),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_19),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_19),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_20),
.B1(n_157),
.B2(n_126),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_157),
.Y(n_162)
);


endmodule