module fake_jpeg_10743_n_503 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_6),
.B(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_51),
.B(n_61),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_8),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_33),
.B(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_14),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_8),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_85),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_84),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_7),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_90),
.Y(n_119)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_95),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_7),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_28),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_52),
.B(n_20),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_105),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_114),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_54),
.A2(n_21),
.B1(n_43),
.B2(n_44),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_147),
.B1(n_78),
.B2(n_76),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_61),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_38),
.B(n_37),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_154),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_62),
.A2(n_20),
.B1(n_43),
.B2(n_44),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_116),
.A2(n_41),
.B(n_47),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_49),
.A2(n_21),
.B1(n_20),
.B2(n_43),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_125),
.B1(n_81),
.B2(n_79),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_56),
.A2(n_21),
.B1(n_30),
.B2(n_45),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_85),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_130),
.B(n_24),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_38),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_145),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_93),
.A2(n_92),
.B1(n_88),
.B2(n_84),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_46),
.B1(n_34),
.B2(n_31),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_63),
.B(n_30),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_64),
.A2(n_74),
.B1(n_65),
.B2(n_72),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_42),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_42),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

HAxp5_ASAP7_75t_SL g154 ( 
.A(n_87),
.B(n_41),
.CON(n_154),
.SN(n_154)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_161),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_190),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_167),
.B(n_197),
.Y(n_249)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_147),
.B1(n_113),
.B2(n_133),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_98),
.B(n_45),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_171),
.B(n_177),
.Y(n_222)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_174),
.Y(n_263)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_176),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_34),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_178),
.A2(n_186),
.B1(n_187),
.B2(n_137),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_111),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_181),
.A2(n_185),
.B1(n_198),
.B2(n_201),
.Y(n_221)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_111),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_121),
.A2(n_46),
.B1(n_25),
.B2(n_31),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_125),
.A2(n_26),
.B1(n_25),
.B2(n_47),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_26),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_188),
.B(n_204),
.Y(n_230)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_109),
.Y(n_191)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_191),
.Y(n_256)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_192),
.Y(n_261)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_101),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_155),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_142),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_202),
.A2(n_208),
.B1(n_212),
.B2(n_137),
.Y(n_246)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_206),
.Y(n_251)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_207),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_102),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_209),
.B(n_210),
.Y(n_259)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_118),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_213),
.Y(n_231)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_140),
.B(n_9),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_148),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_214),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_157),
.B(n_41),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_219),
.B(n_10),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_225),
.A2(n_228),
.B1(n_245),
.B2(n_252),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_103),
.C(n_128),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_242),
.C(n_258),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_176),
.A2(n_156),
.B1(n_106),
.B2(n_143),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_227),
.A2(n_181),
.B1(n_185),
.B2(n_202),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_184),
.A2(n_141),
.B1(n_136),
.B2(n_133),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_160),
.B(n_143),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_244),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_164),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_165),
.B(n_127),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_127),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_162),
.B(n_190),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_162),
.B(n_106),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_257),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_170),
.A2(n_148),
.B1(n_129),
.B2(n_47),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_183),
.B(n_0),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_203),
.B(n_129),
.C(n_47),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_201),
.B(n_7),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_3),
.C(n_4),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_218),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_270),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_271),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_228),
.A2(n_179),
.B1(n_163),
.B2(n_159),
.Y(n_268)
);

OAI22x1_ASAP7_75t_L g310 ( 
.A1(n_268),
.A2(n_306),
.B1(n_254),
.B2(n_215),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_251),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_242),
.B(n_214),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_223),
.A2(n_175),
.B1(n_192),
.B2(n_173),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_273),
.A2(n_294),
.B1(n_216),
.B2(n_233),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_274),
.B(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_172),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_285),
.Y(n_320)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_279),
.Y(n_318)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_244),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_282),
.A2(n_283),
.B(n_290),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_182),
.B(n_207),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_212),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_198),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_292),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_219),
.B(n_199),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_289),
.C(n_258),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_226),
.A2(n_199),
.B(n_180),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_288),
.A2(n_303),
.B(n_235),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_222),
.B(n_174),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_221),
.A2(n_169),
.B(n_1),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_291),
.B(n_295),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_249),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_249),
.A2(n_166),
.B1(n_161),
.B2(n_0),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_296),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_237),
.B(n_3),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_298),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_259),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_224),
.B(n_3),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_301),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_224),
.B(n_16),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_235),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_249),
.A2(n_4),
.B(n_5),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_238),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_304),
.Y(n_333)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_236),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_308),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_250),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_236),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_289),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_234),
.C(n_241),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_327),
.Y(n_351)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_267),
.A2(n_230),
.A3(n_231),
.B1(n_245),
.B2(n_225),
.C1(n_252),
.C2(n_261),
.Y(n_321)
);

AOI21xp33_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_344),
.B(n_311),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_261),
.B(n_234),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_266),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_324),
.A2(n_331),
.B1(n_279),
.B2(n_284),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_307),
.A2(n_231),
.B1(n_230),
.B2(n_220),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_326),
.A2(n_291),
.B1(n_299),
.B2(n_296),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_253),
.C(n_243),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_271),
.B(n_243),
.C(n_239),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_337),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_269),
.A2(n_273),
.B1(n_294),
.B2(n_302),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_300),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_336),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_301),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_271),
.B(n_239),
.C(n_263),
.Y(n_337)
);

OA22x2_ASAP7_75t_L g338 ( 
.A1(n_282),
.A2(n_250),
.B1(n_215),
.B2(n_263),
.Y(n_338)
);

AOI22x1_ASAP7_75t_L g379 ( 
.A1(n_338),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_267),
.B(n_248),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_340),
.B(n_304),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_271),
.B(n_233),
.C(n_216),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_287),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_276),
.A2(n_216),
.B1(n_254),
.B2(n_248),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_342),
.A2(n_346),
.B1(n_302),
.B2(n_277),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_265),
.A2(n_232),
.B1(n_9),
.B2(n_11),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_264),
.A2(n_232),
.B1(n_11),
.B2(n_13),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_347),
.Y(n_358)
);

AO22x1_ASAP7_75t_L g348 ( 
.A1(n_292),
.A2(n_5),
.B1(n_11),
.B2(n_13),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_348),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_350),
.A2(n_371),
.B1(n_378),
.B2(n_379),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_339),
.A2(n_290),
.B(n_288),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_353),
.A2(n_356),
.B(n_361),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_366),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_355),
.B(n_368),
.C(n_319),
.Y(n_395)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_334),
.Y(n_359)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_359),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_313),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_360),
.B(n_364),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_339),
.A2(n_283),
.B(n_292),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_362),
.B(n_319),
.Y(n_400)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_363),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_313),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_320),
.A2(n_265),
.B1(n_272),
.B2(n_285),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_365),
.A2(n_367),
.B1(n_369),
.B2(n_375),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_297),
.C(n_303),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_309),
.B(n_272),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_320),
.A2(n_286),
.B1(n_270),
.B2(n_298),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_275),
.Y(n_370)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_293),
.Y(n_373)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_373),
.Y(n_403)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_312),
.Y(n_374)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_374),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_328),
.A2(n_295),
.B1(n_281),
.B2(n_279),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_313),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_376),
.Y(n_397)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_312),
.Y(n_377)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_322),
.A2(n_305),
.B1(n_308),
.B2(n_14),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_325),
.B(n_15),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_380),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_328),
.A2(n_15),
.B1(n_16),
.B2(n_344),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_381),
.A2(n_333),
.B1(n_329),
.B2(n_343),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_355),
.B(n_314),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_387),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_368),
.B(n_327),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_356),
.A2(n_311),
.B1(n_324),
.B2(n_322),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_389),
.A2(n_370),
.B1(n_349),
.B2(n_365),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_352),
.A2(n_317),
.B1(n_333),
.B2(n_346),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_316),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_396),
.C(n_399),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_351),
.B(n_330),
.C(n_337),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_352),
.A2(n_342),
.B1(n_329),
.B2(n_343),
.Y(n_398)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_398),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_311),
.C(n_341),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_406),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_349),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_338),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_362),
.B(n_345),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_357),
.B(n_345),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_409),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_367),
.A2(n_369),
.B1(n_381),
.B2(n_375),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_408),
.A2(n_386),
.B1(n_383),
.B2(n_403),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_357),
.B(n_335),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_410),
.A2(n_422),
.B1(n_408),
.B2(n_397),
.Y(n_437)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_412),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_394),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_416),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_372),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g444 ( 
.A(n_415),
.Y(n_444)
);

FAx1_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_353),
.CI(n_361),
.CON(n_417),
.SN(n_417)
);

AOI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_417),
.A2(n_406),
.B(n_409),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_391),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_419),
.B(n_429),
.Y(n_439)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_392),
.Y(n_420)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_420),
.Y(n_450)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_424),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_383),
.A2(n_363),
.B1(n_373),
.B2(n_358),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_402),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_433),
.B1(n_385),
.B2(n_404),
.Y(n_434)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_402),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_428),
.Y(n_436)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_382),
.B(n_380),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_382),
.B(n_371),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_430),
.B(n_432),
.Y(n_438)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_405),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_386),
.A2(n_378),
.B1(n_310),
.B2(n_379),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_434),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_437),
.A2(n_442),
.B1(n_443),
.B2(n_447),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_396),
.C(n_384),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_448),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_423),
.A2(n_393),
.B1(n_399),
.B2(n_401),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_410),
.A2(n_393),
.B1(n_379),
.B2(n_388),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_445),
.B(n_449),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_423),
.A2(n_407),
.B(n_395),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_446),
.A2(n_452),
.B(n_411),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_418),
.A2(n_335),
.B1(n_338),
.B2(n_318),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_387),
.C(n_400),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_338),
.C(n_323),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_424),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_412),
.A2(n_323),
.B(n_348),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_418),
.A2(n_318),
.B1(n_348),
.B2(n_15),
.Y(n_453)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_453),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_431),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_466),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_448),
.B(n_411),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_455),
.B(n_457),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_446),
.C(n_426),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_458),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_460),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_425),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_462),
.B(n_451),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_434),
.A2(n_414),
.B1(n_415),
.B2(n_417),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_464),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_451),
.A2(n_417),
.B1(n_433),
.B2(n_432),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_465),
.B(n_468),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_426),
.Y(n_468)
);

XOR2x2_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_435),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_465),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_459),
.A2(n_445),
.B(n_444),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_474),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_461),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_473),
.B(n_476),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_439),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_437),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_478),
.A2(n_464),
.B1(n_443),
.B2(n_460),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_456),
.C(n_457),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_487),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_484),
.A2(n_488),
.B(n_470),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_480),
.A2(n_467),
.B1(n_435),
.B2(n_438),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_485),
.B(n_486),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_468),
.Y(n_486)
);

O2A1O1Ixp33_ASAP7_75t_SL g487 ( 
.A1(n_480),
.A2(n_440),
.B(n_450),
.C(n_438),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_483),
.B(n_475),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_486),
.C(n_475),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_491),
.B(n_493),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_481),
.A2(n_479),
.B(n_477),
.Y(n_493)
);

NAND4xp25_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_490),
.C(n_469),
.D(n_484),
.Y(n_498)
);

OAI321xp33_ASAP7_75t_L g496 ( 
.A1(n_490),
.A2(n_487),
.A3(n_436),
.B1(n_428),
.B2(n_492),
.C(n_482),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_496),
.A2(n_436),
.B1(n_494),
.B2(n_450),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_497),
.B(n_498),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_499),
.A2(n_427),
.B(n_470),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_452),
.B(n_447),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_501),
.B(n_453),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_455),
.B(n_16),
.Y(n_503)
);


endmodule