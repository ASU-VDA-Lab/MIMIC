module fake_jpeg_27662_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_0),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_47),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_60),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_59),
.B(n_21),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_26),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_24),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_73),
.Y(n_122)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_70),
.Y(n_102)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_75),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_33),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_82),
.Y(n_107)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_78),
.B(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_26),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_86),
.Y(n_104)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_17),
.B1(n_32),
.B2(n_33),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_92),
.B1(n_93),
.B2(n_28),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_32),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_31),
.Y(n_86)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_31),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_35),
.B1(n_40),
.B2(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_58),
.B1(n_61),
.B2(n_57),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_17),
.B1(n_32),
.B2(n_35),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_17),
.B1(n_28),
.B2(n_16),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_44),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_17),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_18),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_27),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_28),
.B1(n_39),
.B2(n_40),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_101),
.B(n_100),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_116),
.B1(n_121),
.B2(n_69),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_18),
.B1(n_34),
.B2(n_31),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_89),
.B1(n_94),
.B2(n_70),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_18),
.Y(n_115)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_88),
.A2(n_25),
.B1(n_22),
.B2(n_16),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_71),
.A2(n_25),
.B1(n_22),
.B2(n_16),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

BUFx2_ASAP7_75t_SL g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_27),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_96),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_79),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_71),
.Y(n_136)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_136),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_141),
.Y(n_181)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_139),
.B(n_147),
.Y(n_187)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_100),
.B1(n_67),
.B2(n_73),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_152),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_73),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_86),
.B1(n_69),
.B2(n_74),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_159),
.B1(n_112),
.B2(n_128),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_154),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_106),
.B(n_129),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_155),
.B(n_122),
.Y(n_165)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_69),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_85),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_110),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_95),
.Y(n_157)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_114),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_133),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_141),
.B(n_137),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_166),
.Y(n_214)
);

OAI22x1_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_125),
.B1(n_101),
.B2(n_106),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_170),
.B1(n_171),
.B2(n_182),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_180),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_125),
.B1(n_105),
.B2(n_111),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_172),
.Y(n_220)
);

AO22x1_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_121),
.B1(n_116),
.B2(n_100),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_141),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_110),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_194),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_144),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_105),
.B1(n_111),
.B2(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_184),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_141),
.B1(n_137),
.B2(n_145),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_185),
.A2(n_191),
.B1(n_82),
.B2(n_85),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_189),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_127),
.B1(n_124),
.B2(n_77),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_132),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_123),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_136),
.B(n_21),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_195),
.A2(n_201),
.B(n_212),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_196),
.B(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_204),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_158),
.B(n_142),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_20),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_1),
.C(n_2),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_205),
.B(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_178),
.C(n_163),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_211),
.C(n_170),
.Y(n_232)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_187),
.B(n_25),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_210),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_140),
.C(n_138),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_167),
.A2(n_137),
.B(n_57),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_181),
.A2(n_51),
.B(n_72),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_216),
.B(n_224),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_51),
.B(n_124),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_162),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_219),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_171),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_31),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_85),
.B(n_87),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_SL g225 ( 
.A(n_173),
.B(n_20),
.Y(n_225)
);

AOI32xp33_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_30),
.A3(n_27),
.B1(n_23),
.B2(n_164),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_230),
.B(n_234),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_216),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_195),
.A2(n_186),
.B1(n_185),
.B2(n_174),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_233),
.A2(n_206),
.B1(n_197),
.B2(n_29),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_207),
.B(n_20),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_175),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_241),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_202),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_175),
.C(n_164),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_246),
.C(n_223),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_30),
.C(n_27),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_30),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_247),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_214),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_214),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_262),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_256),
.C(n_242),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_218),
.C(n_200),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_258),
.C(n_263),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_R g257 ( 
.A(n_240),
.B(n_220),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_270),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_234),
.C(n_230),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_238),
.A2(n_208),
.B1(n_204),
.B2(n_224),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_233),
.B1(n_238),
.B2(n_231),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_212),
.B(n_203),
.C(n_213),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_198),
.C(n_197),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_266),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_269),
.A2(n_227),
.B1(n_236),
.B2(n_235),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_237),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_29),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_275),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_282),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_259),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_271),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_228),
.C(n_236),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_285),
.C(n_286),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_248),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_228),
.B1(n_248),
.B2(n_226),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_239),
.C(n_229),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_226),
.C(n_229),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_250),
.C(n_30),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_252),
.C(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_283),
.A2(n_264),
.B1(n_261),
.B2(n_267),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_293),
.A2(n_303),
.B1(n_4),
.B2(n_5),
.Y(n_313)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_4),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_272),
.A2(n_266),
.B(n_265),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_293),
.B(n_304),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_2),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_301),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_23),
.C(n_29),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_299),
.C(n_298),
.Y(n_307)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_276),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_279),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_288),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_286),
.A2(n_22),
.B1(n_23),
.B2(n_6),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_291),
.B(n_287),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_277),
.B1(n_278),
.B2(n_289),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_312),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_292),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_297),
.A2(n_278),
.B1(n_23),
.B2(n_6),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_314),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_291),
.A2(n_300),
.B1(n_295),
.B2(n_290),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_292),
.C(n_9),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_303),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_10),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_320),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_307),
.C(n_312),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_8),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_316),
.Y(n_326)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_324),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_322),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_325),
.B(n_323),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_317),
.C(n_313),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_329),
.A2(n_321),
.B(n_305),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_333),
.A3(n_330),
.B1(n_328),
.B2(n_14),
.C1(n_11),
.C2(n_13),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_12),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_12),
.B(n_13),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_15),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_340)
);


endmodule