module real_jpeg_24361_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_179;
wire n_167;
wire n_244;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_3),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_3),
.A2(n_28),
.B1(n_52),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_28),
.B1(n_33),
.B2(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_3),
.A2(n_28),
.B1(n_58),
.B2(n_60),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_54),
.B(n_161),
.C(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_3),
.B(n_57),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_60),
.B(n_78),
.C(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_3),
.B(n_22),
.C(n_36),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_3),
.B(n_76),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_3),
.B(n_119),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_3),
.B(n_38),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_4),
.A2(n_33),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_4),
.A2(n_43),
.B1(n_58),
.B2(n_60),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_43),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_4),
.A2(n_43),
.B1(n_51),
.B2(n_55),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_51),
.B1(n_52),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_8),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_58),
.B1(n_60),
.B2(n_104),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_8),
.A2(n_33),
.B1(n_37),
.B2(n_104),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_8),
.A2(n_22),
.B1(n_27),
.B2(n_104),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_10),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_10),
.A2(n_40),
.B1(n_58),
.B2(n_60),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_10),
.A2(n_22),
.B1(n_27),
.B2(n_40),
.Y(n_115)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_11),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_11),
.B(n_216),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_130),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_128),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_105),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_15),
.B(n_105),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_85),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_65),
.B2(n_66),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_20),
.A2(n_29),
.B1(n_45),
.B2(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_20),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_20),
.A2(n_45),
.B1(n_186),
.B2(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_26),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_21),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_21),
.B(n_26),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_21),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_22),
.B(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_24),
.Y(n_165)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_28),
.A2(n_53),
.B(n_60),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_28),
.A2(n_37),
.B(n_79),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_29),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_39),
.B(n_41),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_30),
.A2(n_69),
.B(n_71),
.Y(n_142)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_31),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_31),
.B(n_70),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_31),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_33),
.A2(n_37),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_33),
.B(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_38),
.B(n_191),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_39),
.A2(n_71),
.B(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_41),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_41),
.B(n_190),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_61),
.B(n_62),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_49),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_49),
.B(n_63),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_57),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_52),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_63),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_57),
.B(n_127),
.Y(n_156)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_60),
.B1(n_78),
.B2(n_79),
.Y(n_82)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_74),
.B(n_84),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_68),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_73),
.B(n_201),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_80),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_76),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_83),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_81),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_77),
.B(n_123),
.Y(n_154)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_80),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_81),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.C(n_99),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_87),
.B(n_92),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_88),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_90),
.A2(n_115),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_90),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_99),
.B1(n_100),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_152),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_96),
.B(n_145),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.C(n_111),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_106),
.B(n_109),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_111),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_122),
.C(n_124),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_112),
.A2(n_113),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_120),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_120),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_117),
.B(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_121),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_122),
.A2(n_124),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_122),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_124),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_266),
.B(n_270),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_179),
.B(n_252),
.C(n_265),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_167),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_133),
.B(n_167),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_149),
.B2(n_166),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_147),
.B2(n_148),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_136),
.B(n_148),
.C(n_166),
.Y(n_253)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_139),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_159),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_150)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_151),
.B(n_158),
.C(n_159),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_155),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_164),
.Y(n_173)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.C(n_174),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_168),
.A2(n_169),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_174),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.C(n_177),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_251),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_195),
.B(n_250),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_192),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_182),
.B(n_192),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_188),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_183),
.B(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_185),
.B(n_188),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_186),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_245),
.B(n_249),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_236),
.B(n_244),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_218),
.B(n_235),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_199),
.B(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_202),
.B1(n_203),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_212),
.B2(n_217),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_208),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_211),
.C(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_224),
.B(n_234),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_230),
.B(n_233),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_231),
.B(n_232),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_237),
.B(n_238),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_254),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_264),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_262),
.B2(n_263),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_263),
.C(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);


endmodule