module fake_jpeg_28652_n_518 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_518);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_518;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_61),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_20),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_64),
.Y(n_105)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_20),
.B(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_17),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_71),
.B(n_74),
.Y(n_156)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_17),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_80),
.B(n_82),
.Y(n_157)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_10),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_90),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_24),
.B(n_10),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_96),
.Y(n_118)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_29),
.B(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_44),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_94),
.B(n_102),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_37),
.B(n_8),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_36),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_37),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_125),
.B(n_144),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_131),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_90),
.A2(n_28),
.B1(n_49),
.B2(n_40),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_139),
.A2(n_38),
.B1(n_24),
.B2(n_33),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_58),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_145),
.Y(n_178)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_142),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_66),
.A2(n_28),
.B1(n_43),
.B2(n_47),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_61),
.B1(n_78),
.B2(n_95),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_68),
.B(n_40),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_63),
.Y(n_145)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

AND2x4_ASAP7_75t_SL g159 ( 
.A(n_100),
.B(n_43),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_98),
.Y(n_188)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_55),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_57),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_38),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_166),
.B(n_197),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_167),
.Y(n_252)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx4_ASAP7_75t_SL g235 ( 
.A(n_168),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_72),
.B1(n_92),
.B2(n_93),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_187),
.B1(n_194),
.B2(n_199),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_170),
.A2(n_202),
.B1(n_207),
.B2(n_131),
.Y(n_226)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_173),
.Y(n_249)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_175),
.Y(n_251)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_147),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_181),
.B(n_200),
.Y(n_241)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

NAND2x1_ASAP7_75t_SL g186 ( 
.A(n_113),
.B(n_43),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_141),
.A2(n_28),
.B1(n_45),
.B2(n_48),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_45),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_196),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_103),
.B1(n_97),
.B2(n_59),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_48),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_52),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_43),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_201),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_156),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_113),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_137),
.A2(n_65),
.B1(n_60),
.B2(n_76),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_105),
.B(n_52),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_208),
.Y(n_248)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_124),
.A2(n_84),
.B1(n_57),
.B2(n_43),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_206),
.A2(n_134),
.B1(n_107),
.B2(n_108),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_128),
.A2(n_73),
.B1(n_87),
.B2(n_91),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_105),
.B(n_33),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_154),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_211),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_152),
.A2(n_39),
.B1(n_47),
.B2(n_35),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_215),
.B1(n_130),
.B2(n_162),
.Y(n_243)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

CKINVDCx12_ASAP7_75t_R g214 ( 
.A(n_104),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_214),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_129),
.A2(n_150),
.B1(n_162),
.B2(n_136),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_221),
.B(n_227),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_155),
.B1(n_138),
.B2(n_132),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_219),
.A2(n_179),
.B1(n_183),
.B2(n_195),
.Y(n_273)
);

OAI22x1_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_159),
.B1(n_143),
.B2(n_104),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_158),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_223),
.B(n_229),
.C(n_254),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_107),
.B(n_134),
.C(n_25),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_225),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_219),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_117),
.C(n_120),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_220),
.B1(n_136),
.B2(n_150),
.Y(n_264)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

AOI21xp33_ASAP7_75t_L g247 ( 
.A1(n_197),
.A2(n_32),
.B(n_31),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_247),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_172),
.Y(n_250)
);

INVx11_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_18),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_267),
.B1(n_269),
.B2(n_275),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_241),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_285),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_208),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_261),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_186),
.Y(n_261)
);

BUFx24_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

CKINVDCx10_ASAP7_75t_R g263 ( 
.A(n_235),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_264),
.A2(n_273),
.B1(n_280),
.B2(n_250),
.Y(n_305)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_226),
.A2(n_202),
.B1(n_199),
.B2(n_207),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_200),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_224),
.B(n_218),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_181),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_276),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_189),
.B1(n_179),
.B2(n_132),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_217),
.B(n_178),
.Y(n_276)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_278),
.Y(n_320)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_235),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_203),
.B1(n_165),
.B2(n_180),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_239),
.A2(n_123),
.B1(n_210),
.B2(n_173),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_283),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_229),
.A2(n_123),
.B1(n_165),
.B2(n_177),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_287),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_218),
.B(n_183),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_253),
.A2(n_168),
.B1(n_174),
.B2(n_110),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_286),
.A2(n_290),
.B(n_182),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_184),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_225),
.B(n_209),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_288),
.B(n_283),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_289),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_253),
.A2(n_174),
.B1(n_213),
.B2(n_171),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_228),
.B(n_205),
.C(n_195),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_234),
.C(n_237),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_293),
.B(n_307),
.C(n_309),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_312),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_245),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_319),
.Y(n_338)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_277),
.A2(n_228),
.B(n_233),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_314),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_305),
.A2(n_322),
.B1(n_282),
.B2(n_263),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_277),
.A2(n_250),
.B1(n_238),
.B2(n_246),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_306),
.A2(n_313),
.B1(n_321),
.B2(n_323),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_260),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_233),
.C(n_242),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_288),
.A2(n_238),
.B(n_182),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_310),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_242),
.C(n_244),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_262),
.A2(n_238),
.B1(n_167),
.B2(n_222),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_261),
.A2(n_244),
.B(n_230),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_270),
.B(n_163),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_291),
.Y(n_328)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_281),
.A2(n_287),
.A3(n_288),
.B1(n_262),
.B2(n_267),
.Y(n_316)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_257),
.Y(n_317)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_272),
.B(n_234),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_262),
.A2(n_249),
.B1(n_108),
.B2(n_127),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_269),
.A2(n_127),
.B1(n_240),
.B2(n_255),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_289),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_348),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_327),
.A2(n_351),
.B1(n_353),
.B2(n_324),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_315),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_292),
.B(n_276),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_329),
.B(n_331),
.Y(n_358)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_330),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_292),
.B(n_285),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_269),
.B1(n_258),
.B2(n_273),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_333),
.A2(n_337),
.B1(n_346),
.B2(n_340),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_302),
.B(n_270),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_334),
.B(n_335),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_302),
.B(n_265),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_296),
.A2(n_258),
.B1(n_280),
.B2(n_265),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_300),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_339),
.B(n_343),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_251),
.Y(n_343)
);

AND2x6_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_279),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_357),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_296),
.A2(n_278),
.B1(n_268),
.B2(n_289),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_298),
.B(n_266),
.Y(n_350)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_301),
.A2(n_305),
.B1(n_313),
.B2(n_306),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_295),
.B(n_274),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_352),
.B(n_323),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_316),
.A2(n_274),
.B1(n_251),
.B2(n_236),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_255),
.Y(n_354)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_303),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_356),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_294),
.B(n_31),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_317),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_307),
.C(n_309),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_368),
.C(n_374),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_329),
.A2(n_324),
.B1(n_304),
.B2(n_314),
.Y(n_360)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_372),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_362),
.A2(n_332),
.B1(n_326),
.B2(n_25),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_335),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_364),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_353),
.A2(n_310),
.B1(n_312),
.B2(n_293),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_365),
.A2(n_366),
.B1(n_47),
.B2(n_41),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_318),
.B1(n_322),
.B2(n_321),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_337),
.A2(n_311),
.B1(n_299),
.B2(n_320),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_367),
.B(n_381),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_299),
.C(n_297),
.Y(n_368)
);

NOR3xp33_ASAP7_75t_SL g369 ( 
.A(n_338),
.B(n_318),
.C(n_297),
.Y(n_369)
);

NOR3xp33_ASAP7_75t_SL g414 ( 
.A(n_369),
.B(n_375),
.C(n_382),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_164),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_357),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_338),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_377),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_175),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_126),
.C(n_119),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_331),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_379),
.A2(n_384),
.B1(n_351),
.B2(n_341),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_333),
.A2(n_236),
.B1(n_25),
.B2(n_27),
.Y(n_381)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_348),
.A2(n_35),
.B(n_27),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_386),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_383),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_336),
.A2(n_34),
.B1(n_27),
.B2(n_31),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_334),
.B(n_32),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_376),
.A2(n_352),
.B(n_344),
.Y(n_391)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_391),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_359),
.B(n_342),
.C(n_350),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_400),
.C(n_407),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_395),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_394),
.A2(n_399),
.B1(n_408),
.B2(n_412),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_358),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_378),
.A2(n_341),
.B1(n_356),
.B2(n_340),
.Y(n_396)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_361),
.B(n_354),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_398),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_379),
.A2(n_346),
.B1(n_347),
.B2(n_355),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_347),
.C(n_332),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_406),
.A2(n_413),
.B1(n_381),
.B2(n_380),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_326),
.C(n_116),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_367),
.A2(n_176),
.B1(n_41),
.B2(n_47),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_387),
.Y(n_409)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_409),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_171),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_411),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_365),
.B(n_171),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_414),
.A2(n_380),
.B1(n_35),
.B2(n_34),
.Y(n_432)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_375),
.Y(n_416)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_416),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_401),
.A2(n_373),
.B(n_382),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_417),
.A2(n_7),
.B(n_14),
.Y(n_456)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_402),
.Y(n_423)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_423),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_389),
.B(n_388),
.C(n_385),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_424),
.B(n_429),
.Y(n_445)
);

AOI21xp33_ASAP7_75t_L g426 ( 
.A1(n_405),
.A2(n_385),
.B(n_388),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_426),
.A2(n_8),
.B(n_15),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_390),
.B(n_374),
.C(n_362),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_433),
.C(n_407),
.Y(n_448)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_406),
.Y(n_429)
);

FAx1_ASAP7_75t_SL g430 ( 
.A(n_397),
.B(n_366),
.CI(n_384),
.CON(n_430),
.SN(n_430)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_432),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_434),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_41),
.C(n_171),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_399),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_7),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_413),
.A2(n_394),
.B1(n_414),
.B2(n_411),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_438),
.A2(n_439),
.B1(n_84),
.B2(n_34),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_418),
.B(n_415),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_453),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_428),
.A2(n_393),
.B(n_412),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_442),
.A2(n_455),
.B(n_456),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_437),
.B(n_403),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_450),
.Y(n_467)
);

MAJx2_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_392),
.C(n_400),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_447),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_403),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_452),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_427),
.B(n_398),
.C(n_410),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_437),
.C(n_433),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_L g450 ( 
.A1(n_428),
.A2(n_412),
.B(n_408),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_421),
.B(n_32),
.Y(n_453)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_454),
.Y(n_459)
);

XOR2x1_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_7),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_14),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_436),
.A2(n_7),
.B(n_14),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_458),
.B(n_14),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_462),
.B(n_469),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_419),
.C(n_438),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_443),
.C(n_422),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_421),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_468),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_429),
.Y(n_469)
);

INVx11_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_470),
.B(n_474),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_422),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_4),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_472),
.B(n_473),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_451),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_420),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_447),
.B(n_431),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_475),
.B(n_462),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_461),
.Y(n_477)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_463),
.A2(n_449),
.B(n_417),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_478),
.A2(n_488),
.B(n_460),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_483),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_470),
.A2(n_439),
.B(n_455),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_480),
.A2(n_467),
.B(n_464),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_452),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_489),
.C(n_464),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_461),
.A2(n_450),
.B1(n_456),
.B2(n_430),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_484),
.B(n_471),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_486),
.B(n_459),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_463),
.A2(n_4),
.B(n_13),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_0),
.C(n_1),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_491),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_494),
.Y(n_503)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_496),
.B(n_497),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_485),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_495),
.B(n_499),
.C(n_486),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_4),
.C(n_12),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_489),
.B(n_3),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_0),
.C(n_1),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_504),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_498),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_12),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_500),
.A2(n_480),
.B1(n_487),
.B2(n_483),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_495),
.A2(n_481),
.B1(n_3),
.B2(n_11),
.Y(n_506)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_506),
.Y(n_510)
);

A2O1A1Ixp33_ASAP7_75t_L g509 ( 
.A1(n_503),
.A2(n_496),
.B(n_499),
.C(n_3),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_509),
.B(n_511),
.C(n_507),
.Y(n_513)
);

BUFx24_ASAP7_75t_SL g512 ( 
.A(n_508),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_513),
.B(n_505),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_510),
.B1(n_502),
.B2(n_16),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_0),
.B(n_2),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_516),
.B(n_2),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_517),
.A2(n_2),
.B(n_428),
.Y(n_518)
);


endmodule