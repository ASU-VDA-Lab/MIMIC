module fake_jpeg_19481_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

INVx4_ASAP7_75t_SL g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_3),
.B(n_2),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_12),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_7),
.A2(n_0),
.B1(n_3),
.B2(n_6),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_0),
.B(n_7),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_6),
.C(n_8),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_13),
.C(n_11),
.Y(n_33)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_29),
.B(n_23),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_11),
.B1(n_25),
.B2(n_13),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_14),
.B(n_19),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_13),
.C(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_7),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_28),
.B(n_27),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_39),
.C(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_37),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_41),
.B(n_36),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_32),
.C(n_11),
.Y(n_43)
);


endmodule