module real_jpeg_15672_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_286;
wire n_288;
wire n_292;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_258;
wire n_110;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_295;
wire n_167;
wire n_213;
wire n_179;
wire n_133;
wire n_202;
wire n_216;
wire n_138;
wire n_257;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

AND2x4_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_0),
.B(n_61),
.Y(n_60)
);

AND2x4_ASAP7_75t_SL g72 ( 
.A(n_0),
.B(n_73),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_0),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_0),
.B(n_55),
.Y(n_116)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_0),
.Y(n_139)
);

NAND2x1p5_ASAP7_75t_L g180 ( 
.A(n_0),
.B(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_301),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_1),
.B(n_302),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_3),
.Y(n_257)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_4),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_5),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_5),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_5),
.B(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_6),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_6),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_7),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_7),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_7),
.B(n_39),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_7),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_7),
.B(n_181),
.Y(n_240)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_8),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_9),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_9),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_9),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_9),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_9),
.B(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_11),
.Y(n_136)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

BUFx4f_ASAP7_75t_L g225 ( 
.A(n_12),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_13),
.Y(n_181)
);

BUFx8_ASAP7_75t_L g219 ( 
.A(n_13),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_269),
.Y(n_15)
);

INVxp67_ASAP7_75t_SL g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_231),
.B(n_263),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_196),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_158),
.B(n_195),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_125),
.B(n_157),
.Y(n_21)
);

OAI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_95),
.B(n_124),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_77),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_24),
.B(n_77),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_56),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_26),
.B(n_42),
.C(n_56),
.Y(n_126)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_28),
.B(n_34),
.C(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_28),
.B(n_44),
.C(n_169),
.Y(n_281)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_34),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_34),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_34),
.B(n_256),
.C(n_259),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_34),
.B(n_217),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_37),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_37),
.A2(n_154),
.B1(n_168),
.B2(n_174),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_40),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.C(n_52),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_44),
.B1(n_52),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_43),
.A2(n_44),
.B1(n_169),
.B2(n_173),
.Y(n_247)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_44),
.B(n_208),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g243 ( 
.A1(n_44),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_48),
.B1(n_79),
.B2(n_81),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_47),
.A2(n_48),
.B1(n_147),
.B2(n_150),
.Y(n_146)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_48),
.A2(n_107),
.B(n_116),
.C(n_148),
.Y(n_164)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_52),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_52),
.A2(n_80),
.B1(n_131),
.B2(n_143),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_52),
.B(n_293),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_89),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_53),
.B(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_58),
.A2(n_113),
.B(n_117),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_58),
.A2(n_69),
.B(n_76),
.Y(n_144)
);

NOR2x1_ASAP7_75t_R g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_59),
.A2(n_60),
.B1(n_87),
.B2(n_88),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_72),
.B(n_74),
.Y(n_71)
);

NAND2x1p5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_72),
.Y(n_74)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_98),
.B(n_101),
.C(n_107),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_98),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_69),
.A2(n_75),
.B1(n_98),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_71),
.A2(n_76),
.B1(n_137),
.B2(n_138),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_83),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_72),
.B(n_102),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_72),
.A2(n_93),
.B1(n_102),
.B2(n_105),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_72),
.A2(n_102),
.B(n_240),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_74),
.B(n_131),
.C(n_138),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.C(n_91),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_80),
.B(n_143),
.C(n_203),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_83),
.B(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_87),
.A2(n_88),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_88),
.B(n_218),
.C(n_222),
.Y(n_259)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_111),
.B(n_123),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_108),
.Y(n_96)
);

NOR2xp67_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_108),
.Y(n_123)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_98),
.B(n_115),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_98),
.B(n_116),
.C(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_98),
.A2(n_121),
.B1(n_207),
.B2(n_211),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_98),
.B(n_209),
.Y(n_245)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_102),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_102),
.A2(n_105),
.B1(n_169),
.B2(n_173),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_102),
.B(n_154),
.C(n_169),
.Y(n_228)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_119),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_118),
.B(n_122),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_115),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_116),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_121),
.B(n_208),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_127),
.Y(n_157)
);

XOR2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_145),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_144),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_129),
.B(n_144),
.C(n_145),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_137),
.B1(n_138),
.B2(n_143),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_151),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_152),
.C(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

AO22x1_ASAP7_75t_L g293 ( 
.A1(n_148),
.A2(n_149),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_194),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_194),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_175),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_162),
.C(n_175),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_167),
.C(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_166),
.B(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_193),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_183),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_183),
.C(n_193),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_182),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_190),
.B(n_192),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_190),
.Y(n_192)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_197),
.B(n_198),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_214),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_199),
.B(n_215),
.C(n_230),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_212),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_205),
.C(n_212),
.Y(n_233)
);

XNOR2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_230),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_226),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_228),
.C(n_229),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_262),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_262),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_236),
.C(n_248),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_248),
.B2(n_249),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_246),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_242),
.B2(n_243),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_243),
.C(n_246),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_260),
.B2(n_261),
.Y(n_251)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_261),
.C(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_253),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_299),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_272),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_287),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_286),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_284),
.B2(n_285),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);


endmodule