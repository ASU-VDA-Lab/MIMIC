module fake_ariane_622_n_1733 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1733);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1733;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_65),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_44),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_28),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_51),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_42),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_111),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_79),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_55),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_32),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_82),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_39),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_114),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_42),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_34),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_13),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_146),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_35),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_43),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_117),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_48),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_59),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_9),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_10),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

BUFx8_ASAP7_75t_SL g187 ( 
.A(n_151),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_61),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_57),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_20),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_37),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_17),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_120),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_149),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_136),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_2),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_69),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_3),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_80),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_121),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_13),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_70),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_1),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_52),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_28),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_49),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_9),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_19),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_22),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_107),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_115),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_37),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_132),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_128),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_21),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_22),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_125),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_112),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_25),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_50),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_25),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_38),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_38),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_104),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_23),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_40),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_1),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_91),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_83),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_84),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_29),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_145),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_41),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_16),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_63),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_11),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_4),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_12),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_137),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_92),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_75),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_2),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_73),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_60),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_20),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_105),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_66),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_144),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_71),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_135),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_139),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_4),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_96),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_19),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_68),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_47),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_15),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_64),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_32),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_103),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_141),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_74),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_77),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_90),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_47),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_31),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_102),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_72),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_54),
.Y(n_277)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_113),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_27),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_88),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_133),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_43),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_26),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_18),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_8),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_34),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_30),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_93),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_150),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_100),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_5),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_18),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_45),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_108),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_148),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_29),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_24),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_21),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_101),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_119),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_8),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_11),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_172),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_182),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_180),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_162),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_179),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_173),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_187),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_173),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_153),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_264),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_249),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_189),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_182),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_229),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_162),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_181),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_240),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_219),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_247),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_181),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_276),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_229),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_281),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_158),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_161),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_184),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_193),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_191),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_201),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_198),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_171),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_198),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_157),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_214),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_199),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_204),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_206),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_200),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_200),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_192),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_222),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_232),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_234),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_175),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_201),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_238),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_252),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_211),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_218),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_259),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_226),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_233),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_283),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_154),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_160),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_168),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_177),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_214),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g374 ( 
.A(n_262),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_178),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_256),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_244),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_183),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_306),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_287),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_306),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_323),
.B(n_287),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_306),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_257),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_163),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_305),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_331),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_332),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_307),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_308),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_312),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_308),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_329),
.A2(n_190),
.B(n_186),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_312),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_310),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_310),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_302),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_329),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_328),
.B(n_203),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_185),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_333),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_343),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_343),
.Y(n_407)
);

AND2x6_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_221),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_302),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_344),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_336),
.Y(n_411)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_166),
.C(n_157),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_317),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_351),
.A2(n_227),
.B(n_207),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_315),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

BUFx8_ASAP7_75t_L g420 ( 
.A(n_328),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_309),
.B(n_258),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_375),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_342),
.B(n_236),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_317),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_313),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_357),
.A2(n_223),
.B1(n_212),
.B2(n_241),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_372),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_324),
.B(n_197),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_372),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_378),
.B(n_185),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_317),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_342),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_358),
.B(n_196),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_326),
.B(n_185),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_334),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_339),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_317),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_340),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_317),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_317),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_314),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_317),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_358),
.B(n_237),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_327),
.B(n_196),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_314),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_381),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_429),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_404),
.B(n_317),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_SL g451 ( 
.A(n_438),
.B(n_230),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_404),
.B(n_317),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_397),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_384),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_388),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_404),
.B(n_335),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_341),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_432),
.B(n_376),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_397),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_408),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_432),
.B(n_348),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_394),
.B(n_346),
.Y(n_466)
);

BUFx4f_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_429),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_433),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_410),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_384),
.B(n_349),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_418),
.B(n_304),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_410),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g475 ( 
.A(n_421),
.B(n_361),
.C(n_350),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_387),
.B(n_362),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_436),
.B(n_364),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_387),
.B(n_221),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_398),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_446),
.A2(n_311),
.B1(n_354),
.B2(n_347),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_381),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_436),
.B(n_365),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_398),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_383),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_433),
.Y(n_487)
);

BUFx6f_ASAP7_75t_SL g488 ( 
.A(n_446),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_383),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_391),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_433),
.B(n_278),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_379),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_391),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_436),
.B(n_377),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_431),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_386),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_394),
.B(n_373),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_446),
.B(n_337),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_446),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_446),
.B(n_387),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_393),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_380),
.B(n_353),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_393),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_435),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_421),
.B(n_353),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_434),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_379),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_393),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_440),
.B(n_155),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_399),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_399),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_399),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_385),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_434),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_390),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_434),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_386),
.Y(n_520)
);

BUFx8_ASAP7_75t_SL g521 ( 
.A(n_411),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_435),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_379),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_385),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_435),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_379),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_428),
.A2(n_243),
.B1(n_169),
.B2(n_209),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_385),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_401),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_385),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_SL g531 ( 
.A1(n_396),
.A2(n_368),
.B(n_360),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_440),
.B(n_155),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_385),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_435),
.B(n_355),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_435),
.B(n_380),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_382),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_385),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_420),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_380),
.B(n_355),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_385),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_412),
.B(n_156),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_401),
.Y(n_542)
);

INVxp33_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

NOR3xp33_ASAP7_75t_L g544 ( 
.A(n_412),
.B(n_245),
.C(n_176),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_382),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_392),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_402),
.B(n_338),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_392),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_382),
.B(n_176),
.C(n_166),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_380),
.B(n_360),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_408),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_SL g552 ( 
.A(n_380),
.B(n_228),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_403),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_392),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_430),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_400),
.B(n_221),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_400),
.A2(n_359),
.B1(n_356),
.B2(n_243),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_392),
.Y(n_559)
);

OAI21xp33_ASAP7_75t_SL g560 ( 
.A1(n_396),
.A2(n_368),
.B(n_367),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_392),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_392),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_405),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_402),
.B(n_363),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_423),
.B(n_363),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_405),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_392),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_400),
.B(n_366),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_395),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_395),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_406),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_395),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_395),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_395),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_406),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_400),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_SL g577 ( 
.A(n_400),
.B(n_228),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_409),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_425),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_409),
.B(n_366),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_395),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_395),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_433),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_437),
.Y(n_584)
);

BUFx4f_ASAP7_75t_L g585 ( 
.A(n_416),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_409),
.B(n_156),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_407),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_407),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_409),
.B(n_367),
.Y(n_589)
);

AO21x2_ASAP7_75t_L g590 ( 
.A1(n_396),
.A2(n_267),
.B(n_289),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_409),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_419),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_414),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_439),
.B(n_278),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_419),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_413),
.Y(n_596)
);

INVx8_ASAP7_75t_L g597 ( 
.A(n_408),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_448),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_456),
.B(n_443),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_496),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_L g601 ( 
.A(n_496),
.B(n_428),
.C(n_284),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_454),
.B(n_420),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_500),
.B(n_420),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_500),
.B(n_420),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_450),
.B(n_439),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_502),
.B(n_420),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_448),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_564),
.B(n_419),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_596),
.Y(n_609)
);

O2A1O1Ixp33_ASAP7_75t_L g610 ( 
.A1(n_508),
.A2(n_539),
.B(n_589),
.C(n_550),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_552),
.A2(n_416),
.B1(n_422),
.B2(n_419),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_452),
.B(n_439),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_565),
.B(n_419),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_458),
.B(n_583),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_L g615 ( 
.A(n_466),
.B(n_284),
.C(n_282),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_547),
.B(n_422),
.Y(n_616)
);

NAND3xp33_ASAP7_75t_L g617 ( 
.A(n_475),
.B(n_285),
.C(n_282),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_458),
.B(n_439),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_520),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_498),
.B(n_591),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_472),
.B(n_423),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_458),
.B(n_439),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_486),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_456),
.B(n_443),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_591),
.B(n_422),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_583),
.B(n_413),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_453),
.B(n_422),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_486),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_463),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_489),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_596),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_488),
.A2(n_422),
.B1(n_414),
.B2(n_417),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_461),
.B(n_445),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_463),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_457),
.B(n_445),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_583),
.B(n_413),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_521),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_456),
.B(n_447),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_457),
.B(n_415),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_576),
.B(n_424),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_483),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_507),
.B(n_415),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_552),
.A2(n_416),
.B1(n_417),
.B2(n_426),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_501),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_489),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_507),
.B(n_426),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_522),
.B(n_427),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_522),
.B(n_427),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_488),
.A2(n_280),
.B1(n_288),
.B2(n_295),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_L g650 ( 
.A(n_520),
.B(n_292),
.C(n_299),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_483),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_456),
.A2(n_291),
.B1(n_299),
.B2(n_298),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_455),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_455),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_459),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_576),
.B(n_578),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_490),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_525),
.B(n_424),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_525),
.B(n_424),
.Y(n_659)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_509),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_545),
.B(n_285),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_505),
.B(n_441),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_459),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_505),
.B(n_441),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_490),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_568),
.B(n_441),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_576),
.B(n_442),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_568),
.B(n_442),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_580),
.B(n_449),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_580),
.B(n_442),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_577),
.A2(n_416),
.B1(n_265),
.B2(n_215),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_480),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_503),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_545),
.B(n_316),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_503),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_578),
.B(n_444),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_596),
.B(n_444),
.Y(n_677)
);

AO221x1_ASAP7_75t_L g678 ( 
.A1(n_451),
.A2(n_253),
.B1(n_221),
.B2(n_260),
.C(n_242),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_578),
.B(n_444),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_R g680 ( 
.A(n_579),
.B(n_291),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_501),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_468),
.B(n_164),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_480),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_SL g684 ( 
.A(n_521),
.B(n_215),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_476),
.A2(n_298),
.B1(n_292),
.B2(n_296),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_577),
.A2(n_265),
.B1(n_215),
.B2(n_231),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_501),
.B(n_316),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_485),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_465),
.B(n_296),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_518),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_477),
.B(n_263),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_467),
.B(n_159),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_467),
.B(n_159),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_467),
.B(n_165),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_495),
.B(n_165),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_504),
.Y(n_696)
);

AND2x2_ASAP7_75t_SL g697 ( 
.A(n_585),
.B(n_248),
.Y(n_697)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_484),
.B(n_272),
.C(n_273),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_494),
.B(n_275),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_R g700 ( 
.A(n_579),
.B(n_167),
.Y(n_700)
);

O2A1O1Ixp5_ASAP7_75t_L g701 ( 
.A1(n_541),
.A2(n_294),
.B(n_290),
.C(n_322),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_585),
.B(n_167),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_485),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_518),
.B(n_318),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_499),
.B(n_170),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_497),
.B(n_303),
.C(n_279),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_535),
.B(n_170),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_553),
.B(n_174),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_504),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_585),
.B(n_174),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_471),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_529),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_554),
.B(n_280),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_460),
.B(n_288),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_506),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_506),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_512),
.B(n_295),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_563),
.B(n_300),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_529),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_593),
.B(n_300),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_473),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_584),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_542),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_596),
.B(n_301),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_493),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_493),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_518),
.B(n_318),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_542),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_566),
.B(n_571),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_566),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_488),
.A2(n_265),
.B1(n_231),
.B2(n_408),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_571),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_575),
.B(n_301),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_511),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_575),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_511),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_587),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_596),
.B(n_278),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_587),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_478),
.B(n_278),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_482),
.B(n_319),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_532),
.B(n_231),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_478),
.B(n_278),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_588),
.B(n_188),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_479),
.B(n_194),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_479),
.B(n_195),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_592),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_479),
.A2(n_251),
.B1(n_205),
.B2(n_208),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_513),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_584),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_479),
.B(n_202),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_478),
.B(n_530),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_479),
.B(n_210),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_509),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_549),
.B(n_213),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_595),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_534),
.B(n_216),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_470),
.B(n_217),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_597),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_478),
.B(n_278),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_595),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_513),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_487),
.B(n_220),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_514),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_722),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_653),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_598),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_598),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_654),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_599),
.B(n_462),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_607),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_635),
.B(n_514),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_655),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_SL g775 ( 
.A1(n_756),
.A2(n_526),
.B(n_510),
.C(n_469),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_663),
.B(n_515),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_600),
.B(n_619),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_672),
.B(n_515),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_607),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_683),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_605),
.A2(n_560),
.B(n_531),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_688),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_637),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_703),
.B(n_519),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_711),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_712),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_751),
.B(n_543),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_629),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_621),
.A2(n_594),
.B(n_491),
.C(n_544),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_755),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_SL g791 ( 
.A(n_685),
.B(n_586),
.C(n_268),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_599),
.B(n_462),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_629),
.Y(n_793)
);

OR2x6_ASAP7_75t_L g794 ( 
.A(n_721),
.B(n_597),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_624),
.B(n_558),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_700),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_719),
.B(n_469),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_614),
.A2(n_491),
.B(n_594),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_634),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_615),
.B(n_556),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_723),
.B(n_469),
.Y(n_801)
);

AO21x2_ASAP7_75t_L g802 ( 
.A1(n_692),
.A2(n_590),
.B(n_540),
.Y(n_802)
);

AO22x1_ASAP7_75t_L g803 ( 
.A1(n_601),
.A2(n_557),
.B1(n_527),
.B2(n_474),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_728),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_697),
.A2(n_557),
.B1(n_517),
.B2(n_548),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_624),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_SL g807 ( 
.A(n_697),
.B(n_538),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_730),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_732),
.B(n_481),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_661),
.B(n_474),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_735),
.B(n_481),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_687),
.B(n_517),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_737),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_739),
.B(n_481),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_700),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_SL g816 ( 
.A1(n_686),
.A2(n_325),
.B1(n_322),
.B2(n_321),
.Y(n_816)
);

BUFx5_ASAP7_75t_L g817 ( 
.A(n_765),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_623),
.B(n_492),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_624),
.B(n_538),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_638),
.B(n_557),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_644),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_641),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_680),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_638),
.A2(n_557),
.B1(n_548),
.B2(n_582),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_641),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_651),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_760),
.B(n_464),
.Y(n_827)
);

INVx5_ASAP7_75t_L g828 ( 
.A(n_760),
.Y(n_828)
);

NOR3xp33_ASAP7_75t_SL g829 ( 
.A(n_652),
.B(n_239),
.C(n_224),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_628),
.B(n_492),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_630),
.B(n_492),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_704),
.B(n_510),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_645),
.B(n_510),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_760),
.B(n_464),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_727),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_SL g836 ( 
.A(n_681),
.B(n_690),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_725),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_638),
.Y(n_838)
);

AND3x2_ASAP7_75t_SL g839 ( 
.A(n_684),
.B(n_582),
.C(n_516),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_651),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_644),
.B(n_557),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_620),
.B(n_523),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_725),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_755),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_714),
.B(n_523),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_602),
.B(n_478),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_674),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_741),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_726),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_633),
.B(n_530),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_729),
.B(n_610),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_755),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_662),
.B(n_523),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_755),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_664),
.B(n_526),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_691),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_666),
.B(n_526),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_609),
.Y(n_858)
);

AND2x6_ASAP7_75t_SL g859 ( 
.A(n_689),
.B(n_699),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_639),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_649),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_726),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_682),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_668),
.B(n_548),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_698),
.B(n_557),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_734),
.Y(n_866)
);

NOR3xp33_ASAP7_75t_SL g867 ( 
.A(n_617),
.B(n_269),
.C(n_235),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_742),
.B(n_516),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_657),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_656),
.B(n_319),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_609),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_670),
.B(n_734),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_669),
.B(n_530),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_736),
.B(n_524),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_745),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_606),
.B(n_530),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_665),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_614),
.A2(n_528),
.B(n_533),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_736),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_750),
.B(n_524),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_750),
.B(n_528),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_717),
.A2(n_567),
.B1(n_540),
.B2(n_546),
.Y(n_882)
);

NOR2x1p5_ASAP7_75t_L g883 ( 
.A(n_706),
.B(n_320),
.Y(n_883)
);

NAND3xp33_ASAP7_75t_L g884 ( 
.A(n_650),
.B(n_573),
.C(n_574),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_665),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_609),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_695),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_763),
.B(n_533),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_632),
.B(n_530),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_707),
.B(n_320),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_671),
.A2(n_597),
.B1(n_590),
.B2(n_562),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_763),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_609),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_616),
.B(n_537),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_656),
.A2(n_660),
.B1(n_733),
.B2(n_642),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_631),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_631),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_631),
.Y(n_898)
);

AND2x6_ASAP7_75t_L g899 ( 
.A(n_631),
.B(n_537),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_705),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_646),
.A2(n_555),
.B1(n_546),
.B2(n_559),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_673),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_708),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_643),
.A2(n_597),
.B1(n_590),
.B2(n_555),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_748),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_608),
.B(n_559),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_613),
.B(n_562),
.Y(n_907)
);

INVx3_ASAP7_75t_SL g908 ( 
.A(n_724),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_713),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_673),
.B(n_675),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_718),
.B(n_567),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_675),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_640),
.B(n_321),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_647),
.B(n_325),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_757),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_696),
.B(n_570),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_762),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_627),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_658),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_696),
.Y(n_920)
);

NOR2xp67_ASAP7_75t_L g921 ( 
.A(n_720),
.B(n_570),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_709),
.B(n_572),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_648),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_640),
.B(n_572),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_709),
.B(n_573),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_744),
.B(n_561),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_715),
.B(n_574),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_715),
.Y(n_928)
);

AND2x2_ASAP7_75t_SL g929 ( 
.A(n_731),
.B(n_221),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_625),
.A2(n_0),
.B(n_3),
.C(n_5),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_716),
.B(n_581),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_758),
.B(n_0),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_716),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_659),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_738),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_724),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_611),
.B(n_581),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_753),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_759),
.B(n_581),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_618),
.A2(n_581),
.B(n_569),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_677),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_738),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_764),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_761),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_605),
.B(n_581),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_667),
.B(n_676),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_753),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_R g948 ( 
.A(n_677),
.B(n_569),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_768),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_767),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_851),
.A2(n_612),
.B(n_622),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_851),
.A2(n_612),
.B(n_622),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_798),
.A2(n_618),
.B(n_636),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_860),
.B(n_692),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_861),
.A2(n_667),
.B1(n_676),
.B2(n_679),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_909),
.B(n_777),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_810),
.B(n_693),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_943),
.B(n_693),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_876),
.A2(n_694),
.B(n_702),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_856),
.B(n_815),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_823),
.B(n_603),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_859),
.B(n_702),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_770),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_894),
.A2(n_626),
.B(n_636),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_899),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_SL g966 ( 
.A(n_807),
.B(n_604),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_894),
.A2(n_626),
.B(n_710),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_785),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_906),
.A2(n_710),
.B(n_679),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_906),
.A2(n_761),
.B(n_743),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_819),
.B(n_749),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_774),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_789),
.A2(n_752),
.B1(n_747),
.B2(n_746),
.Y(n_973)
);

CKINVDCx8_ASAP7_75t_R g974 ( 
.A(n_766),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_787),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_847),
.B(n_678),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_780),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_782),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_903),
.B(n_803),
.C(n_800),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_819),
.B(n_754),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_899),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_858),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_848),
.B(n_569),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_786),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_804),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_781),
.A2(n_743),
.B(n_740),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_907),
.A2(n_740),
.B(n_701),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_835),
.B(n_6),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_932),
.A2(n_6),
.B(n_7),
.C(n_10),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_923),
.B(n_569),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_812),
.B(n_569),
.Y(n_991)
);

AOI221xp5_ASAP7_75t_L g992 ( 
.A1(n_887),
.A2(n_254),
.B1(n_277),
.B2(n_274),
.C(n_271),
.Y(n_992)
);

NOR2xp67_ASAP7_75t_L g993 ( 
.A(n_796),
.B(n_561),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_863),
.B(n_806),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_838),
.B(n_561),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_907),
.A2(n_561),
.B(n_225),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_858),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_783),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_832),
.A2(n_270),
.B(n_250),
.C(n_255),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_820),
.B(n_551),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_872),
.A2(n_246),
.B(n_464),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_769),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_858),
.Y(n_1003)
);

NAND2x1p5_ASAP7_75t_L g1004 ( 
.A(n_821),
.B(n_464),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_872),
.A2(n_551),
.B(n_464),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_773),
.A2(n_551),
.B1(n_253),
.B2(n_14),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_841),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_773),
.B(n_7),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_808),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_845),
.A2(n_551),
.B(n_253),
.Y(n_1010)
);

AO32x1_ASAP7_75t_L g1011 ( 
.A1(n_890),
.A2(n_408),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_SL g1012 ( 
.A(n_829),
.B(n_253),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_930),
.A2(n_12),
.B(n_17),
.C(n_23),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_836),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_934),
.B(n_24),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_875),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_813),
.A2(n_26),
.B(n_27),
.C(n_30),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_852),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_784),
.A2(n_31),
.B(n_33),
.C(n_36),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_868),
.A2(n_253),
.B(n_551),
.C(n_278),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_908),
.Y(n_1021)
);

BUFx12f_ASAP7_75t_L g1022 ( 
.A(n_841),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_899),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_807),
.B(n_408),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_842),
.A2(n_855),
.B(n_853),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_842),
.A2(n_81),
.B(n_89),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_853),
.A2(n_76),
.B(n_87),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_905),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_883),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_790),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_795),
.B(n_33),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_870),
.B(n_36),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_895),
.B(n_828),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_929),
.A2(n_408),
.B1(n_278),
.B2(n_41),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_828),
.B(n_39),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_828),
.B(n_40),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_898),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_918),
.B(n_44),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_794),
.B(n_408),
.Y(n_1039)
);

AO21x2_ASAP7_75t_L g1040 ( 
.A1(n_846),
.A2(n_408),
.B(n_86),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_899),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_772),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_855),
.A2(n_45),
.B(n_46),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_857),
.A2(n_95),
.B(n_53),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_828),
.B(n_48),
.Y(n_1045)
);

AOI21x1_ASAP7_75t_L g1046 ( 
.A1(n_939),
.A2(n_56),
.B(n_58),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_914),
.B(n_62),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_936),
.B(n_67),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_816),
.A2(n_85),
.B1(n_116),
.B2(n_122),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_776),
.A2(n_123),
.B1(n_127),
.B2(n_131),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_915),
.Y(n_1051)
);

BUFx12f_ASAP7_75t_L g1052 ( 
.A(n_790),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_870),
.B(n_138),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_914),
.B(n_140),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_784),
.A2(n_791),
.B(n_914),
.C(n_775),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_790),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_936),
.B(n_771),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_SL g1058 ( 
.A(n_884),
.B(n_797),
.C(n_809),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_857),
.A2(n_864),
.B(n_926),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_776),
.A2(n_778),
.B(n_873),
.C(n_850),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_917),
.Y(n_1061)
);

OAI21xp33_ASAP7_75t_L g1062 ( 
.A1(n_781),
.A2(n_778),
.B(n_867),
.Y(n_1062)
);

AO21x1_ASAP7_75t_L g1063 ( 
.A1(n_889),
.A2(n_911),
.B(n_946),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_792),
.B(n_946),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_779),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_837),
.B(n_843),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_797),
.A2(n_833),
.B(n_831),
.C(n_830),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_849),
.B(n_862),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_801),
.A2(n_818),
.B(n_811),
.C(n_833),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_844),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_SL g1071 ( 
.A(n_941),
.B(n_794),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_864),
.A2(n_878),
.B(n_940),
.Y(n_1072)
);

BUFx10_ASAP7_75t_L g1073 ( 
.A(n_865),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_945),
.A2(n_919),
.B(n_931),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_935),
.A2(n_942),
.B(n_944),
.C(n_866),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_945),
.A2(n_931),
.B(n_831),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_913),
.A2(n_865),
.B1(n_879),
.B2(n_892),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_893),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_794),
.B(n_844),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_913),
.A2(n_788),
.B1(n_793),
.B2(n_799),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_SL g1081 ( 
.A1(n_886),
.A2(n_896),
.B(n_809),
.C(n_801),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_941),
.B(n_844),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_SL g1083 ( 
.A(n_811),
.B(n_830),
.C(n_818),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_928),
.B(n_933),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_854),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_901),
.A2(n_814),
.B(n_874),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_938),
.B(n_947),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_814),
.A2(n_888),
.B(n_881),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_886),
.B(n_896),
.C(n_921),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_854),
.B(n_898),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_898),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_938),
.B(n_947),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_941),
.A2(n_805),
.B1(n_824),
.B2(n_893),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1031),
.A2(n_882),
.B(n_937),
.C(n_941),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1034),
.A2(n_881),
.B1(n_880),
.B2(n_874),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1025),
.A2(n_880),
.B(n_888),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1062),
.B(n_1066),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_1023),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1088),
.A2(n_871),
.B(n_897),
.Y(n_1099)
);

AND2x6_ASAP7_75t_SL g1100 ( 
.A(n_962),
.B(n_924),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_989),
.B(n_947),
.C(n_938),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1062),
.B(n_817),
.Y(n_1102)
);

AOI211x1_ASAP7_75t_L g1103 ( 
.A1(n_1043),
.A2(n_927),
.B(n_916),
.C(n_922),
.Y(n_1103)
);

O2A1O1Ixp5_ASAP7_75t_L g1104 ( 
.A1(n_1012),
.A2(n_927),
.B(n_925),
.C(n_922),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1072),
.A2(n_925),
.B(n_916),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1068),
.B(n_817),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_968),
.Y(n_1107)
);

NAND3x1_ASAP7_75t_L g1108 ( 
.A(n_979),
.B(n_839),
.C(n_910),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_1023),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_953),
.A2(n_1059),
.B(n_1076),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_955),
.B(n_817),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_950),
.Y(n_1112)
);

AOI221x1_ASAP7_75t_L g1113 ( 
.A1(n_1006),
.A2(n_839),
.B1(n_920),
.B2(n_822),
.C(n_825),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_955),
.B(n_1008),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_958),
.B(n_854),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1032),
.B(n_877),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_975),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_SL g1118 ( 
.A(n_992),
.B(n_948),
.C(n_891),
.Y(n_1118)
);

AO32x2_ASAP7_75t_L g1119 ( 
.A1(n_1093),
.A2(n_802),
.A3(n_817),
.B1(n_924),
.B2(n_885),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_956),
.B(n_924),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_994),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_986),
.A2(n_904),
.B(n_912),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1074),
.A2(n_902),
.B(n_869),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_1016),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_SL g1125 ( 
.A(n_965),
.B(n_817),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_957),
.B(n_826),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1084),
.B(n_840),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1067),
.A2(n_802),
.B(n_834),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_967),
.A2(n_827),
.B(n_834),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_969),
.A2(n_827),
.B(n_970),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1021),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_991),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1002),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1086),
.A2(n_959),
.B(n_987),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_973),
.A2(n_1020),
.A3(n_1075),
.B(n_964),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_1022),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1034),
.A2(n_1015),
.B1(n_1009),
.B2(n_978),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1052),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1083),
.B(n_963),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_974),
.B(n_960),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1018),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_972),
.B(n_977),
.Y(n_1142)
);

OA22x2_ASAP7_75t_L g1143 ( 
.A1(n_1077),
.A2(n_1029),
.B1(n_984),
.B2(n_985),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_951),
.A2(n_952),
.B(n_1046),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1010),
.A2(n_1069),
.B(n_1060),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1064),
.B(n_1077),
.Y(n_1146)
);

OAI22x1_ASAP7_75t_L g1147 ( 
.A1(n_1057),
.A2(n_1054),
.B1(n_1051),
.B2(n_1061),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1081),
.A2(n_1033),
.B(n_1055),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1028),
.B(n_1042),
.Y(n_1149)
);

AO21x1_ASAP7_75t_L g1150 ( 
.A1(n_966),
.A2(n_1013),
.B(n_1047),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_988),
.B(n_998),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1065),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1026),
.A2(n_1027),
.B(n_1044),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1082),
.A2(n_1001),
.B(n_1005),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1087),
.B(n_1092),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_996),
.A2(n_1050),
.A3(n_954),
.B(n_999),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_983),
.A2(n_1038),
.A3(n_1041),
.B(n_990),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1048),
.A2(n_1056),
.B(n_980),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1017),
.A2(n_1019),
.B(n_1045),
.C(n_1036),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_SL g1160 ( 
.A1(n_976),
.A2(n_1053),
.B(n_995),
.Y(n_1160)
);

NAND3x1_ASAP7_75t_L g1161 ( 
.A(n_1089),
.B(n_1014),
.C(n_1056),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_966),
.A2(n_1024),
.B(n_965),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1041),
.A2(n_1070),
.A3(n_1040),
.B(n_1011),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1078),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_SL g1165 ( 
.A1(n_1085),
.A2(n_1049),
.B(n_1080),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_965),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1058),
.B(n_1071),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1090),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1030),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_961),
.A2(n_1035),
.B(n_971),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_SL g1171 ( 
.A(n_1007),
.B(n_1071),
.C(n_1024),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1073),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_993),
.A2(n_1039),
.B(n_981),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_981),
.A2(n_1011),
.B(n_1040),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_981),
.A2(n_1039),
.B(n_1000),
.C(n_997),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1004),
.A2(n_1073),
.B(n_1079),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1000),
.A2(n_982),
.B(n_997),
.C(n_1003),
.Y(n_1177)
);

NAND2x1_ASAP7_75t_L g1178 ( 
.A(n_982),
.B(n_997),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1079),
.B(n_1003),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1003),
.Y(n_1180)
);

NAND2x1_ASAP7_75t_L g1181 ( 
.A(n_1037),
.B(n_1091),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1079),
.Y(n_1182)
);

AO32x2_ASAP7_75t_L g1183 ( 
.A1(n_1011),
.A2(n_1093),
.A3(n_848),
.B1(n_973),
.B2(n_1006),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1037),
.A2(n_1063),
.A3(n_1025),
.B(n_973),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_1091),
.B(n_579),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1032),
.B(n_536),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_951),
.A2(n_789),
.B(n_952),
.Y(n_1187)
);

NAND3xp33_ASAP7_75t_L g1188 ( 
.A(n_1031),
.B(n_989),
.C(n_742),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1032),
.B(n_536),
.Y(n_1189)
);

AND3x1_ASAP7_75t_L g1190 ( 
.A(n_962),
.B(n_684),
.C(n_473),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_1025),
.A2(n_1072),
.B(n_1074),
.Y(n_1191)
);

NOR4xp25_ASAP7_75t_L g1192 ( 
.A(n_989),
.B(n_1013),
.C(n_1019),
.D(n_1017),
.Y(n_1192)
);

AO21x1_ASAP7_75t_L g1193 ( 
.A1(n_1034),
.A2(n_1031),
.B(n_1055),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_950),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1025),
.A2(n_851),
.B(n_1072),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_956),
.A2(n_584),
.B1(n_579),
.B2(n_722),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_950),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_950),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1025),
.A2(n_851),
.B(n_1088),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1062),
.B(n_773),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1062),
.B(n_773),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1063),
.A2(n_1025),
.A3(n_973),
.B(n_1072),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1072),
.A2(n_1025),
.B(n_1059),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1072),
.A2(n_959),
.B(n_1033),
.Y(n_1204)
);

AOI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1072),
.A2(n_959),
.B(n_1033),
.Y(n_1205)
);

INVxp67_ASAP7_75t_SL g1206 ( 
.A(n_994),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1062),
.B(n_773),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_968),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1062),
.B(n_773),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_974),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1025),
.A2(n_851),
.B(n_1088),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1025),
.A2(n_851),
.B(n_1088),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_950),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_949),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1031),
.A2(n_428),
.B1(n_313),
.B2(n_334),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1072),
.A2(n_1025),
.B(n_1059),
.Y(n_1216)
);

CKINVDCx11_ASAP7_75t_R g1217 ( 
.A(n_974),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_950),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1022),
.Y(n_1219)
);

NAND2xp33_ASAP7_75t_L g1220 ( 
.A(n_1083),
.B(n_722),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_950),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1031),
.A2(n_958),
.B(n_1034),
.C(n_1062),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1034),
.A2(n_851),
.B1(n_957),
.B2(n_1008),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1031),
.B(n_989),
.C(n_742),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_951),
.A2(n_789),
.B(n_952),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_950),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_SL g1227 ( 
.A1(n_1222),
.A2(n_1114),
.B(n_1223),
.C(n_1200),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1223),
.A2(n_1224),
.B(n_1188),
.Y(n_1228)
);

NAND2xp33_ASAP7_75t_R g1229 ( 
.A(n_1162),
.B(n_1167),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1137),
.A2(n_1193),
.B1(n_1215),
.B2(n_1114),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1168),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1113),
.A2(n_1174),
.A3(n_1128),
.B(n_1137),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1139),
.A2(n_1196),
.B1(n_1101),
.B2(n_1097),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1217),
.Y(n_1234)
);

OAI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1139),
.A2(n_1097),
.B1(n_1146),
.B2(n_1206),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1185),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1142),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1126),
.B(n_1107),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1220),
.A2(n_1159),
.B(n_1192),
.C(n_1201),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1179),
.B(n_1182),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1107),
.B(n_1208),
.Y(n_1241)
);

INVx6_ASAP7_75t_L g1242 ( 
.A(n_1138),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1118),
.A2(n_1143),
.B1(n_1095),
.B2(n_1146),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_SL g1244 ( 
.A1(n_1200),
.A2(n_1209),
.B(n_1201),
.C(n_1207),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1190),
.A2(n_1120),
.B1(n_1189),
.B2(n_1186),
.Y(n_1245)
);

OAI21xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1106),
.A2(n_1209),
.B(n_1207),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1110),
.A2(n_1130),
.B(n_1195),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1143),
.A2(n_1095),
.B1(n_1147),
.B2(n_1150),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1142),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1208),
.B(n_1167),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1154),
.A2(n_1105),
.B(n_1211),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1199),
.A2(n_1212),
.B(n_1145),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_SL g1253 ( 
.A1(n_1170),
.A2(n_1148),
.B(n_1106),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1153),
.A2(n_1096),
.B(n_1225),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1096),
.A2(n_1225),
.B(n_1187),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1151),
.B(n_1116),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1111),
.A2(n_1125),
.B1(n_1198),
.B2(n_1213),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1121),
.B(n_1117),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1187),
.A2(n_1122),
.B(n_1129),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1099),
.A2(n_1174),
.B(n_1148),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1160),
.A2(n_1104),
.B(n_1203),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1210),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1112),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1203),
.A2(n_1216),
.B(n_1102),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1202),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1192),
.A2(n_1111),
.B(n_1170),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1102),
.A2(n_1094),
.B(n_1132),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1140),
.A2(n_1124),
.B1(n_1161),
.B2(n_1155),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1182),
.B(n_1175),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1158),
.A2(n_1127),
.B(n_1149),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1194),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1115),
.A2(n_1108),
.B(n_1125),
.Y(n_1272)
);

BUFx8_ASAP7_75t_L g1273 ( 
.A(n_1138),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1155),
.A2(n_1131),
.B1(n_1103),
.B2(n_1109),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1197),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1164),
.B(n_1141),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1218),
.Y(n_1277)
);

INVx6_ASAP7_75t_L g1278 ( 
.A(n_1138),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1216),
.A2(n_1123),
.B(n_1098),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1173),
.A2(n_1176),
.B(n_1165),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1127),
.A2(n_1149),
.B(n_1226),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1221),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1180),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1133),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1152),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1214),
.A2(n_1171),
.B1(n_1169),
.B2(n_1219),
.Y(n_1286)
);

BUFx12f_ASAP7_75t_L g1287 ( 
.A(n_1136),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1136),
.A2(n_1219),
.B1(n_1172),
.B2(n_1134),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1136),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1178),
.A2(n_1181),
.B(n_1191),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1100),
.B(n_1219),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1191),
.A2(n_1202),
.B(n_1184),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1177),
.A2(n_1157),
.B(n_1156),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1202),
.A2(n_1184),
.B(n_1135),
.Y(n_1294)
);

AO32x2_ASAP7_75t_L g1295 ( 
.A1(n_1119),
.A2(n_1183),
.A3(n_1184),
.B1(n_1157),
.B2(n_1163),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1135),
.A2(n_1163),
.B(n_1157),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1135),
.A2(n_1163),
.B(n_1156),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1183),
.A2(n_1119),
.B(n_1156),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1166),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1119),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1183),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1180),
.A2(n_1144),
.B(n_1204),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1180),
.A2(n_1211),
.B(n_1199),
.Y(n_1303)
);

OAI221xp5_ASAP7_75t_L g1304 ( 
.A1(n_1188),
.A2(n_1224),
.B1(n_1192),
.B2(n_1222),
.C(n_1223),
.Y(n_1304)
);

AO32x2_ASAP7_75t_L g1305 ( 
.A1(n_1223),
.A2(n_1137),
.A3(n_1095),
.B1(n_1093),
.B2(n_1119),
.Y(n_1305)
);

AO32x2_ASAP7_75t_L g1306 ( 
.A1(n_1223),
.A2(n_1137),
.A3(n_1095),
.B1(n_1093),
.B2(n_1119),
.Y(n_1306)
);

AOI221xp5_ASAP7_75t_L g1307 ( 
.A1(n_1223),
.A2(n_1137),
.B1(n_384),
.B2(n_1224),
.C(n_1188),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1188),
.A2(n_722),
.B1(n_900),
.B2(n_887),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1126),
.B(n_1107),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1144),
.A2(n_1205),
.B(n_1204),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1144),
.A2(n_1205),
.B(n_1204),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1137),
.A2(n_1223),
.B1(n_428),
.B2(n_1188),
.Y(n_1312)
);

NAND2xp33_ASAP7_75t_R g1313 ( 
.A(n_1162),
.B(n_1083),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1222),
.A2(n_1114),
.B(n_1223),
.C(n_1081),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1142),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1188),
.A2(n_722),
.B1(n_900),
.B2(n_887),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1202),
.Y(n_1317)
);

NAND2x1p5_ASAP7_75t_L g1318 ( 
.A(n_1166),
.B(n_965),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1199),
.A2(n_1212),
.B(n_1211),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_SL g1320 ( 
.A1(n_1222),
.A2(n_1114),
.B(n_1223),
.C(n_1081),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1182),
.B(n_1179),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1202),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1199),
.A2(n_1212),
.B(n_1211),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_SL g1324 ( 
.A1(n_1222),
.A2(n_1114),
.B(n_1223),
.C(n_1081),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1166),
.B(n_965),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_SL g1326 ( 
.A(n_1137),
.B(n_1223),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1142),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1166),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1144),
.A2(n_1205),
.B(n_1204),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1199),
.A2(n_1212),
.B(n_1211),
.Y(n_1330)
);

AOI222xp33_ASAP7_75t_L g1331 ( 
.A1(n_1215),
.A2(n_428),
.B1(n_1137),
.B2(n_171),
.C1(n_197),
.C2(n_223),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1222),
.A2(n_1034),
.B(n_1137),
.C(n_1223),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1137),
.A2(n_1223),
.B1(n_428),
.B2(n_1188),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1144),
.A2(n_1205),
.B(n_1204),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1168),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1166),
.B(n_965),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1142),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1137),
.A2(n_1223),
.B1(n_428),
.B2(n_1188),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1185),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1123),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1168),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1142),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1260),
.A2(n_1323),
.B(n_1319),
.Y(n_1343)
);

AOI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1312),
.A2(n_1333),
.B1(n_1338),
.B2(n_1230),
.C(n_1307),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1330),
.A2(n_1292),
.B(n_1297),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1301),
.B(n_1305),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1236),
.Y(n_1347)
);

O2A1O1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1332),
.A2(n_1304),
.B(n_1228),
.C(n_1312),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1250),
.B(n_1237),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1301),
.B(n_1305),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1333),
.A2(n_1338),
.B1(n_1332),
.B2(n_1230),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1241),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1305),
.B(n_1306),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1233),
.A2(n_1239),
.B(n_1235),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1250),
.B(n_1249),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1305),
.B(n_1306),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1321),
.B(n_1269),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1306),
.B(n_1266),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1298),
.B(n_1326),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1227),
.A2(n_1324),
.B(n_1314),
.C(n_1320),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1227),
.A2(n_1324),
.B(n_1314),
.C(n_1320),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1239),
.A2(n_1268),
.B(n_1272),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1257),
.A2(n_1267),
.B(n_1274),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1283),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1243),
.A2(n_1316),
.B1(n_1308),
.B2(n_1248),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1315),
.Y(n_1366)
);

AOI211xp5_ASAP7_75t_L g1367 ( 
.A1(n_1326),
.A2(n_1257),
.B(n_1246),
.C(n_1244),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1243),
.A2(n_1248),
.B1(n_1245),
.B2(n_1339),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1327),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1321),
.B(n_1269),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1303),
.A2(n_1255),
.B(n_1244),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1321),
.B(n_1240),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1238),
.A2(n_1309),
.B1(n_1242),
.B2(n_1278),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1267),
.A2(n_1336),
.B(n_1325),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1254),
.A2(n_1252),
.B(n_1296),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1261),
.A2(n_1247),
.B(n_1294),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1337),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1267),
.A2(n_1336),
.B(n_1318),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1271),
.A2(n_1275),
.B1(n_1277),
.B2(n_1282),
.C(n_1342),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1264),
.A2(n_1293),
.B(n_1251),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1242),
.A2(n_1278),
.B1(n_1286),
.B2(n_1256),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1234),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1331),
.A2(n_1253),
.B(n_1258),
.C(n_1265),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1265),
.B(n_1317),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1281),
.B(n_1276),
.Y(n_1385)
);

O2A1O1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1322),
.A2(n_1289),
.B(n_1335),
.C(n_1291),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1278),
.A2(n_1286),
.B1(n_1231),
.B2(n_1341),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1290),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1295),
.B(n_1298),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1234),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1287),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1302),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1281),
.B(n_1240),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1231),
.A2(n_1341),
.B1(n_1288),
.B2(n_1287),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1295),
.B(n_1298),
.Y(n_1395)
);

INVxp67_ASAP7_75t_SL g1396 ( 
.A(n_1270),
.Y(n_1396)
);

CKINVDCx16_ASAP7_75t_R g1397 ( 
.A(n_1313),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1273),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1295),
.B(n_1232),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1295),
.B(n_1232),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1232),
.B(n_1270),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1313),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1229),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1310),
.A2(n_1334),
.B(n_1329),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1232),
.B(n_1300),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1311),
.A2(n_1279),
.B(n_1259),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1262),
.A2(n_1273),
.B1(n_1328),
.B2(n_1299),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1299),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1284),
.A2(n_1285),
.B1(n_1340),
.B2(n_1280),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1301),
.B(n_1306),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1263),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1312),
.A2(n_1333),
.B1(n_1338),
.B2(n_1332),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1326),
.A2(n_1332),
.B(n_1223),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1301),
.B(n_1306),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1312),
.A2(n_1338),
.B1(n_1333),
.B2(n_1304),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1260),
.A2(n_1323),
.B(n_1319),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1326),
.A2(n_1332),
.B(n_1223),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1263),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1299),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1250),
.B(n_1237),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1263),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1301),
.B(n_1306),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1260),
.A2(n_1323),
.B(n_1319),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1250),
.B(n_1237),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1250),
.B(n_1237),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1250),
.B(n_1237),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1234),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1401),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1388),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1403),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1388),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1359),
.B(n_1358),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1359),
.B(n_1358),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1401),
.Y(n_1434)
);

AO21x2_ASAP7_75t_L g1435 ( 
.A1(n_1363),
.A2(n_1396),
.B(n_1371),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1363),
.A2(n_1399),
.B(n_1400),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1413),
.A2(n_1417),
.B(n_1400),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1385),
.Y(n_1438)
);

AO21x1_ASAP7_75t_SL g1439 ( 
.A1(n_1367),
.A2(n_1418),
.B(n_1411),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1421),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1405),
.B(n_1353),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1393),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1399),
.A2(n_1354),
.B(n_1409),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1353),
.B(n_1356),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1366),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1374),
.B(n_1378),
.Y(n_1446)
);

INVxp67_ASAP7_75t_R g1447 ( 
.A(n_1407),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1405),
.B(n_1356),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1346),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1389),
.B(n_1395),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1351),
.A2(n_1412),
.B(n_1389),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1415),
.A2(n_1344),
.B1(n_1365),
.B2(n_1397),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1346),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1368),
.A2(n_1402),
.B1(n_1348),
.B2(n_1410),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1362),
.B(n_1369),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1395),
.B(n_1350),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1350),
.B(n_1422),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1377),
.B(n_1410),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1392),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1360),
.A2(n_1361),
.B(n_1414),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1384),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1392),
.A2(n_1416),
.B(n_1343),
.Y(n_1462)
);

OAI321xp33_ASAP7_75t_L g1463 ( 
.A1(n_1383),
.A2(n_1381),
.A3(n_1387),
.B1(n_1373),
.B2(n_1426),
.C(n_1349),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1352),
.B(n_1424),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1380),
.B(n_1416),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1380),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1355),
.B(n_1425),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1357),
.B(n_1370),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1380),
.B(n_1416),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1376),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1345),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1420),
.B(n_1379),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1456),
.B(n_1423),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1457),
.B(n_1345),
.Y(n_1474)
);

NOR2xp67_ASAP7_75t_L g1475 ( 
.A(n_1429),
.B(n_1370),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1468),
.B(n_1357),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1431),
.Y(n_1477)
);

INVx1_ASAP7_75t_SL g1478 ( 
.A(n_1430),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1457),
.B(n_1437),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1442),
.B(n_1364),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1455),
.B(n_1347),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1442),
.B(n_1386),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1440),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1452),
.A2(n_1394),
.B1(n_1370),
.B2(n_1372),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1470),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1440),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1468),
.B(n_1372),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1451),
.B(n_1430),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1470),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1451),
.B(n_1375),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1432),
.B(n_1406),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1437),
.B(n_1406),
.Y(n_1492)
);

NOR2x1_ASAP7_75t_L g1493 ( 
.A(n_1435),
.B(n_1419),
.Y(n_1493)
);

NOR2x1_ASAP7_75t_L g1494 ( 
.A(n_1435),
.B(n_1455),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1437),
.B(n_1406),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1470),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1437),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1452),
.A2(n_1427),
.B1(n_1390),
.B2(n_1382),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1437),
.B(n_1404),
.Y(n_1499)
);

NAND2x1p5_ASAP7_75t_L g1500 ( 
.A(n_1437),
.B(n_1404),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1451),
.B(n_1408),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1484),
.A2(n_1451),
.B1(n_1436),
.B2(n_1443),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1478),
.B(n_1445),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1498),
.A2(n_1451),
.B1(n_1454),
.B2(n_1436),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1483),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1483),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_R g1507 ( 
.A(n_1498),
.B(n_1382),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1476),
.B(n_1468),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1483),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1478),
.B(n_1432),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1501),
.B(n_1432),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1482),
.B(n_1445),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1479),
.A2(n_1436),
.B1(n_1443),
.B2(n_1434),
.Y(n_1513)
);

OAI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1488),
.A2(n_1454),
.B1(n_1472),
.B2(n_1433),
.C(n_1438),
.Y(n_1514)
);

OAI211xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1494),
.A2(n_1472),
.B(n_1471),
.C(n_1459),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1501),
.B(n_1433),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_1497),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1481),
.Y(n_1518)
);

AOI21xp33_ASAP7_75t_L g1519 ( 
.A1(n_1494),
.A2(n_1443),
.B(n_1463),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1488),
.A2(n_1436),
.B1(n_1443),
.B2(n_1439),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1490),
.A2(n_1463),
.B1(n_1434),
.B2(n_1428),
.C(n_1466),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_R g1522 ( 
.A(n_1481),
.B(n_1390),
.Y(n_1522)
);

NOR4xp25_ASAP7_75t_SL g1523 ( 
.A(n_1477),
.B(n_1427),
.C(n_1466),
.D(n_1431),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_L g1524 ( 
.A(n_1480),
.B(n_1460),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1486),
.Y(n_1525)
);

AOI322xp5_ASAP7_75t_L g1526 ( 
.A1(n_1479),
.A2(n_1448),
.A3(n_1441),
.B1(n_1428),
.B2(n_1444),
.C1(n_1438),
.C2(n_1453),
.Y(n_1526)
);

AOI33xp33_ASAP7_75t_L g1527 ( 
.A1(n_1479),
.A2(n_1461),
.A3(n_1453),
.B1(n_1449),
.B2(n_1469),
.B3(n_1465),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1487),
.B(n_1450),
.Y(n_1528)
);

OR2x6_ASAP7_75t_L g1529 ( 
.A(n_1493),
.B(n_1446),
.Y(n_1529)
);

OAI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1490),
.A2(n_1433),
.B1(n_1466),
.B2(n_1467),
.C(n_1464),
.Y(n_1530)
);

NOR3xp33_ASAP7_75t_L g1531 ( 
.A(n_1497),
.B(n_1469),
.C(n_1465),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_R g1532 ( 
.A(n_1479),
.B(n_1398),
.Y(n_1532)
);

NOR4xp25_ASAP7_75t_SL g1533 ( 
.A(n_1477),
.B(n_1431),
.C(n_1408),
.D(n_1439),
.Y(n_1533)
);

OAI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1484),
.A2(n_1447),
.B1(n_1450),
.B2(n_1467),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1480),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1484),
.A2(n_1447),
.B1(n_1444),
.B2(n_1458),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1482),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1519),
.A2(n_1497),
.B(n_1499),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1524),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1521),
.A2(n_1435),
.B(n_1497),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1502),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1511),
.B(n_1491),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1516),
.B(n_1491),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1505),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1520),
.A2(n_1499),
.B(n_1495),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1506),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1509),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1531),
.B(n_1474),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1517),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1508),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1517),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1508),
.B(n_1475),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1529),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1527),
.B(n_1473),
.Y(n_1554)
);

OA21x2_ASAP7_75t_L g1555 ( 
.A1(n_1520),
.A2(n_1499),
.B(n_1495),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1525),
.Y(n_1556)
);

INVxp67_ASAP7_75t_SL g1557 ( 
.A(n_1531),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1537),
.Y(n_1558)
);

NAND3xp33_ASAP7_75t_SL g1559 ( 
.A(n_1513),
.B(n_1495),
.C(n_1492),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1518),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1504),
.A2(n_1492),
.B(n_1499),
.Y(n_1561)
);

OAI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1504),
.A2(n_1500),
.B(n_1462),
.Y(n_1562)
);

NOR3xp33_ASAP7_75t_L g1563 ( 
.A(n_1515),
.B(n_1492),
.C(n_1493),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1550),
.B(n_1528),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1550),
.B(n_1526),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1560),
.B(n_1534),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1544),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1560),
.B(n_1512),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1544),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1546),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1545),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1559),
.B(n_1491),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1558),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1550),
.B(n_1533),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1558),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1545),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1557),
.B(n_1535),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1557),
.B(n_1546),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1550),
.B(n_1523),
.Y(n_1579)
);

CKINVDCx16_ASAP7_75t_R g1580 ( 
.A(n_1559),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1545),
.Y(n_1581)
);

NAND3xp33_ASAP7_75t_L g1582 ( 
.A(n_1561),
.B(n_1513),
.C(n_1515),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1548),
.B(n_1503),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1561),
.B(n_1563),
.Y(n_1584)
);

NAND2xp67_ASAP7_75t_L g1585 ( 
.A(n_1541),
.B(n_1485),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1548),
.B(n_1474),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1554),
.A2(n_1532),
.B1(n_1514),
.B2(n_1534),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1556),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1556),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1548),
.B(n_1460),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1554),
.B(n_1530),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1562),
.A2(n_1496),
.B(n_1489),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1547),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1563),
.B(n_1460),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_L g1596 ( 
.A(n_1540),
.B(n_1536),
.C(n_1489),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1547),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1547),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_L g1599 ( 
.A(n_1545),
.B(n_1477),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1573),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

NOR2x1p5_ASAP7_75t_SL g1602 ( 
.A(n_1571),
.B(n_1549),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1580),
.B(n_1576),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1594),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1573),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1580),
.B(n_1576),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1571),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1594),
.Y(n_1608)
);

INVxp67_ASAP7_75t_SL g1609 ( 
.A(n_1575),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1591),
.B(n_1545),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1597),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1597),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1584),
.B(n_1565),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1566),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1598),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1568),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1577),
.B(n_1510),
.Y(n_1617)
);

AOI31xp33_ASAP7_75t_L g1618 ( 
.A1(n_1584),
.A2(n_1541),
.A3(n_1552),
.B(n_1553),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1588),
.B(n_1541),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1584),
.B(n_1565),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1584),
.B(n_1552),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1564),
.B(n_1545),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1578),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1564),
.B(n_1555),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1578),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1598),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1579),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1599),
.B(n_1555),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1599),
.B(n_1555),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1588),
.B(n_1541),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1567),
.B(n_1591),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1569),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1592),
.B(n_1555),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1582),
.A2(n_1555),
.B1(n_1538),
.B2(n_1460),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1604),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1628),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1604),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1608),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1601),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1601),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1605),
.B(n_1571),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1608),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1611),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1605),
.B(n_1574),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1610),
.B(n_1582),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1634),
.B(n_1587),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1610),
.A2(n_1581),
.B1(n_1555),
.B2(n_1596),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1600),
.B(n_1596),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1609),
.B(n_1581),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1616),
.B(n_1595),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1621),
.B(n_1574),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1614),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1613),
.B(n_1581),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1621),
.B(n_1579),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1603),
.B(n_1592),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1612),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1612),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1628),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1640),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1656),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1646),
.A2(n_1634),
.B1(n_1606),
.B2(n_1613),
.C(n_1620),
.Y(n_1662)
);

INVxp67_ASAP7_75t_SL g1663 ( 
.A(n_1640),
.Y(n_1663)
);

AOI222xp33_ASAP7_75t_L g1664 ( 
.A1(n_1647),
.A2(n_1606),
.B1(n_1620),
.B2(n_1629),
.C1(n_1602),
.C2(n_1624),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1645),
.A2(n_1603),
.B1(n_1572),
.B2(n_1629),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1653),
.B(n_1623),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1656),
.B(n_1631),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1645),
.A2(n_1627),
.B1(n_1622),
.B2(n_1624),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1644),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1644),
.Y(n_1670)
);

OAI32xp33_ASAP7_75t_L g1671 ( 
.A1(n_1648),
.A2(n_1633),
.A3(n_1572),
.B1(n_1654),
.B2(n_1636),
.Y(n_1671)
);

OAI32xp33_ASAP7_75t_L g1672 ( 
.A1(n_1636),
.A2(n_1633),
.A3(n_1623),
.B1(n_1630),
.B2(n_1619),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1637),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1659),
.A2(n_1618),
.B1(n_1590),
.B2(n_1622),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1637),
.Y(n_1675)
);

OAI222xp33_ASAP7_75t_L g1676 ( 
.A1(n_1649),
.A2(n_1659),
.B1(n_1641),
.B2(n_1625),
.C1(n_1651),
.C2(n_1539),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1652),
.Y(n_1677)
);

INVxp33_ASAP7_75t_L g1678 ( 
.A(n_1652),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1660),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1662),
.A2(n_1607),
.B1(n_1655),
.B2(n_1538),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1670),
.B(n_1639),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1669),
.B(n_1617),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1663),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1663),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1661),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1666),
.B(n_1655),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1678),
.B(n_1677),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1673),
.Y(n_1688)
);

AOI222xp33_ASAP7_75t_L g1689 ( 
.A1(n_1665),
.A2(n_1602),
.B1(n_1676),
.B2(n_1671),
.C1(n_1666),
.C2(n_1674),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1667),
.B(n_1632),
.Y(n_1690)
);

AOI211x1_ASAP7_75t_L g1691 ( 
.A1(n_1686),
.A2(n_1676),
.B(n_1672),
.C(n_1675),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1680),
.A2(n_1664),
.B1(n_1607),
.B2(n_1538),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_SL g1693 ( 
.A1(n_1689),
.A2(n_1668),
.B(n_1657),
.Y(n_1693)
);

AOI22x1_ASAP7_75t_L g1694 ( 
.A1(n_1679),
.A2(n_1638),
.B1(n_1650),
.B2(n_1643),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1690),
.B(n_1679),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1687),
.Y(n_1696)
);

OAI211xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1680),
.A2(n_1658),
.B(n_1650),
.C(n_1643),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1682),
.A2(n_1607),
.B1(n_1538),
.B2(n_1593),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1683),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1681),
.A2(n_1642),
.B(n_1638),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1696),
.B(n_1690),
.Y(n_1701)
);

OAI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1691),
.A2(n_1684),
.B(n_1685),
.C(n_1688),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1692),
.A2(n_1583),
.B1(n_1607),
.B2(n_1632),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1695),
.B(n_1642),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1694),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1701),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1705),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1704),
.B(n_1699),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1702),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1703),
.B(n_1697),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1701),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1708),
.Y(n_1712)
);

NAND2x1p5_ASAP7_75t_L g1713 ( 
.A(n_1707),
.B(n_1391),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1706),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1709),
.A2(n_1693),
.B1(n_1698),
.B2(n_1700),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1711),
.B(n_1635),
.Y(n_1716)
);

NAND4xp75_ASAP7_75t_L g1717 ( 
.A(n_1712),
.B(n_1710),
.C(n_1658),
.D(n_1626),
.Y(n_1717)
);

XNOR2x1_ASAP7_75t_L g1718 ( 
.A(n_1715),
.B(n_1710),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_SL g1719 ( 
.A(n_1713),
.B(n_1539),
.C(n_1522),
.Y(n_1719)
);

NOR2xp67_ASAP7_75t_L g1720 ( 
.A(n_1719),
.B(n_1714),
.Y(n_1720)
);

A2O1A1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1716),
.B(n_1718),
.C(n_1717),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1593),
.B1(n_1538),
.B2(n_1626),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1721),
.B(n_1615),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1723),
.B(n_1615),
.Y(n_1724)
);

AOI22x1_ASAP7_75t_L g1725 ( 
.A1(n_1722),
.A2(n_1589),
.B1(n_1569),
.B2(n_1570),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1724),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1725),
.Y(n_1727)
);

BUFx2_ASAP7_75t_SL g1728 ( 
.A(n_1726),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1728),
.A2(n_1727),
.B1(n_1593),
.B2(n_1538),
.Y(n_1729)
);

NAND2x1p5_ASAP7_75t_L g1730 ( 
.A(n_1729),
.B(n_1570),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_R g1731 ( 
.A(n_1730),
.B(n_1585),
.C(n_1507),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1589),
.B1(n_1549),
.B2(n_1551),
.C(n_1586),
.Y(n_1732)
);

AOI211xp5_ASAP7_75t_L g1733 ( 
.A1(n_1732),
.A2(n_1447),
.B(n_1551),
.C(n_1549),
.Y(n_1733)
);


endmodule