module real_jpeg_19963_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_57;
wire n_73;
wire n_65;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_52;
wire n_31;
wire n_67;
wire n_58;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_47;
wire n_14;
wire n_11;
wire n_71;
wire n_45;
wire n_25;
wire n_51;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_40;
wire n_36;
wire n_70;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_0),
.A2(n_32),
.B1(n_37),
.B2(n_64),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_1),
.A2(n_17),
.B1(n_20),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_1),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_2),
.A2(n_17),
.B1(n_20),
.B2(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_3),
.A2(n_14),
.B1(n_18),
.B2(n_22),
.Y(n_13)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_32),
.B1(n_37),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_5),
.A2(n_17),
.B1(n_20),
.B2(n_41),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_6),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_21),
.B1(n_32),
.B2(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_17),
.B(n_30),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_28),
.B1(n_32),
.B2(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_15),
.B1(n_46),
.B2(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_62),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_54),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_42),
.B(n_53),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_25),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_25),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_15),
.A2(n_19),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_15),
.A2(n_23),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_17),
.A2(n_20),
.B1(n_29),
.B2(n_30),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_33),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_47),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_35),
.A2(n_38),
.B1(n_40),
.B2(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_48),
.B(n_52),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_73),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_58),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);


endmodule