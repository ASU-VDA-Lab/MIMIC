module fake_ibex_1251_n_6695 (n_151, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_1060, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_1067, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1061, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_1056, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_1051, n_854, n_1008, n_458, n_244, n_73, n_1053, n_343, n_310, n_714, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_1055, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_1025, n_465, n_1057, n_1068, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_1052, n_852, n_789, n_880, n_654, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_1070, n_1074, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_1064, n_1071, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_1066, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1062, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_1072, n_82, n_263, n_1069, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_1063, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_1054, n_44, n_672, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_1049, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_1065, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_1059, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_1073, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_1048, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_1058, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_1050, n_6695);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_1060;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_1067;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1061;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_1056;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_1051;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_1053;
input n_343;
input n_310;
input n_714;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_1055;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_1057;
input n_1068;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_1052;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_1070;
input n_1074;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_1064;
input n_1071;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_1066;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1062;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_1072;
input n_82;
input n_263;
input n_1069;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_1063;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_1054;
input n_44;
input n_672;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_1049;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_1065;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_1059;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_1073;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_1058;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;
input n_1050;

output n_6695;

wire n_4557;
wire n_6210;
wire n_5285;
wire n_6516;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_6537;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_6616;
wire n_4371;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_6567;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_6229;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_6639;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_6658;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_6517;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_6530;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_6602;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_6562;
wire n_3979;
wire n_3714;
wire n_6534;
wire n_6629;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_4854;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_6674;
wire n_6486;
wire n_5261;
wire n_5895;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_1078;
wire n_4422;
wire n_5743;
wire n_1865;
wire n_5033;
wire n_6491;
wire n_4842;
wire n_4786;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_6580;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_6078;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_6625;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_6638;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_6485;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_6114;
wire n_1121;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_6606;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_5252;
wire n_6209;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_6011;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_6533;
wire n_3859;
wire n_6540;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2924;
wire n_2456;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_6691;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6124;
wire n_3352;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_6136;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_5859;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6128;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_6379;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_6570;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_6507;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_3796;
wire n_5719;
wire n_6544;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_6605;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_6527;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_6626;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_6528;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_1095;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_6652;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_6531;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_6502;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_6646;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_3339;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_6595;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_1517;
wire n_5973;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_5770;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_6682;
wire n_2959;
wire n_2420;
wire n_2380;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_6553;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_6543;
wire n_5566;
wire n_6185;
wire n_5342;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_5787;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_5843;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_1278;
wire n_2059;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_6591;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_5824;
wire n_6280;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_6656;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_4919;
wire n_4200;
wire n_4111;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_6637;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_6577;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_6641;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_6556;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_6152;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_6416;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_2266;
wire n_4473;
wire n_6673;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_6482;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_6483;
wire n_4686;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_6598;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6499;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_6594;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_6621;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3919;
wire n_3683;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4962;
wire n_1082;
wire n_4797;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_5384;
wire n_6550;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5265;
wire n_5087;
wire n_4401;
wire n_4727;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_6176;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6662;
wire n_6461;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_6617;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_6549;
wire n_5097;
wire n_4688;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_6607;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_6564;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_6566;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_6496;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5319;
wire n_5543;
wire n_4721;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_5631;
wire n_5983;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_6021;
wire n_3221;
wire n_3210;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_4067;
wire n_4997;
wire n_5906;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_5916;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_6476;
wire n_5828;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_6669;
wire n_5357;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_1709;
wire n_6655;
wire n_6541;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_6497;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_6535;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6676;
wire n_6117;
wire n_6563;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_6448;
wire n_3684;
wire n_6667;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_6552;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2573;
wire n_1793;
wire n_2424;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_6653;
wire n_3098;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_6539;
wire n_4330;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_6560;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_6519;
wire n_3703;
wire n_5116;
wire n_6635;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_6661;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_1593;
wire n_1775;
wire n_6361;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_6523;
wire n_5746;
wire n_5883;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_6062;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_6252;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_2463;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_6630;
wire n_6631;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_6489;
wire n_1251;
wire n_6657;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_6481;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_6694;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_6597;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_6647;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4924;
wire n_2238;
wire n_6398;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_1294;
wire n_1351;
wire n_6679;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_6660;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_5096;
wire n_6480;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_6693;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_6615;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5862;
wire n_5869;
wire n_1238;
wire n_3959;
wire n_4288;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_5277;
wire n_5900;
wire n_3647;
wire n_6240;
wire n_3928;
wire n_3619;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_6498;
wire n_1669;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_6574;
wire n_2756;
wire n_1175;
wire n_4408;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_5645;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_6139;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_6494;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_6380;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_6526;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_6520;
wire n_4906;
wire n_4257;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_6444;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_6648;
wire n_2408;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_6622;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_6488;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_6692;
wire n_6590;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_6501;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_6551;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_5644;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_5700;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_6579;
wire n_4018;
wire n_2609;
wire n_6633;
wire n_4613;
wire n_5940;
wire n_6614;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_3261;
wire n_5324;
wire n_6547;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_6589;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_6583;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_6310;
wire n_1506;
wire n_5061;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_6618;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_6249;
wire n_3559;
wire n_5184;
wire n_6440;
wire n_5747;
wire n_6575;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_6584;
wire n_6689;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_6643;
wire n_6569;
wire n_3132;
wire n_5618;
wire n_6596;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_5464;
wire n_6548;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_2565;
wire n_4201;
wire n_6634;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_6478;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_6056;
wire n_2873;
wire n_1576;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_6375;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_6025;
wire n_6168;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_2275;
wire n_1853;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_6525;
wire n_1764;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_6675;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_5123;
wire n_6160;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_6678;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_6561;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_6557;
wire n_2748;
wire n_5359;
wire n_6503;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5999;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_6140;
wire n_5903;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_6663;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_6620;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_6529;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_6554;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_6585;
wire n_5985;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_6473;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_6651;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_6490;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_6558;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_6500;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_6518;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_6578;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_6049;
wire n_2419;
wire n_6671;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_5724;
wire n_6610;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_6576;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_6260;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_6624;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_6687;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_6088;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_4163;
wire n_2831;
wire n_6504;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_1587;
wire n_2555;
wire n_6356;
wire n_6640;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_6521;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_6582;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_6623;
wire n_1880;
wire n_6225;
wire n_1642;
wire n_5744;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6493;
wire n_6364;
wire n_5715;
wire n_6665;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_6649;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_2157;
wire n_6546;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_6555;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_6532;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_6677;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_6524;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_6514;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_6685;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_6609;
wire n_5853;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_6627;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_6162;
wire n_5592;
wire n_5484;
wire n_6650;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_6592;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_6512;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_6522;
wire n_4907;
wire n_4659;
wire n_2128;
wire n_1697;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_6613;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_6538;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_6505;
wire n_3989;
wire n_6581;
wire n_5565;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_6484;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_6573;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_5500;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_6568;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6167;
wire n_6189;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_6611;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_6588;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5984;
wire n_6385;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_6586;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_6479;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_2374;
wire n_1614;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6612;
wire n_6376;
wire n_2571;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_6132;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6089;
wire n_5211;
wire n_1668;
wire n_5861;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6175;
wire n_5279;
wire n_6506;
wire n_6690;
wire n_4650;
wire n_6415;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_6644;
wire n_1588;
wire n_2579;
wire n_6688;
wire n_2876;
wire n_6670;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_6680;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_6046;
wire n_4981;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_6329;
wire n_4755;
wire n_6355;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_1106;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1985;
wire n_1140;
wire n_4740;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_6632;
wire n_2717;
wire n_1589;
wire n_5720;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_6654;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_6672;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_5682;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1566;
wire n_1464;
wire n_6565;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_6601;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_3331;
wire n_2999;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6513;
wire n_6214;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_6559;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_6683;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5819;
wire n_5855;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6608;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_6593;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_6542;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_5604;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_6515;
wire n_6619;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_6664;
wire n_5992;
wire n_5105;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_6599;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_6099;
wire n_5939;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_3747;
wire n_1323;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1458;
wire n_1694;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_5780;
wire n_2642;
wire n_5485;
wire n_5737;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_6571;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_6509;
wire n_6642;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_6636;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_6492;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_6545;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_6250;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_1167;
wire n_3231;
wire n_6423;
wire n_6659;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6668;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_2345;
wire n_1139;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_6510;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_6353;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_6686;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_1088;
wire n_6666;
wire n_6075;
wire n_1102;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_6317;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_1542;
wire n_1547;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_6511;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_6603;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_6587;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_6487;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_6495;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_6194;
wire n_1911;
wire n_6381;
wire n_2870;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_6628;
wire n_5283;
wire n_1419;
wire n_4738;
wire n_6604;
wire n_1193;
wire n_3557;
wire n_2928;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_2668;
wire n_6684;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_6261;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_6645;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_6572;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_6508;
wire n_6536;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_6681;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_6600;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_248),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_116),
.Y(n_1076)
);

CKINVDCx16_ASAP7_75t_R g1077 ( 
.A(n_820),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_461),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_4),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_940),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_422),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_325),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_387),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_576),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_395),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_83),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_716),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_1009),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_21),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_814),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_620),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_125),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_474),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_939),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_340),
.Y(n_1095)
);

BUFx5_ASAP7_75t_L g1096 ( 
.A(n_1008),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_363),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_24),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_384),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_558),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_992),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1023),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_781),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_607),
.Y(n_1104)
);

BUFx10_ASAP7_75t_L g1105 ( 
.A(n_111),
.Y(n_1105)
);

BUFx10_ASAP7_75t_L g1106 ( 
.A(n_231),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_826),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_865),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_325),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1039),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_102),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_198),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_752),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_963),
.Y(n_1114)
);

BUFx10_ASAP7_75t_L g1115 ( 
.A(n_314),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_497),
.Y(n_1116)
);

CKINVDCx14_ASAP7_75t_R g1117 ( 
.A(n_302),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_103),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_231),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_77),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_919),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_550),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_486),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_663),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_789),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_255),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_207),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_57),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_304),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_652),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_649),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_713),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_683),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_921),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_782),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_236),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_784),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_792),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_669),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1021),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1029),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_770),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_574),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1035),
.Y(n_1144)
);

BUFx10_ASAP7_75t_L g1145 ( 
.A(n_991),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_905),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_57),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_136),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_599),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_832),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1015),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1010),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_721),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_786),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_432),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_551),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1036),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_419),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_415),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_78),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_435),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1028),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_715),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_701),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_752),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_661),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_147),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_597),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_987),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_797),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_109),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_341),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_112),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_386),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_440),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_650),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_404),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_949),
.Y(n_1178)
);

BUFx5_ASAP7_75t_L g1179 ( 
.A(n_763),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_149),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_460),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_187),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_965),
.Y(n_1183)
);

CKINVDCx16_ASAP7_75t_R g1184 ( 
.A(n_854),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_294),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_181),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_101),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_591),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_988),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_285),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1024),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_699),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1037),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_192),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_56),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_595),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_5),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_209),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_652),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_974),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_137),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_33),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_756),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_138),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_993),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_547),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_251),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_105),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1010),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_104),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_320),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_510),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_973),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_490),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_877),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_79),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_594),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_943),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_982),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_325),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_305),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_694),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1043),
.Y(n_1223)
);

BUFx5_ASAP7_75t_L g1224 ( 
.A(n_908),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_601),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_700),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_989),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_255),
.Y(n_1228)
);

CKINVDCx16_ASAP7_75t_R g1229 ( 
.A(n_1032),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1039),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_255),
.Y(n_1231)
);

CKINVDCx16_ASAP7_75t_R g1232 ( 
.A(n_181),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_718),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_799),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_645),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_550),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_289),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_160),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_745),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_500),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1030),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_812),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_973),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_362),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_575),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1073),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_42),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_676),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_762),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_486),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_876),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1033),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_753),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_783),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1036),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_247),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1006),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_156),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_57),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_246),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_456),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_948),
.Y(n_1262)
);

INVxp33_ASAP7_75t_L g1263 ( 
.A(n_302),
.Y(n_1263)
);

BUFx2_ASAP7_75t_SL g1264 ( 
.A(n_1017),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_235),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_578),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_576),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_561),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_616),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_283),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_176),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_940),
.Y(n_1272)
);

BUFx10_ASAP7_75t_L g1273 ( 
.A(n_15),
.Y(n_1273)
);

CKINVDCx16_ASAP7_75t_R g1274 ( 
.A(n_203),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_763),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1031),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1008),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_60),
.Y(n_1278)
);

BUFx8_ASAP7_75t_SL g1279 ( 
.A(n_1016),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_281),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_324),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_181),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1025),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_464),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1003),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_328),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_445),
.Y(n_1287)
);

BUFx8_ASAP7_75t_SL g1288 ( 
.A(n_775),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_518),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1026),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_326),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_444),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_404),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_291),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_200),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_59),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_534),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1049),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_679),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1016),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_919),
.Y(n_1301)
);

BUFx8_ASAP7_75t_SL g1302 ( 
.A(n_277),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1051),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_997),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_337),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_980),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_696),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_164),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_731),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_398),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_680),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_232),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_518),
.Y(n_1313)
);

BUFx10_ASAP7_75t_L g1314 ( 
.A(n_371),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_433),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_872),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_412),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_953),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_958),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1044),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_619),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_969),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_855),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_815),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_975),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_632),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_303),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_380),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_238),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_623),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_745),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_90),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_294),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_208),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1073),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_380),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_672),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_437),
.Y(n_1338)
);

BUFx5_ASAP7_75t_L g1339 ( 
.A(n_673),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_962),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_995),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_974),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_738),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_713),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_503),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_688),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_352),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_121),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_505),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_243),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_572),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_357),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_909),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_100),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1014),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_715),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1002),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_312),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_302),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1070),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1024),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_526),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_936),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_348),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_34),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_326),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_978),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_534),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_675),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1013),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_806),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_516),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_982),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_456),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_64),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_424),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_426),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_756),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_456),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_986),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_486),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_956),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_854),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_648),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_610),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_239),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_318),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_645),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1058),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_167),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_627),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_299),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_216),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1041),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_509),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_506),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_330),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_258),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_304),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_351),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_871),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_284),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_448),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_996),
.Y(n_1404)
);

BUFx5_ASAP7_75t_L g1405 ( 
.A(n_158),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_397),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_264),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_526),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_980),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_803),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_869),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_517),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_588),
.Y(n_1413)
);

BUFx8_ASAP7_75t_SL g1414 ( 
.A(n_705),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_395),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1007),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_339),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1037),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_953),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_638),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_985),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_406),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1050),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_60),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_296),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1012),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_130),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_942),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_789),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_407),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_260),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_917),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_398),
.Y(n_1433)
);

INVxp67_ASAP7_75t_L g1434 ( 
.A(n_1052),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_480),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1046),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1053),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_171),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1020),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_28),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_153),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_403),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_381),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_213),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_996),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1043),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_412),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_834),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_79),
.Y(n_1449)
);

CKINVDCx14_ASAP7_75t_R g1450 ( 
.A(n_169),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_1047),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_595),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_338),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_206),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_329),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_516),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_377),
.Y(n_1457)
);

BUFx5_ASAP7_75t_L g1458 ( 
.A(n_78),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_548),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_734),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_333),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_72),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_806),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_565),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_71),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_800),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_13),
.Y(n_1467)
);

BUFx2_ASAP7_75t_SL g1468 ( 
.A(n_895),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_352),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_226),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_999),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_27),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_928),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_417),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_676),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_53),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_123),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_469),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_310),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_508),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_211),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_639),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_48),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_69),
.Y(n_1484)
);

BUFx10_ASAP7_75t_L g1485 ( 
.A(n_341),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_491),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_864),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_102),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1009),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_284),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_331),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_713),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_378),
.Y(n_1493)
);

CKINVDCx16_ASAP7_75t_R g1494 ( 
.A(n_41),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1027),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_336),
.Y(n_1496)
);

BUFx5_ASAP7_75t_L g1497 ( 
.A(n_166),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_494),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_371),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_699),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_990),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_628),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1049),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1003),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_866),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1034),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1049),
.Y(n_1507)
);

BUFx5_ASAP7_75t_L g1508 ( 
.A(n_171),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_743),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_880),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_512),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_643),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_29),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1004),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_983),
.Y(n_1515)
);

INVxp67_ASAP7_75t_SL g1516 ( 
.A(n_417),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_51),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_588),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_642),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_14),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_662),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_551),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_706),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_110),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_17),
.Y(n_1525)
);

CKINVDCx14_ASAP7_75t_R g1526 ( 
.A(n_794),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_140),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_722),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_881),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_400),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_408),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_501),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_455),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1005),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_114),
.Y(n_1535)
);

CKINVDCx16_ASAP7_75t_R g1536 ( 
.A(n_1031),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_875),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_421),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_712),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_8),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_27),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_526),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_783),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_338),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_608),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_133),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_361),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_143),
.Y(n_1548)
);

BUFx10_ASAP7_75t_L g1549 ( 
.A(n_769),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_293),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_93),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_225),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1054),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_284),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_357),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_939),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1040),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_911),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_939),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_768),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_761),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_105),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1009),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_96),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1035),
.Y(n_1565)
);

CKINVDCx16_ASAP7_75t_R g1566 ( 
.A(n_981),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_17),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_812),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1053),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_758),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_9),
.Y(n_1571)
);

BUFx5_ASAP7_75t_L g1572 ( 
.A(n_1003),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_340),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_545),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_967),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_853),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1011),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_812),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_669),
.Y(n_1579)
);

CKINVDCx20_ASAP7_75t_R g1580 ( 
.A(n_598),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_849),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_462),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_422),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1007),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_64),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_984),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1069),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_663),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_605),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_502),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_479),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_480),
.Y(n_1592)
);

CKINVDCx14_ASAP7_75t_R g1593 ( 
.A(n_470),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_954),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_226),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_742),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1001),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_505),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_129),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1030),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_421),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_310),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_940),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_761),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_863),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_924),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1028),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_979),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_172),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_553),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_674),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_767),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_694),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_349),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_25),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_399),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_744),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1002),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_474),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_144),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_899),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_48),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_725),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_983),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1027),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_369),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_80),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1042),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1038),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_994),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_166),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_510),
.Y(n_1632)
);

BUFx5_ASAP7_75t_L g1633 ( 
.A(n_942),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_162),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_299),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1018),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_261),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_84),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1019),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_241),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_510),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_88),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_327),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_778),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_132),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_966),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_792),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_768),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1022),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_490),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_947),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_496),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_492),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_188),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_254),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_554),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1053),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_424),
.Y(n_1658)
);

CKINVDCx16_ASAP7_75t_R g1659 ( 
.A(n_995),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_738),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_539),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_421),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_153),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_164),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_881),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_222),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_120),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_703),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_395),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_614),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_894),
.Y(n_1671)
);

CKINVDCx16_ASAP7_75t_R g1672 ( 
.A(n_58),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_924),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_995),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_313),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_878),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_615),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_677),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_631),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1031),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_761),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_766),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_998),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_986),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1045),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_854),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_707),
.Y(n_1687)
);

CKINVDCx16_ASAP7_75t_R g1688 ( 
.A(n_1048),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_563),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_973),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1000),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_440),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_569),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_266),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_717),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1064),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_542),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_276),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_901),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_844),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_210),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1043),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1273),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_1117),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1273),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1472),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1273),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1259),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1567),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1120),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1494),
.Y(n_1711)
);

INVxp67_ASAP7_75t_SL g1712 ( 
.A(n_1098),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1672),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1117),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1197),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1450),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1216),
.Y(n_1717)
);

INVxp67_ASAP7_75t_SL g1718 ( 
.A(n_1098),
.Y(n_1718)
);

CKINVDCx14_ASAP7_75t_R g1719 ( 
.A(n_1450),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1195),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1526),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1458),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1484),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1526),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1279),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1517),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1540),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_1279),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1615),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1585),
.Y(n_1730)
);

CKINVDCx16_ASAP7_75t_R g1731 ( 
.A(n_1077),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1182),
.Y(n_1732)
);

INVxp33_ASAP7_75t_L g1733 ( 
.A(n_1091),
.Y(n_1733)
);

INVxp67_ASAP7_75t_SL g1734 ( 
.A(n_1195),
.Y(n_1734)
);

INVxp67_ASAP7_75t_SL g1735 ( 
.A(n_1296),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1222),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1593),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_1288),
.Y(n_1738)
);

CKINVDCx16_ASAP7_75t_R g1739 ( 
.A(n_1184),
.Y(n_1739)
);

INVxp67_ASAP7_75t_SL g1740 ( 
.A(n_1296),
.Y(n_1740)
);

INVxp33_ASAP7_75t_SL g1741 ( 
.A(n_1108),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1329),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1593),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1348),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1251),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1376),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1076),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1137),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1394),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_1288),
.Y(n_1750)
);

NOR2xp67_ASAP7_75t_L g1751 ( 
.A(n_1457),
.B(n_0),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1417),
.Y(n_1752)
);

INVxp33_ASAP7_75t_L g1753 ( 
.A(n_1312),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1655),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1699),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1302),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1272),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1294),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1590),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1263),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1601),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1457),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1302),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1489),
.Y(n_1764)
);

CKINVDCx20_ASAP7_75t_R g1765 ( 
.A(n_1414),
.Y(n_1765)
);

INVxp67_ASAP7_75t_SL g1766 ( 
.A(n_1263),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1147),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1694),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1458),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1458),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1414),
.Y(n_1771)
);

INVxp33_ASAP7_75t_SL g1772 ( 
.A(n_1079),
.Y(n_1772)
);

INVxp67_ASAP7_75t_SL g1773 ( 
.A(n_1424),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1089),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1458),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1458),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1458),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1202),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1458),
.Y(n_1779)
);

CKINVDCx20_ASAP7_75t_R g1780 ( 
.A(n_1160),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1100),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1101),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1109),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1112),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1113),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1247),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1116),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1125),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1278),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1127),
.Y(n_1790)
);

CKINVDCx16_ASAP7_75t_R g1791 ( 
.A(n_1229),
.Y(n_1791)
);

INVxp33_ASAP7_75t_L g1792 ( 
.A(n_1128),
.Y(n_1792)
);

CKINVDCx14_ASAP7_75t_R g1793 ( 
.A(n_1105),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1375),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1132),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1136),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1141),
.Y(n_1797)
);

CKINVDCx14_ASAP7_75t_R g1798 ( 
.A(n_1105),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1365),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1424),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1142),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1143),
.Y(n_1802)
);

CKINVDCx20_ASAP7_75t_R g1803 ( 
.A(n_1462),
.Y(n_1803)
);

INVxp67_ASAP7_75t_SL g1804 ( 
.A(n_1082),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1144),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1148),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1232),
.B(n_0),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1153),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1158),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1161),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1164),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1274),
.B(n_1451),
.Y(n_1812)
);

INVxp33_ASAP7_75t_L g1813 ( 
.A(n_1128),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1181),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1096),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1190),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1082),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1440),
.Y(n_1818)
);

CKINVDCx20_ASAP7_75t_R g1819 ( 
.A(n_1622),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1192),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1193),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1096),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1204),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1207),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1096),
.Y(n_1825)
);

INVxp33_ASAP7_75t_SL g1826 ( 
.A(n_1449),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1209),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1212),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1214),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1223),
.Y(n_1830)
);

INVxp33_ASAP7_75t_SL g1831 ( 
.A(n_1465),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1467),
.Y(n_1832)
);

INVxp67_ASAP7_75t_SL g1833 ( 
.A(n_1122),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1225),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1228),
.Y(n_1835)
);

BUFx3_ASAP7_75t_L g1836 ( 
.A(n_1799),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1767),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1730),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1760),
.B(n_1105),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1743),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1722),
.Y(n_1841)
);

BUFx12f_ASAP7_75t_L g1842 ( 
.A(n_1713),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1760),
.B(n_1476),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1710),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1766),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1815),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1715),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1770),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1717),
.Y(n_1849)
);

BUFx12f_ASAP7_75t_L g1850 ( 
.A(n_1756),
.Y(n_1850)
);

CKINVDCx6p67_ASAP7_75t_R g1851 ( 
.A(n_1731),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1723),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_L g1853 ( 
.A(n_1726),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1822),
.Y(n_1854)
);

OA21x2_ASAP7_75t_L g1855 ( 
.A1(n_1769),
.A2(n_1121),
.B(n_1093),
.Y(n_1855)
);

BUFx6f_ASAP7_75t_L g1856 ( 
.A(n_1727),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1729),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1793),
.Y(n_1858)
);

INVx5_ASAP7_75t_L g1859 ( 
.A(n_1757),
.Y(n_1859)
);

BUFx3_ASAP7_75t_L g1860 ( 
.A(n_1832),
.Y(n_1860)
);

CKINVDCx16_ASAP7_75t_R g1861 ( 
.A(n_1798),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1766),
.B(n_1106),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1708),
.B(n_1106),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1733),
.B(n_1106),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1712),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1825),
.A2(n_1121),
.B(n_1093),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1712),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1716),
.B(n_1513),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1721),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1734),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1762),
.Y(n_1871)
);

OAI22x1_ASAP7_75t_SL g1872 ( 
.A1(n_1780),
.A2(n_1803),
.B1(n_1819),
.B2(n_1794),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1720),
.B(n_1774),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1734),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1772),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1735),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1778),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1732),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1736),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1735),
.Y(n_1880)
);

INVx2_ASAP7_75t_SL g1881 ( 
.A(n_1786),
.Y(n_1881)
);

OAI22x1_ASAP7_75t_SL g1882 ( 
.A1(n_1725),
.A2(n_1386),
.B1(n_1111),
.B2(n_1149),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1711),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1742),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1826),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1747),
.B(n_1122),
.Y(n_1886)
);

BUFx12f_ASAP7_75t_L g1887 ( 
.A(n_1763),
.Y(n_1887)
);

OA21x2_ASAP7_75t_L g1888 ( 
.A1(n_1775),
.A2(n_1777),
.B(n_1776),
.Y(n_1888)
);

BUFx6f_ASAP7_75t_L g1889 ( 
.A(n_1744),
.Y(n_1889)
);

INVx5_ASAP7_75t_L g1890 ( 
.A(n_1739),
.Y(n_1890)
);

OAI21x1_ASAP7_75t_L g1891 ( 
.A1(n_1779),
.A2(n_1156),
.B(n_1154),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1720),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1746),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1749),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1812),
.A2(n_1525),
.B1(n_1541),
.B2(n_1520),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1789),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1706),
.Y(n_1897)
);

OA21x2_ASAP7_75t_L g1898 ( 
.A1(n_1740),
.A2(n_1156),
.B(n_1154),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1740),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1833),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1747),
.B(n_1748),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1752),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1833),
.Y(n_1903)
);

BUFx12f_ASAP7_75t_L g1904 ( 
.A(n_1818),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1831),
.Y(n_1905)
);

AND2x4_ASAP7_75t_L g1906 ( 
.A(n_1748),
.B(n_1758),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1754),
.Y(n_1907)
);

AND2x6_ASAP7_75t_L g1908 ( 
.A(n_1703),
.B(n_1129),
.Y(n_1908)
);

INVx5_ASAP7_75t_L g1909 ( 
.A(n_1791),
.Y(n_1909)
);

INVx5_ASAP7_75t_L g1910 ( 
.A(n_1751),
.Y(n_1910)
);

INVx5_ASAP7_75t_L g1911 ( 
.A(n_1753),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1755),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1817),
.B(n_1571),
.Y(n_1913)
);

INVx5_ASAP7_75t_L g1914 ( 
.A(n_1741),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1759),
.B(n_1761),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1705),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_L g1917 ( 
.A1(n_1707),
.A2(n_1782),
.B(n_1781),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1783),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1745),
.Y(n_1919)
);

INVx6_ASAP7_75t_L g1920 ( 
.A(n_1719),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1764),
.B(n_1129),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1709),
.B(n_1115),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1817),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1784),
.Y(n_1924)
);

AND2x6_ASAP7_75t_L g1925 ( 
.A(n_1768),
.B(n_1155),
.Y(n_1925)
);

BUFx8_ASAP7_75t_L g1926 ( 
.A(n_1728),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1718),
.B(n_1627),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1704),
.B(n_1155),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1785),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1773),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1787),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1773),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1714),
.B(n_1176),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1724),
.A2(n_1536),
.B1(n_1659),
.B2(n_1566),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1788),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1737),
.B(n_1804),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1800),
.B(n_1688),
.Y(n_1937)
);

OAI21x1_ASAP7_75t_L g1938 ( 
.A1(n_1790),
.A2(n_1185),
.B(n_1169),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1800),
.B(n_1075),
.Y(n_1939)
);

INVxp67_ASAP7_75t_L g1940 ( 
.A(n_1807),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1795),
.Y(n_1941)
);

BUFx6f_ASAP7_75t_L g1942 ( 
.A(n_1796),
.Y(n_1942)
);

INVxp67_ASAP7_75t_L g1943 ( 
.A(n_1835),
.Y(n_1943)
);

CKINVDCx16_ASAP7_75t_R g1944 ( 
.A(n_1738),
.Y(n_1944)
);

CKINVDCx20_ASAP7_75t_R g1945 ( 
.A(n_1750),
.Y(n_1945)
);

INVx5_ASAP7_75t_L g1946 ( 
.A(n_1792),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1797),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1801),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1802),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1805),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1806),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1808),
.B(n_1115),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1809),
.Y(n_1953)
);

INVxp67_ASAP7_75t_L g1954 ( 
.A(n_1810),
.Y(n_1954)
);

INVx5_ASAP7_75t_L g1955 ( 
.A(n_1813),
.Y(n_1955)
);

CKINVDCx16_ASAP7_75t_R g1956 ( 
.A(n_1765),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1811),
.Y(n_1957)
);

AOI22x1_ASAP7_75t_SL g1958 ( 
.A1(n_1771),
.A2(n_1386),
.B1(n_1150),
.B2(n_1196),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1814),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1816),
.B(n_1078),
.Y(n_1960)
);

BUFx3_ASAP7_75t_L g1961 ( 
.A(n_1820),
.Y(n_1961)
);

OAI22x1_ASAP7_75t_SL g1962 ( 
.A1(n_1821),
.A2(n_1198),
.B1(n_1203),
.B2(n_1095),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1823),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1824),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1827),
.A2(n_1081),
.B1(n_1084),
.B2(n_1083),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1828),
.Y(n_1966)
);

BUFx8_ASAP7_75t_SL g1967 ( 
.A(n_1829),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1830),
.B(n_1115),
.Y(n_1968)
);

BUFx12f_ASAP7_75t_L g1969 ( 
.A(n_1834),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1710),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1767),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1767),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1793),
.Y(n_1973)
);

INVx5_ASAP7_75t_L g1974 ( 
.A(n_1757),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1722),
.Y(n_1975)
);

INVx5_ASAP7_75t_L g1976 ( 
.A(n_1757),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1722),
.Y(n_1977)
);

BUFx2_ASAP7_75t_L g1978 ( 
.A(n_1767),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1722),
.Y(n_1979)
);

BUFx2_ASAP7_75t_L g1980 ( 
.A(n_1767),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1767),
.Y(n_1981)
);

INVx6_ASAP7_75t_L g1982 ( 
.A(n_1731),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1799),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1710),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1760),
.B(n_1085),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1722),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1760),
.B(n_1176),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1760),
.B(n_1325),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1710),
.Y(n_1989)
);

CKINVDCx16_ASAP7_75t_R g1990 ( 
.A(n_1793),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1760),
.B(n_1325),
.Y(n_1991)
);

BUFx6f_ASAP7_75t_L g1992 ( 
.A(n_1710),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1722),
.Y(n_1993)
);

BUFx12f_ASAP7_75t_L g1994 ( 
.A(n_1713),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1710),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_L g1996 ( 
.A1(n_1710),
.A2(n_1185),
.B(n_1169),
.Y(n_1996)
);

BUFx8_ASAP7_75t_SL g1997 ( 
.A(n_1725),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1710),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1722),
.Y(n_1999)
);

BUFx2_ASAP7_75t_L g2000 ( 
.A(n_1767),
.Y(n_2000)
);

BUFx12f_ASAP7_75t_L g2001 ( 
.A(n_1713),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1710),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1716),
.B(n_1221),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1767),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1760),
.B(n_1086),
.Y(n_2005)
);

INVx5_ASAP7_75t_L g2006 ( 
.A(n_1757),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1760),
.Y(n_2007)
);

BUFx8_ASAP7_75t_SL g2008 ( 
.A(n_1725),
.Y(n_2008)
);

INVx3_ASAP7_75t_L g2009 ( 
.A(n_1767),
.Y(n_2009)
);

BUFx8_ASAP7_75t_SL g2010 ( 
.A(n_1725),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1799),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1710),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1722),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1767),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1767),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_1760),
.B(n_1336),
.Y(n_2016)
);

CKINVDCx20_ASAP7_75t_R g2017 ( 
.A(n_1780),
.Y(n_2017)
);

INVx5_ASAP7_75t_L g2018 ( 
.A(n_1757),
.Y(n_2018)
);

INVx3_ASAP7_75t_L g2019 ( 
.A(n_1767),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1760),
.B(n_1145),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1760),
.B(n_1145),
.Y(n_2021)
);

BUFx12f_ASAP7_75t_L g2022 ( 
.A(n_1713),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1741),
.A2(n_1087),
.B1(n_1090),
.B2(n_1088),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1722),
.Y(n_2024)
);

INVx3_ASAP7_75t_L g2025 ( 
.A(n_1767),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1767),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1760),
.B(n_1145),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1760),
.Y(n_2028)
);

INVx5_ASAP7_75t_L g2029 ( 
.A(n_1757),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1722),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_1760),
.B(n_1336),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1760),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1716),
.B(n_1313),
.Y(n_2033)
);

BUFx6f_ASAP7_75t_L g2034 ( 
.A(n_1710),
.Y(n_2034)
);

BUFx6f_ASAP7_75t_L g2035 ( 
.A(n_1710),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1760),
.B(n_1092),
.Y(n_2036)
);

AND2x6_ASAP7_75t_L g2037 ( 
.A(n_1703),
.B(n_1353),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1760),
.B(n_1250),
.Y(n_2038)
);

BUFx8_ASAP7_75t_L g2039 ( 
.A(n_1713),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_1710),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1710),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1793),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1722),
.Y(n_2043)
);

BUFx2_ASAP7_75t_L g2044 ( 
.A(n_1767),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1722),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1760),
.Y(n_2046)
);

BUFx12f_ASAP7_75t_L g2047 ( 
.A(n_1713),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1722),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1760),
.B(n_1353),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1815),
.Y(n_2050)
);

AND2x4_ASAP7_75t_L g2051 ( 
.A(n_1760),
.B(n_1370),
.Y(n_2051)
);

BUFx12f_ASAP7_75t_L g2052 ( 
.A(n_1713),
.Y(n_2052)
);

INVx5_ASAP7_75t_L g2053 ( 
.A(n_1757),
.Y(n_2053)
);

INVx4_ASAP7_75t_L g2054 ( 
.A(n_1743),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_1767),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1710),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1722),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1716),
.B(n_1434),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1722),
.Y(n_2059)
);

INVx4_ASAP7_75t_L g2060 ( 
.A(n_1743),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1952),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1837),
.B(n_1250),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1952),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1968),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1938),
.Y(n_2065)
);

INVxp67_ASAP7_75t_L g2066 ( 
.A(n_1971),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1855),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1837),
.B(n_1978),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1996),
.Y(n_2069)
);

INVxp67_ASAP7_75t_L g2070 ( 
.A(n_1972),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1968),
.Y(n_2071)
);

AND2x4_ASAP7_75t_L g2072 ( 
.A(n_1981),
.B(n_1516),
.Y(n_2072)
);

NOR3xp33_ASAP7_75t_L g2073 ( 
.A(n_1978),
.B(n_1146),
.C(n_1080),
.Y(n_2073)
);

OR2x6_ASAP7_75t_L g2074 ( 
.A(n_1980),
.B(n_1264),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1980),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1932),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_2000),
.Y(n_2077)
);

HB1xp67_ASAP7_75t_L g2078 ( 
.A(n_2004),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1932),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_2000),
.Y(n_2080)
);

INVx3_ASAP7_75t_L g2081 ( 
.A(n_2009),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_2044),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_2044),
.Y(n_2083)
);

NAND2xp33_ASAP7_75t_SL g2084 ( 
.A(n_2014),
.B(n_1094),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1839),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1839),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_2015),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_R g2088 ( 
.A(n_1858),
.B(n_1261),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_2055),
.Y(n_2089)
);

BUFx6f_ASAP7_75t_L g2090 ( 
.A(n_1855),
.Y(n_2090)
);

BUFx6f_ASAP7_75t_L g2091 ( 
.A(n_1866),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1891),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1913),
.B(n_1483),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_2019),
.B(n_1370),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1943),
.B(n_1950),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1898),
.Y(n_2096)
);

BUFx6f_ASAP7_75t_L g2097 ( 
.A(n_2025),
.Y(n_2097)
);

BUFx6f_ASAP7_75t_L g2098 ( 
.A(n_2026),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1862),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1954),
.B(n_1096),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1862),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2020),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1898),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1861),
.Y(n_2104)
);

CKINVDCx20_ASAP7_75t_R g2105 ( 
.A(n_2017),
.Y(n_2105)
);

INVx4_ASAP7_75t_L g2106 ( 
.A(n_1969),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1844),
.Y(n_2107)
);

INVx3_ASAP7_75t_L g2108 ( 
.A(n_1836),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1990),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2020),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1864),
.B(n_1250),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_2054),
.B(n_1097),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_1911),
.Y(n_2113)
);

INVx3_ASAP7_75t_L g2114 ( 
.A(n_1860),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2021),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_2039),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2021),
.Y(n_2117)
);

CKINVDCx20_ASAP7_75t_R g2118 ( 
.A(n_1875),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2027),
.Y(n_2119)
);

CKINVDCx20_ASAP7_75t_R g2120 ( 
.A(n_1885),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2027),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_1911),
.Y(n_2122)
);

AND3x2_ASAP7_75t_L g2123 ( 
.A(n_1896),
.B(n_1410),
.C(n_1293),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_1905),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2038),
.Y(n_2125)
);

AND2x6_ASAP7_75t_L g2126 ( 
.A(n_1922),
.B(n_1482),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1851),
.Y(n_2127)
);

NAND2xp33_ASAP7_75t_R g2128 ( 
.A(n_1973),
.B(n_1099),
.Y(n_2128)
);

INVxp67_ASAP7_75t_L g2129 ( 
.A(n_1883),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_1997),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_1983),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2038),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1864),
.B(n_1314),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1930),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1893),
.Y(n_2135)
);

BUFx2_ASAP7_75t_L g2136 ( 
.A(n_2011),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1907),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1912),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1879),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1838),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1922),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_2008),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_2010),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1878),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1863),
.B(n_1314),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1844),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1884),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1879),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1843),
.B(n_1096),
.Y(n_2149)
);

AND2x6_ASAP7_75t_L g2150 ( 
.A(n_1863),
.B(n_1482),
.Y(n_2150)
);

BUFx6f_ASAP7_75t_L g2151 ( 
.A(n_1888),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1847),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_1872),
.Y(n_2153)
);

NOR2xp67_ASAP7_75t_L g2154 ( 
.A(n_1890),
.B(n_0),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1847),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1892),
.B(n_1096),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_2042),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1927),
.B(n_1096),
.Y(n_2158)
);

BUFx6f_ASAP7_75t_L g2159 ( 
.A(n_1888),
.Y(n_2159)
);

CKINVDCx20_ASAP7_75t_R g2160 ( 
.A(n_1896),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1873),
.B(n_1179),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1842),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_L g2163 ( 
.A(n_1917),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_L g2164 ( 
.A(n_1953),
.B(n_1179),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1849),
.Y(n_2165)
);

CKINVDCx5p33_ASAP7_75t_R g2166 ( 
.A(n_1994),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1889),
.Y(n_2167)
);

HB1xp67_ASAP7_75t_L g2168 ( 
.A(n_1919),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1849),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_2001),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1889),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1923),
.B(n_1179),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_2022),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_1897),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1894),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1894),
.Y(n_2176)
);

CKINVDCx20_ASAP7_75t_R g2177 ( 
.A(n_1945),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1902),
.Y(n_2178)
);

AND2x4_ASAP7_75t_L g2179 ( 
.A(n_1886),
.B(n_1584),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1902),
.Y(n_2180)
);

BUFx10_ASAP7_75t_L g2181 ( 
.A(n_1982),
.Y(n_2181)
);

INVxp67_ASAP7_75t_L g2182 ( 
.A(n_1901),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1852),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_2047),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1871),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_2052),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_1904),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_1845),
.B(n_1584),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1939),
.B(n_1179),
.Y(n_2189)
);

CKINVDCx5p33_ASAP7_75t_R g2190 ( 
.A(n_1850),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_1887),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1926),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1961),
.Y(n_2193)
);

BUFx10_ASAP7_75t_L g2194 ( 
.A(n_1982),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1852),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1865),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1853),
.Y(n_2197)
);

BUFx3_ASAP7_75t_L g2198 ( 
.A(n_1920),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_1877),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_1944),
.Y(n_2200)
);

CKINVDCx20_ASAP7_75t_R g2201 ( 
.A(n_1956),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1853),
.Y(n_2202)
);

CKINVDCx20_ASAP7_75t_R g2203 ( 
.A(n_1890),
.Y(n_2203)
);

INVx6_ASAP7_75t_L g2204 ( 
.A(n_1909),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1867),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1958),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1870),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_R g2208 ( 
.A(n_1920),
.B(n_1432),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1874),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1958),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_1946),
.Y(n_2211)
);

CKINVDCx20_ASAP7_75t_R g2212 ( 
.A(n_1909),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1856),
.Y(n_2213)
);

CKINVDCx11_ASAP7_75t_R g2214 ( 
.A(n_1906),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_2007),
.B(n_1646),
.Y(n_2215)
);

XOR2xp5_ASAP7_75t_L g2216 ( 
.A(n_1882),
.B(n_1488),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_1914),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1987),
.B(n_1179),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_1856),
.Y(n_2219)
);

BUFx10_ASAP7_75t_L g2220 ( 
.A(n_1915),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1914),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_1967),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1876),
.Y(n_2223)
);

BUFx2_ASAP7_75t_L g2224 ( 
.A(n_1881),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1880),
.Y(n_2225)
);

CKINVDCx5p33_ASAP7_75t_R g2226 ( 
.A(n_1962),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_1988),
.B(n_1314),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1899),
.Y(n_2228)
);

CKINVDCx20_ASAP7_75t_R g2229 ( 
.A(n_2023),
.Y(n_2229)
);

CKINVDCx16_ASAP7_75t_R g2230 ( 
.A(n_1934),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1916),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1857),
.Y(n_2232)
);

HB1xp67_ASAP7_75t_L g2233 ( 
.A(n_1859),
.Y(n_2233)
);

CKINVDCx16_ASAP7_75t_R g2234 ( 
.A(n_2060),
.Y(n_2234)
);

CKINVDCx20_ASAP7_75t_R g2235 ( 
.A(n_1859),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_1937),
.B(n_1485),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1900),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_1974),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_1974),
.Y(n_2239)
);

CKINVDCx5p33_ASAP7_75t_R g2240 ( 
.A(n_1976),
.Y(n_2240)
);

INVx3_ASAP7_75t_L g2241 ( 
.A(n_1946),
.Y(n_2241)
);

CKINVDCx20_ASAP7_75t_R g2242 ( 
.A(n_1976),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_2006),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1903),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_1857),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1991),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2016),
.Y(n_2247)
);

HB1xp67_ASAP7_75t_L g2248 ( 
.A(n_2006),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_2018),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2031),
.B(n_1179),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2018),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2049),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2051),
.B(n_1179),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1918),
.Y(n_2254)
);

CKINVDCx20_ASAP7_75t_R g2255 ( 
.A(n_2029),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_1970),
.Y(n_2256)
);

INVx3_ASAP7_75t_L g2257 ( 
.A(n_1955),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1869),
.B(n_1485),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_2029),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1970),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_2053),
.Y(n_2261)
);

HB1xp67_ASAP7_75t_L g2262 ( 
.A(n_2053),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_1955),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1918),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1984),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1984),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1989),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1929),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_1989),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1992),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_2028),
.B(n_1646),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1929),
.Y(n_2272)
);

INVxp67_ASAP7_75t_SL g2273 ( 
.A(n_1992),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_1931),
.Y(n_2274)
);

HB1xp67_ASAP7_75t_L g2275 ( 
.A(n_1840),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1985),
.B(n_2005),
.Y(n_2276)
);

CKINVDCx20_ASAP7_75t_R g2277 ( 
.A(n_1965),
.Y(n_2277)
);

CKINVDCx20_ASAP7_75t_R g2278 ( 
.A(n_1895),
.Y(n_2278)
);

INVx3_ASAP7_75t_L g2279 ( 
.A(n_1931),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1935),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_1925),
.Y(n_2281)
);

AND2x4_ASAP7_75t_L g2282 ( 
.A(n_2032),
.B(n_1230),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_1868),
.B(n_1102),
.Y(n_2283)
);

INVx3_ASAP7_75t_L g2284 ( 
.A(n_1935),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1942),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2036),
.B(n_1224),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1995),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1942),
.Y(n_2288)
);

OAI21x1_ASAP7_75t_L g2289 ( 
.A1(n_1948),
.A2(n_1260),
.B(n_1208),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1995),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_1936),
.B(n_1485),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_R g2292 ( 
.A(n_1925),
.B(n_1492),
.Y(n_2292)
);

INVx4_ASAP7_75t_L g2293 ( 
.A(n_1925),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2046),
.B(n_1549),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1963),
.Y(n_2295)
);

INVxp67_ASAP7_75t_L g2296 ( 
.A(n_2003),
.Y(n_2296)
);

BUFx2_ASAP7_75t_L g2297 ( 
.A(n_1940),
.Y(n_2297)
);

HB1xp67_ASAP7_75t_L g2298 ( 
.A(n_1928),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1998),
.Y(n_2299)
);

CKINVDCx20_ASAP7_75t_R g2300 ( 
.A(n_2033),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_1921),
.B(n_1235),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1963),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1998),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2002),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2002),
.Y(n_2305)
);

INVx5_ASAP7_75t_L g2306 ( 
.A(n_2012),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2012),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_L g2308 ( 
.A(n_2058),
.B(n_1103),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2034),
.Y(n_2309)
);

INVx2_ASAP7_75t_SL g2310 ( 
.A(n_1933),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_1908),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2034),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2035),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_R g2314 ( 
.A(n_1908),
.B(n_1512),
.Y(n_2314)
);

AND2x4_ASAP7_75t_L g2315 ( 
.A(n_1910),
.B(n_1960),
.Y(n_2315)
);

BUFx2_ASAP7_75t_L g2316 ( 
.A(n_1908),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2035),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2040),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_R g2319 ( 
.A(n_2037),
.B(n_1531),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2040),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2041),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_1924),
.B(n_1549),
.Y(n_2322)
);

CKINVDCx16_ASAP7_75t_R g2323 ( 
.A(n_2037),
.Y(n_2323)
);

INVxp67_ASAP7_75t_L g2324 ( 
.A(n_2041),
.Y(n_2324)
);

CKINVDCx5p33_ASAP7_75t_R g2325 ( 
.A(n_2037),
.Y(n_2325)
);

INVx3_ASAP7_75t_L g2326 ( 
.A(n_2056),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_1910),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2056),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_1949),
.B(n_1224),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_1941),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1947),
.Y(n_2331)
);

CKINVDCx20_ASAP7_75t_R g2332 ( 
.A(n_1957),
.Y(n_2332)
);

CKINVDCx5p33_ASAP7_75t_R g2333 ( 
.A(n_1951),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1959),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1964),
.Y(n_2335)
);

BUFx6f_ASAP7_75t_L g2336 ( 
.A(n_1966),
.Y(n_2336)
);

BUFx2_ASAP7_75t_L g2337 ( 
.A(n_1846),
.Y(n_2337)
);

BUFx6f_ASAP7_75t_L g2338 ( 
.A(n_1846),
.Y(n_2338)
);

BUFx2_ASAP7_75t_L g2339 ( 
.A(n_2050),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_2050),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_1854),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_1841),
.B(n_1549),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_1848),
.B(n_1224),
.Y(n_2343)
);

HB1xp67_ASAP7_75t_L g2344 ( 
.A(n_1975),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_1977),
.Y(n_2345)
);

BUFx10_ASAP7_75t_L g2346 ( 
.A(n_1979),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_1986),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1993),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_1999),
.B(n_1224),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2013),
.Y(n_2350)
);

BUFx6f_ASAP7_75t_L g2351 ( 
.A(n_2059),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2024),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_R g2353 ( 
.A(n_2030),
.B(n_1542),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_2043),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2057),
.B(n_1224),
.Y(n_2355)
);

BUFx2_ASAP7_75t_L g2356 ( 
.A(n_2045),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_2048),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1952),
.Y(n_2358)
);

CKINVDCx5p33_ASAP7_75t_R g2359 ( 
.A(n_1837),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_1981),
.B(n_1208),
.Y(n_2360)
);

NOR2x1_ASAP7_75t_L g2361 ( 
.A(n_1981),
.B(n_1243),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1952),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1952),
.Y(n_2363)
);

CKINVDCx5p33_ASAP7_75t_R g2364 ( 
.A(n_1837),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_1938),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2066),
.B(n_2070),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2076),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2067),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2338),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2338),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2338),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2079),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2289),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2103),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2068),
.B(n_1557),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_2087),
.Y(n_2376)
);

INVx2_ASAP7_75t_SL g2377 ( 
.A(n_2097),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2134),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2336),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2336),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2329),
.Y(n_2381)
);

AND3x2_ASAP7_75t_L g2382 ( 
.A(n_2078),
.B(n_1576),
.C(n_1574),
.Y(n_2382)
);

BUFx2_ASAP7_75t_L g2383 ( 
.A(n_2089),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2336),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2096),
.Y(n_2385)
);

INVx3_ASAP7_75t_L g2386 ( 
.A(n_2346),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2129),
.B(n_1580),
.Y(n_2387)
);

BUFx6f_ASAP7_75t_SL g2388 ( 
.A(n_2181),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_L g2389 ( 
.A(n_2297),
.B(n_1612),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2096),
.Y(n_2390)
);

BUFx10_ASAP7_75t_L g2391 ( 
.A(n_2192),
.Y(n_2391)
);

NAND2xp33_ASAP7_75t_R g2392 ( 
.A(n_2208),
.B(n_2292),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2096),
.Y(n_2393)
);

BUFx3_ASAP7_75t_L g2394 ( 
.A(n_2198),
.Y(n_2394)
);

INVx5_ASAP7_75t_L g2395 ( 
.A(n_2193),
.Y(n_2395)
);

INVxp33_ASAP7_75t_L g2396 ( 
.A(n_2353),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2345),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2174),
.B(n_1620),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2075),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2337),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_2067),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_2067),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2345),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2345),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2351),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2351),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2296),
.B(n_1643),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_2193),
.Y(n_2408)
);

INVx3_ASAP7_75t_L g2409 ( 
.A(n_2193),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2062),
.B(n_2077),
.Y(n_2410)
);

OR2x6_ASAP7_75t_L g2411 ( 
.A(n_2074),
.B(n_1468),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2276),
.B(n_1104),
.Y(n_2412)
);

NAND2xp33_ASAP7_75t_L g2413 ( 
.A(n_2163),
.B(n_1224),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2090),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2339),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2090),
.Y(n_2416)
);

OAI22xp33_ASAP7_75t_SL g2417 ( 
.A1(n_2080),
.A2(n_1110),
.B1(n_1114),
.B2(n_1107),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_SL g2418 ( 
.A(n_2097),
.B(n_1118),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2061),
.Y(n_2419)
);

NAND3xp33_ASAP7_75t_L g2420 ( 
.A(n_2308),
.B(n_1123),
.C(n_1119),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2063),
.Y(n_2421)
);

AOI22xp33_ASAP7_75t_L g2422 ( 
.A1(n_2085),
.A2(n_2099),
.B1(n_2101),
.B2(n_2086),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2082),
.B(n_2083),
.Y(n_2423)
);

INVx2_ASAP7_75t_SL g2424 ( 
.A(n_2098),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2093),
.B(n_1124),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2199),
.B(n_1665),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2090),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2064),
.Y(n_2428)
);

NAND2xp33_ASAP7_75t_L g2429 ( 
.A(n_2163),
.B(n_1224),
.Y(n_2429)
);

OR2x2_ASAP7_75t_L g2430 ( 
.A(n_2359),
.B(n_1171),
.Y(n_2430)
);

HB1xp67_ASAP7_75t_L g2431 ( 
.A(n_2364),
.Y(n_2431)
);

CKINVDCx14_ASAP7_75t_R g2432 ( 
.A(n_2160),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2071),
.Y(n_2433)
);

BUFx6f_ASAP7_75t_SL g2434 ( 
.A(n_2194),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_SL g2435 ( 
.A(n_2098),
.B(n_1130),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2219),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2219),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2219),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2358),
.Y(n_2439)
);

BUFx3_ASAP7_75t_L g2440 ( 
.A(n_2203),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2245),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2362),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2236),
.B(n_2145),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2363),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2245),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2245),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2196),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2322),
.B(n_1131),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2256),
.Y(n_2449)
);

NAND3xp33_ASAP7_75t_L g2450 ( 
.A(n_2073),
.B(n_1134),
.C(n_1133),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2224),
.B(n_1135),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2256),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2256),
.Y(n_2453)
);

INVx1_ASAP7_75t_SL g2454 ( 
.A(n_2136),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2168),
.B(n_2111),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2323),
.B(n_1138),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2269),
.Y(n_2457)
);

INVx4_ASAP7_75t_L g2458 ( 
.A(n_2074),
.Y(n_2458)
);

INVx5_ASAP7_75t_L g2459 ( 
.A(n_2150),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2269),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2269),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2151),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2065),
.Y(n_2463)
);

AND2x4_ASAP7_75t_L g2464 ( 
.A(n_2141),
.B(n_1248),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2069),
.Y(n_2465)
);

BUFx3_ASAP7_75t_L g2466 ( 
.A(n_2212),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2205),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2234),
.B(n_1682),
.Y(n_2468)
);

AND3x2_ASAP7_75t_L g2469 ( 
.A(n_2275),
.B(n_1258),
.C(n_1253),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2116),
.Y(n_2470)
);

INVx2_ASAP7_75t_SL g2471 ( 
.A(n_2220),
.Y(n_2471)
);

HB1xp67_ASAP7_75t_L g2472 ( 
.A(n_2094),
.Y(n_2472)
);

INVx2_ASAP7_75t_SL g2473 ( 
.A(n_2108),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2207),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2365),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2092),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2126),
.B(n_1139),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2126),
.B(n_1140),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2102),
.B(n_1268),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2331),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2126),
.B(n_1151),
.Y(n_2481)
);

BUFx10_ASAP7_75t_L g2482 ( 
.A(n_2127),
.Y(n_2482)
);

AOI22xp5_ASAP7_75t_L g2483 ( 
.A1(n_2278),
.A2(n_1157),
.B1(n_1159),
.B2(n_1152),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2209),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2095),
.B(n_1162),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2151),
.Y(n_2486)
);

AOI22xp5_ASAP7_75t_L g2487 ( 
.A1(n_2332),
.A2(n_1165),
.B1(n_1166),
.B2(n_1163),
.Y(n_2487)
);

HB1xp67_ASAP7_75t_L g2488 ( 
.A(n_2094),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2223),
.Y(n_2489)
);

BUFx6f_ASAP7_75t_SL g2490 ( 
.A(n_2106),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2225),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2228),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2334),
.Y(n_2493)
);

BUFx2_ASAP7_75t_L g2494 ( 
.A(n_2088),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2335),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2237),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2185),
.Y(n_2497)
);

AOI21x1_ASAP7_75t_L g2498 ( 
.A1(n_2149),
.A2(n_1277),
.B(n_1276),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2244),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2340),
.B(n_1167),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2231),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2344),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2342),
.B(n_1168),
.Y(n_2503)
);

CKINVDCx6p67_ASAP7_75t_R g2504 ( 
.A(n_2214),
.Y(n_2504)
);

AOI22xp33_ASAP7_75t_L g2505 ( 
.A1(n_2110),
.A2(n_2115),
.B1(n_2119),
.B2(n_2117),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2189),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2282),
.B(n_1170),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2282),
.B(n_1172),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2121),
.B(n_1173),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2135),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2137),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2138),
.Y(n_2512)
);

INVxp67_ASAP7_75t_SL g2513 ( 
.A(n_2114),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2125),
.B(n_1174),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2163),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2132),
.B(n_1175),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2348),
.Y(n_2517)
);

INVx4_ASAP7_75t_L g2518 ( 
.A(n_2204),
.Y(n_2518)
);

INVx2_ASAP7_75t_SL g2519 ( 
.A(n_2131),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2350),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2356),
.Y(n_2521)
);

NAND3xp33_ASAP7_75t_L g2522 ( 
.A(n_2283),
.B(n_1178),
.C(n_1177),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2352),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_2306),
.Y(n_2524)
);

OR2x6_ASAP7_75t_L g2525 ( 
.A(n_2204),
.B(n_1260),
.Y(n_2525)
);

NAND2xp33_ASAP7_75t_L g2526 ( 
.A(n_2150),
.B(n_1339),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2188),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2188),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2072),
.B(n_1180),
.Y(n_2529)
);

AND2x4_ASAP7_75t_L g2530 ( 
.A(n_2315),
.B(n_1280),
.Y(n_2530)
);

CKINVDCx5p33_ASAP7_75t_R g2531 ( 
.A(n_2162),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2151),
.Y(n_2532)
);

AND2x4_ASAP7_75t_L g2533 ( 
.A(n_2315),
.B(n_1283),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2159),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2215),
.Y(n_2535)
);

INVx5_ASAP7_75t_L g2536 ( 
.A(n_2150),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2159),
.Y(n_2537)
);

INVx2_ASAP7_75t_SL g2538 ( 
.A(n_2081),
.Y(n_2538)
);

AND3x1_ASAP7_75t_L g2539 ( 
.A(n_2153),
.B(n_1289),
.C(n_1286),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2159),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2215),
.Y(n_2541)
);

AOI22xp33_ASAP7_75t_L g2542 ( 
.A1(n_2271),
.A2(n_1128),
.B1(n_1405),
.B2(n_1339),
.Y(n_2542)
);

BUFx6f_ASAP7_75t_L g2543 ( 
.A(n_2091),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_2306),
.Y(n_2544)
);

BUFx3_ASAP7_75t_L g2545 ( 
.A(n_2118),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2330),
.B(n_1183),
.Y(n_2546)
);

NOR2xp33_ASAP7_75t_R g2547 ( 
.A(n_2166),
.B(n_1186),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_L g2548 ( 
.A(n_2182),
.B(n_1187),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2156),
.Y(n_2549)
);

BUFx2_ASAP7_75t_L g2550 ( 
.A(n_2120),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_2258),
.B(n_2133),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2091),
.Y(n_2552)
);

INVx8_ASAP7_75t_L g2553 ( 
.A(n_2170),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2091),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2107),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2333),
.B(n_1188),
.Y(n_2556)
);

INVx6_ASAP7_75t_L g2557 ( 
.A(n_2179),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_2173),
.Y(n_2558)
);

AND3x2_ASAP7_75t_L g2559 ( 
.A(n_2130),
.B(n_1309),
.C(n_1291),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2072),
.B(n_1189),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2271),
.Y(n_2561)
);

INVx2_ASAP7_75t_SL g2562 ( 
.A(n_2314),
.Y(n_2562)
);

OR2x6_ASAP7_75t_L g2563 ( 
.A(n_2310),
.B(n_1265),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2112),
.B(n_1191),
.Y(n_2564)
);

INVx3_ASAP7_75t_L g2565 ( 
.A(n_2306),
.Y(n_2565)
);

AND3x2_ASAP7_75t_L g2566 ( 
.A(n_2142),
.B(n_1332),
.C(n_1319),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2146),
.Y(n_2567)
);

BUFx4f_ASAP7_75t_L g2568 ( 
.A(n_2301),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2301),
.B(n_1194),
.Y(n_2569)
);

BUFx3_ASAP7_75t_L g2570 ( 
.A(n_2201),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2218),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2341),
.B(n_1200),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2250),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2253),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2246),
.Y(n_2575)
);

INVxp33_ASAP7_75t_L g2576 ( 
.A(n_2298),
.Y(n_2576)
);

INVx3_ASAP7_75t_L g2577 ( 
.A(n_2274),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2347),
.B(n_2354),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2152),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2155),
.Y(n_2580)
);

INVx2_ASAP7_75t_SL g2581 ( 
.A(n_2319),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2293),
.B(n_1201),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2247),
.Y(n_2583)
);

INVx2_ASAP7_75t_SL g2584 ( 
.A(n_2357),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2161),
.B(n_1205),
.Y(n_2585)
);

NAND2xp33_ASAP7_75t_L g2586 ( 
.A(n_2311),
.B(n_2325),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2252),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2179),
.B(n_1206),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2172),
.B(n_1210),
.Y(n_2589)
);

INVx4_ASAP7_75t_L g2590 ( 
.A(n_2281),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2140),
.Y(n_2591)
);

CKINVDCx20_ASAP7_75t_R g2592 ( 
.A(n_2177),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2286),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2158),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2291),
.B(n_1211),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_2084),
.B(n_1213),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2164),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2165),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2124),
.B(n_1215),
.Y(n_2599)
);

INVxp67_ASAP7_75t_L g2600 ( 
.A(n_2128),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2144),
.B(n_1217),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2169),
.Y(n_2602)
);

BUFx2_ASAP7_75t_L g2603 ( 
.A(n_2105),
.Y(n_2603)
);

CKINVDCx5p33_ASAP7_75t_R g2604 ( 
.A(n_2184),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2316),
.B(n_2147),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2183),
.Y(n_2606)
);

INVx2_ASAP7_75t_SL g2607 ( 
.A(n_2113),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2100),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2360),
.Y(n_2609)
);

INVx1_ASAP7_75t_SL g2610 ( 
.A(n_2235),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2277),
.B(n_1218),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2195),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2197),
.Y(n_2613)
);

INVxp33_ASAP7_75t_L g2614 ( 
.A(n_2122),
.Y(n_2614)
);

INVx3_ASAP7_75t_L g2615 ( 
.A(n_2279),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2300),
.B(n_1219),
.Y(n_2616)
);

INVx5_ASAP7_75t_L g2617 ( 
.A(n_2211),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2361),
.B(n_1220),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_SL g2619 ( 
.A(n_2154),
.B(n_1226),
.Y(n_2619)
);

CKINVDCx20_ASAP7_75t_R g2620 ( 
.A(n_2186),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2324),
.B(n_1227),
.Y(n_2621)
);

NAND2xp33_ASAP7_75t_L g2622 ( 
.A(n_2343),
.B(n_1339),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2202),
.Y(n_2623)
);

INVx2_ASAP7_75t_SL g2624 ( 
.A(n_2327),
.Y(n_2624)
);

AND2x4_ASAP7_75t_L g2625 ( 
.A(n_2227),
.B(n_1335),
.Y(n_2625)
);

INVx5_ASAP7_75t_L g2626 ( 
.A(n_2241),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2213),
.Y(n_2627)
);

CKINVDCx20_ASAP7_75t_R g2628 ( 
.A(n_2187),
.Y(n_2628)
);

INVx3_ASAP7_75t_L g2629 ( 
.A(n_2284),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2230),
.B(n_1231),
.Y(n_2630)
);

NAND2xp33_ASAP7_75t_SL g2631 ( 
.A(n_2229),
.B(n_1233),
.Y(n_2631)
);

NAND2xp33_ASAP7_75t_L g2632 ( 
.A(n_2349),
.B(n_2355),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2294),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2326),
.B(n_1234),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2232),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2123),
.B(n_1238),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2148),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2260),
.Y(n_2638)
);

AOI22xp33_ASAP7_75t_L g2639 ( 
.A1(n_2254),
.A2(n_1128),
.B1(n_1405),
.B2(n_1339),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_2167),
.B(n_1239),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2233),
.B(n_2248),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2171),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2175),
.Y(n_2643)
);

NOR2xp33_ASAP7_75t_L g2644 ( 
.A(n_2251),
.B(n_1240),
.Y(n_2644)
);

INVx8_ASAP7_75t_L g2645 ( 
.A(n_2190),
.Y(n_2645)
);

CKINVDCx6p67_ASAP7_75t_R g2646 ( 
.A(n_2242),
.Y(n_2646)
);

OR2x2_ASAP7_75t_L g2647 ( 
.A(n_2200),
.B(n_1269),
.Y(n_2647)
);

AND2x6_ASAP7_75t_L g2648 ( 
.A(n_2264),
.B(n_2268),
.Y(n_2648)
);

AOI22xp33_ASAP7_75t_L g2649 ( 
.A1(n_2272),
.A2(n_1405),
.B1(n_1497),
.B2(n_1339),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2176),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2265),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2266),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2139),
.B(n_1241),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2273),
.B(n_1242),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2178),
.Y(n_2655)
);

BUFx6f_ASAP7_75t_L g2656 ( 
.A(n_2267),
.Y(n_2656)
);

INVxp33_ASAP7_75t_L g2657 ( 
.A(n_2262),
.Y(n_2657)
);

NAND3xp33_ASAP7_75t_L g2658 ( 
.A(n_2217),
.B(n_1245),
.C(n_1244),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2180),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2280),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2270),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2287),
.Y(n_2662)
);

CKINVDCx5p33_ASAP7_75t_R g2663 ( 
.A(n_2143),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_SL g2664 ( 
.A(n_2290),
.B(n_1246),
.Y(n_2664)
);

BUFx6f_ASAP7_75t_SL g2665 ( 
.A(n_2191),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2285),
.Y(n_2666)
);

INVxp67_ASAP7_75t_SL g2667 ( 
.A(n_2255),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2288),
.Y(n_2668)
);

BUFx3_ASAP7_75t_L g2669 ( 
.A(n_2104),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2299),
.Y(n_2670)
);

CKINVDCx6p67_ASAP7_75t_R g2671 ( 
.A(n_2109),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2295),
.B(n_1249),
.Y(n_2672)
);

AND2x4_ASAP7_75t_L g2673 ( 
.A(n_2257),
.B(n_1338),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2304),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2309),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2318),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2157),
.B(n_2221),
.Y(n_2677)
);

INVx4_ASAP7_75t_L g2678 ( 
.A(n_2238),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2328),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2302),
.Y(n_2680)
);

INVx3_ASAP7_75t_L g2681 ( 
.A(n_2303),
.Y(n_2681)
);

INVx3_ASAP7_75t_L g2682 ( 
.A(n_2305),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2307),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2312),
.B(n_1252),
.Y(n_2684)
);

CKINVDCx20_ASAP7_75t_R g2685 ( 
.A(n_2222),
.Y(n_2685)
);

INVx4_ASAP7_75t_L g2686 ( 
.A(n_2239),
.Y(n_2686)
);

AOI22xp33_ASAP7_75t_L g2687 ( 
.A1(n_2313),
.A2(n_1405),
.B1(n_1497),
.B2(n_1339),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2317),
.Y(n_2688)
);

OR2x2_ASAP7_75t_L g2689 ( 
.A(n_2216),
.B(n_1295),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2320),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2321),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2263),
.B(n_1254),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2240),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2243),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_2249),
.B(n_1255),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_SL g2696 ( 
.A(n_2259),
.B(n_1256),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2261),
.B(n_1257),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2226),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_L g2699 ( 
.A(n_2206),
.B(n_1262),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_SL g2700 ( 
.A(n_2210),
.B(n_1266),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2338),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2066),
.B(n_1270),
.Y(n_2702)
);

AOI22xp33_ASAP7_75t_SL g2703 ( 
.A1(n_2292),
.A2(n_1275),
.B1(n_1281),
.B2(n_1271),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2338),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2338),
.Y(n_2705)
);

BUFx10_ASAP7_75t_L g2706 ( 
.A(n_2192),
.Y(n_2706)
);

NAND2xp33_ASAP7_75t_R g2707 ( 
.A(n_2208),
.B(n_1284),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2066),
.B(n_1285),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2338),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2338),
.Y(n_2710)
);

INVx3_ASAP7_75t_L g2711 ( 
.A(n_2336),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2338),
.Y(n_2712)
);

OAI22xp33_ASAP7_75t_SL g2713 ( 
.A1(n_2075),
.A2(n_1298),
.B1(n_1300),
.B2(n_1299),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2338),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2076),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2076),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_SL g2717 ( 
.A(n_2066),
.B(n_1301),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2076),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2338),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2276),
.B(n_1303),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2338),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2338),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2068),
.B(n_1304),
.Y(n_2723)
);

AOI21x1_ASAP7_75t_L g2724 ( 
.A1(n_2065),
.A2(n_1341),
.B(n_1340),
.Y(n_2724)
);

INVxp67_ASAP7_75t_SL g2725 ( 
.A(n_2078),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_SL g2726 ( 
.A(n_2066),
.B(n_1305),
.Y(n_2726)
);

INVx4_ASAP7_75t_L g2727 ( 
.A(n_2097),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2338),
.Y(n_2728)
);

NAND3xp33_ASAP7_75t_L g2729 ( 
.A(n_2308),
.B(n_1307),
.C(n_1306),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2338),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2076),
.Y(n_2731)
);

BUFx3_ASAP7_75t_L g2732 ( 
.A(n_2198),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2076),
.Y(n_2733)
);

INVx3_ASAP7_75t_L g2734 ( 
.A(n_2336),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_2087),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2076),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2076),
.Y(n_2737)
);

INVx2_ASAP7_75t_SL g2738 ( 
.A(n_2097),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2338),
.Y(n_2739)
);

INVx3_ASAP7_75t_L g2740 ( 
.A(n_2336),
.Y(n_2740)
);

INVx3_ASAP7_75t_L g2741 ( 
.A(n_2336),
.Y(n_2741)
);

NAND3xp33_ASAP7_75t_L g2742 ( 
.A(n_2308),
.B(n_1311),
.C(n_1310),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2076),
.Y(n_2743)
);

BUFx2_ASAP7_75t_L g2744 ( 
.A(n_2087),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2076),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2338),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_2087),
.Y(n_2747)
);

BUFx6f_ASAP7_75t_L g2748 ( 
.A(n_2368),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2447),
.Y(n_2749)
);

BUFx6f_ASAP7_75t_L g2750 ( 
.A(n_2368),
.Y(n_2750)
);

INVx1_ASAP7_75t_SL g2751 ( 
.A(n_2454),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2412),
.B(n_1315),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2720),
.B(n_1316),
.Y(n_2753)
);

INVxp33_ASAP7_75t_L g2754 ( 
.A(n_2468),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2467),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2407),
.B(n_2389),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_SL g2757 ( 
.A(n_2568),
.B(n_1317),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_SL g2758 ( 
.A(n_2459),
.B(n_1320),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2723),
.B(n_1322),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2422),
.B(n_2505),
.Y(n_2760)
);

INVxp67_ASAP7_75t_L g2761 ( 
.A(n_2725),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2367),
.B(n_1323),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2367),
.B(n_1324),
.Y(n_2763)
);

NOR2xp67_ASAP7_75t_L g2764 ( 
.A(n_2376),
.B(n_83),
.Y(n_2764)
);

INVx3_ASAP7_75t_L g2765 ( 
.A(n_2395),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2374),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_L g2767 ( 
.A(n_2426),
.B(n_1326),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2474),
.Y(n_2768)
);

NOR2xp67_ASAP7_75t_L g2769 ( 
.A(n_2735),
.B(n_83),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2502),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_SL g2771 ( 
.A(n_2568),
.B(n_1327),
.Y(n_2771)
);

HB1xp67_ASAP7_75t_L g2772 ( 
.A(n_2383),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_SL g2773 ( 
.A(n_2386),
.B(n_1330),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2372),
.B(n_1331),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2372),
.B(n_1333),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2374),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2378),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2378),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2443),
.B(n_1334),
.Y(n_2779)
);

NAND2xp33_ASAP7_75t_L g2780 ( 
.A(n_2543),
.B(n_1337),
.Y(n_2780)
);

INVxp67_ASAP7_75t_L g2781 ( 
.A(n_2744),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_2386),
.B(n_1342),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2715),
.B(n_1343),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2484),
.Y(n_2784)
);

AO221x1_ASAP7_75t_L g2785 ( 
.A1(n_2494),
.A2(n_1236),
.B1(n_1237),
.B2(n_1199),
.C(n_1126),
.Y(n_2785)
);

BUFx3_ASAP7_75t_L g2786 ( 
.A(n_2394),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2484),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_SL g2788 ( 
.A(n_2584),
.B(n_1344),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2489),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2489),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2491),
.Y(n_2791)
);

BUFx3_ASAP7_75t_L g2792 ( 
.A(n_2732),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_2703),
.B(n_1345),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2491),
.B(n_1346),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2492),
.Y(n_2795)
);

NAND2xp33_ASAP7_75t_L g2796 ( 
.A(n_2543),
.B(n_1347),
.Y(n_2796)
);

A2O1A1Ixp33_ASAP7_75t_L g2797 ( 
.A1(n_2506),
.A2(n_1267),
.B(n_1290),
.C(n_1265),
.Y(n_2797)
);

NOR3xp33_ASAP7_75t_L g2798 ( 
.A(n_2631),
.B(n_1328),
.C(n_1297),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_SL g2799 ( 
.A(n_2747),
.B(n_1352),
.Y(n_2799)
);

OA21x2_ASAP7_75t_L g2800 ( 
.A1(n_2373),
.A2(n_1290),
.B(n_1267),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2492),
.B(n_2496),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2496),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_SL g2803 ( 
.A(n_2578),
.B(n_1356),
.Y(n_2803)
);

CKINVDCx20_ASAP7_75t_R g2804 ( 
.A(n_2504),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2455),
.B(n_1357),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_2423),
.B(n_1362),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_SL g2807 ( 
.A(n_2399),
.B(n_1363),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_L g2808 ( 
.A(n_2387),
.B(n_2410),
.Y(n_2808)
);

AOI22xp33_ASAP7_75t_L g2809 ( 
.A1(n_2611),
.A2(n_1366),
.B1(n_1367),
.B2(n_1364),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2499),
.B(n_1368),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_SL g2811 ( 
.A(n_2430),
.B(n_1374),
.Y(n_2811)
);

NOR2xp33_ASAP7_75t_L g2812 ( 
.A(n_2398),
.B(n_1377),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2499),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2375),
.B(n_2529),
.Y(n_2814)
);

INVxp33_ASAP7_75t_L g2815 ( 
.A(n_2547),
.Y(n_2815)
);

AND2x6_ASAP7_75t_SL g2816 ( 
.A(n_2411),
.B(n_1351),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_L g2817 ( 
.A(n_2616),
.B(n_1379),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_L g2818 ( 
.A(n_2366),
.B(n_1380),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2419),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_SL g2820 ( 
.A(n_2459),
.B(n_1382),
.Y(n_2820)
);

XOR2xp5_ASAP7_75t_L g2821 ( 
.A(n_2620),
.B(n_1384),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_2458),
.B(n_1354),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2421),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2715),
.Y(n_2824)
);

INVx3_ASAP7_75t_L g2825 ( 
.A(n_2395),
.Y(n_2825)
);

AOI221xp5_ASAP7_75t_L g2826 ( 
.A1(n_2417),
.A2(n_1391),
.B1(n_1392),
.B2(n_1389),
.C(n_1387),
.Y(n_2826)
);

BUFx5_ASAP7_75t_L g2827 ( 
.A(n_2390),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2716),
.Y(n_2828)
);

NOR2xp33_ASAP7_75t_L g2829 ( 
.A(n_2431),
.B(n_1393),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2428),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2433),
.B(n_1396),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2458),
.B(n_2576),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2439),
.B(n_1399),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2716),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_2470),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2442),
.Y(n_2836)
);

INVxp67_ASAP7_75t_L g2837 ( 
.A(n_2563),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_SL g2838 ( 
.A(n_2459),
.B(n_1400),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2444),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2718),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_SL g2841 ( 
.A(n_2536),
.B(n_1401),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2564),
.B(n_2425),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2400),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2479),
.B(n_1402),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_SL g2845 ( 
.A(n_2536),
.B(n_1404),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_SL g2846 ( 
.A(n_2536),
.B(n_1406),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2479),
.B(n_1407),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2415),
.Y(n_2848)
);

BUFx6f_ASAP7_75t_SL g2849 ( 
.A(n_2391),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2718),
.B(n_1411),
.Y(n_2850)
);

INVxp67_ASAP7_75t_L g2851 ( 
.A(n_2563),
.Y(n_2851)
);

INVx2_ASAP7_75t_SL g2852 ( 
.A(n_2391),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2510),
.Y(n_2853)
);

AO221x1_ASAP7_75t_L g2854 ( 
.A1(n_2600),
.A2(n_1236),
.B1(n_1237),
.B2(n_1199),
.C(n_1126),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_L g2855 ( 
.A(n_2396),
.B(n_1412),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2551),
.B(n_2557),
.Y(n_2856)
);

NAND2xp33_ASAP7_75t_L g2857 ( 
.A(n_2543),
.B(n_2648),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_SL g2858 ( 
.A(n_2395),
.B(n_1413),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2731),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2731),
.B(n_2733),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_L g2861 ( 
.A(n_2557),
.B(n_1415),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_SL g2862 ( 
.A(n_2599),
.B(n_1416),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2451),
.B(n_1418),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2733),
.Y(n_2864)
);

AOI22xp5_ASAP7_75t_L g2865 ( 
.A1(n_2487),
.A2(n_1422),
.B1(n_1423),
.B2(n_1420),
.Y(n_2865)
);

OR2x2_ASAP7_75t_L g2866 ( 
.A(n_2647),
.B(n_1514),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2736),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2736),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2546),
.B(n_1425),
.Y(n_2869)
);

NOR3xp33_ASAP7_75t_L g2870 ( 
.A(n_2713),
.B(n_1360),
.C(n_1349),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2511),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2737),
.B(n_1426),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2560),
.B(n_1428),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2737),
.B(n_2743),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2480),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2493),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_SL g2877 ( 
.A(n_2556),
.B(n_1431),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2572),
.B(n_1433),
.Y(n_2878)
);

INVxp33_ASAP7_75t_SL g2879 ( 
.A(n_2531),
.Y(n_2879)
);

INVxp67_ASAP7_75t_L g2880 ( 
.A(n_2525),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2743),
.B(n_1436),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_SL g2882 ( 
.A(n_2483),
.B(n_1438),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2745),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2495),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2745),
.B(n_1441),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_SL g2886 ( 
.A(n_2471),
.B(n_1445),
.Y(n_2886)
);

BUFx5_ASAP7_75t_L g2887 ( 
.A(n_2390),
.Y(n_2887)
);

NAND2xp33_ASAP7_75t_L g2888 ( 
.A(n_2648),
.B(n_1448),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2497),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2501),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2507),
.B(n_1452),
.Y(n_2891)
);

NAND2xp33_ASAP7_75t_L g2892 ( 
.A(n_2648),
.B(n_1453),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2500),
.B(n_1454),
.Y(n_2893)
);

BUFx6f_ASAP7_75t_L g2894 ( 
.A(n_2368),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2724),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2512),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2485),
.B(n_1455),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2521),
.Y(n_2898)
);

INVxp33_ASAP7_75t_L g2899 ( 
.A(n_2603),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2702),
.B(n_1456),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_SL g2901 ( 
.A(n_2508),
.B(n_1463),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2517),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2463),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_2448),
.B(n_1464),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2464),
.B(n_1470),
.Y(n_2905)
);

BUFx6f_ASAP7_75t_SL g2906 ( 
.A(n_2706),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2708),
.B(n_1473),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_L g2908 ( 
.A(n_2401),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2465),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2717),
.B(n_1478),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2726),
.B(n_1481),
.Y(n_2911)
);

BUFx2_ASAP7_75t_L g2912 ( 
.A(n_2525),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2520),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_SL g2914 ( 
.A(n_2697),
.B(n_1486),
.Y(n_2914)
);

OR2x6_ASAP7_75t_L g2915 ( 
.A(n_2645),
.B(n_2411),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2523),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2569),
.B(n_1487),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2464),
.B(n_1493),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2509),
.B(n_1495),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_2477),
.B(n_2478),
.Y(n_2920)
);

NOR2x1p5_ASAP7_75t_L g2921 ( 
.A(n_2646),
.B(n_1496),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2575),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2514),
.B(n_1498),
.Y(n_2923)
);

BUFx5_ASAP7_75t_L g2924 ( 
.A(n_2393),
.Y(n_2924)
);

BUFx6f_ASAP7_75t_L g2925 ( 
.A(n_2401),
.Y(n_2925)
);

NOR2xp67_ASAP7_75t_L g2926 ( 
.A(n_2558),
.B(n_2604),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2506),
.B(n_1499),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2593),
.B(n_1500),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2583),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2587),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2630),
.B(n_1501),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2516),
.B(n_1502),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2475),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2481),
.B(n_1503),
.Y(n_2934)
);

INVxp67_ASAP7_75t_L g2935 ( 
.A(n_2707),
.Y(n_2935)
);

NOR3xp33_ASAP7_75t_L g2936 ( 
.A(n_2450),
.B(n_1403),
.C(n_1373),
.Y(n_2936)
);

NOR2xp33_ASAP7_75t_L g2937 ( 
.A(n_2657),
.B(n_1505),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2593),
.B(n_1506),
.Y(n_2938)
);

AND2x2_ASAP7_75t_L g2939 ( 
.A(n_2530),
.B(n_1507),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2527),
.Y(n_2940)
);

NAND2xp33_ASAP7_75t_SL g2941 ( 
.A(n_2392),
.B(n_1685),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2528),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2476),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2591),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2614),
.B(n_1510),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2530),
.B(n_1515),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2535),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_2644),
.B(n_1518),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2498),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_SL g2950 ( 
.A(n_2594),
.B(n_1521),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2533),
.B(n_1523),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2541),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2561),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2637),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2642),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_SL g2956 ( 
.A(n_2594),
.B(n_1524),
.Y(n_2956)
);

INVxp33_ASAP7_75t_L g2957 ( 
.A(n_2550),
.Y(n_2957)
);

NOR3xp33_ASAP7_75t_L g2958 ( 
.A(n_2522),
.B(n_1522),
.C(n_1437),
.Y(n_2958)
);

NOR3xp33_ASAP7_75t_L g2959 ( 
.A(n_2420),
.B(n_1600),
.C(n_1595),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_2503),
.B(n_1528),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2533),
.B(n_1529),
.Y(n_2961)
);

BUFx5_ASAP7_75t_L g2962 ( 
.A(n_2393),
.Y(n_2962)
);

NOR2xp33_ASAP7_75t_L g2963 ( 
.A(n_2595),
.B(n_1530),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2472),
.B(n_1532),
.Y(n_2964)
);

CKINVDCx20_ASAP7_75t_R g2965 ( 
.A(n_2628),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2625),
.B(n_1533),
.Y(n_2966)
);

INVx8_ASAP7_75t_L g2967 ( 
.A(n_2490),
.Y(n_2967)
);

INVxp67_ASAP7_75t_L g2968 ( 
.A(n_2545),
.Y(n_2968)
);

INVxp33_ASAP7_75t_L g2969 ( 
.A(n_2641),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2673),
.Y(n_2970)
);

INVx2_ASAP7_75t_SL g2971 ( 
.A(n_2706),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2625),
.B(n_1534),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2633),
.B(n_1537),
.Y(n_2973)
);

INVxp67_ASAP7_75t_L g2974 ( 
.A(n_2488),
.Y(n_2974)
);

A2O1A1Ixp33_ASAP7_75t_L g2975 ( 
.A1(n_2381),
.A2(n_1318),
.B(n_1321),
.C(n_1292),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2601),
.B(n_1539),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2673),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2469),
.B(n_1543),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2609),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2548),
.B(n_1544),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2588),
.B(n_1545),
.Y(n_2981)
);

NOR3xp33_ASAP7_75t_L g2982 ( 
.A(n_2729),
.B(n_1696),
.C(n_1695),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2381),
.B(n_1547),
.Y(n_2983)
);

INVxp67_ASAP7_75t_L g2984 ( 
.A(n_2490),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2654),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2643),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_2665),
.Y(n_2987)
);

NOR2xp33_ASAP7_75t_L g2988 ( 
.A(n_2562),
.B(n_1548),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2672),
.Y(n_2989)
);

BUFx5_ASAP7_75t_L g2990 ( 
.A(n_2648),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2571),
.B(n_1550),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_SL g2992 ( 
.A(n_2607),
.B(n_1552),
.Y(n_2992)
);

BUFx6f_ASAP7_75t_L g2993 ( 
.A(n_2401),
.Y(n_2993)
);

NAND3xp33_ASAP7_75t_L g2994 ( 
.A(n_2526),
.B(n_1199),
.C(n_1126),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_SL g2995 ( 
.A(n_2473),
.B(n_1553),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2650),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_SL g2997 ( 
.A(n_2519),
.B(n_1554),
.Y(n_2997)
);

AND2x2_ASAP7_75t_L g2998 ( 
.A(n_2636),
.B(n_1555),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2684),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2655),
.Y(n_3000)
);

AOI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2677),
.A2(n_1559),
.B1(n_1561),
.B2(n_1556),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2653),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2659),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2692),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2402),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2660),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_SL g3007 ( 
.A(n_2581),
.B(n_1562),
.Y(n_3007)
);

BUFx5_ASAP7_75t_L g3008 ( 
.A(n_2597),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2573),
.B(n_1564),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2574),
.B(n_1565),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2666),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2668),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2680),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_SL g3014 ( 
.A(n_2597),
.B(n_2658),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2585),
.B(n_1568),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2690),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2513),
.Y(n_3017)
);

NAND2xp33_ASAP7_75t_L g3018 ( 
.A(n_2402),
.B(n_1592),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2618),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2589),
.B(n_2742),
.Y(n_3020)
);

INVx4_ASAP7_75t_L g3021 ( 
.A(n_2388),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2608),
.B(n_1570),
.Y(n_3022)
);

INVx2_ASAP7_75t_SL g3023 ( 
.A(n_2553),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2596),
.B(n_1573),
.Y(n_3024)
);

NOR2xp33_ASAP7_75t_L g3025 ( 
.A(n_2624),
.B(n_1575),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2664),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2634),
.Y(n_3027)
);

NAND3xp33_ASAP7_75t_L g3028 ( 
.A(n_2542),
.B(n_2622),
.C(n_2429),
.Y(n_3028)
);

NAND3xp33_ASAP7_75t_L g3029 ( 
.A(n_2413),
.B(n_1199),
.C(n_1126),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2683),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_L g3031 ( 
.A(n_2456),
.B(n_1577),
.Y(n_3031)
);

NOR2xp33_ASAP7_75t_L g3032 ( 
.A(n_2570),
.B(n_2669),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2418),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2435),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2549),
.B(n_2377),
.Y(n_3035)
);

AND2x6_ASAP7_75t_SL g3036 ( 
.A(n_2432),
.B(n_2592),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2549),
.B(n_1578),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_SL g3038 ( 
.A(n_2727),
.B(n_1582),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2424),
.B(n_1587),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_SL g3040 ( 
.A(n_2727),
.B(n_1588),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2738),
.B(n_1591),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2619),
.B(n_1594),
.Y(n_3042)
);

NAND3xp33_ASAP7_75t_L g3043 ( 
.A(n_2649),
.B(n_1237),
.C(n_1236),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2640),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2688),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2621),
.B(n_1597),
.Y(n_3046)
);

BUFx6f_ASAP7_75t_L g3047 ( 
.A(n_2402),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2691),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2369),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2370),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2582),
.B(n_1598),
.Y(n_3051)
);

OR2x2_ASAP7_75t_L g3052 ( 
.A(n_2689),
.B(n_1604),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2605),
.B(n_1605),
.Y(n_3053)
);

OAI21xp33_ASAP7_75t_L g3054 ( 
.A1(n_2699),
.A2(n_1607),
.B(n_1606),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2678),
.B(n_1608),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2538),
.B(n_1609),
.Y(n_3056)
);

NOR3xp33_ASAP7_75t_L g3057 ( 
.A(n_2700),
.B(n_1358),
.C(n_1355),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2693),
.B(n_1610),
.Y(n_3058)
);

BUFx5_ASAP7_75t_L g3059 ( 
.A(n_2462),
.Y(n_3059)
);

NAND2xp33_ASAP7_75t_L g3060 ( 
.A(n_2462),
.B(n_1613),
.Y(n_3060)
);

INVx3_ASAP7_75t_L g3061 ( 
.A(n_2408),
.Y(n_3061)
);

AOI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2632),
.A2(n_1369),
.B(n_1361),
.Y(n_3062)
);

AO221x1_ASAP7_75t_L g3063 ( 
.A1(n_2382),
.A2(n_1282),
.B1(n_1287),
.B2(n_1237),
.C(n_1236),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2695),
.B(n_2696),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2524),
.Y(n_3065)
);

INVx4_ASAP7_75t_L g3066 ( 
.A(n_2388),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2524),
.Y(n_3067)
);

BUFx5_ASAP7_75t_L g3068 ( 
.A(n_2462),
.Y(n_3068)
);

HB1xp67_ASAP7_75t_L g3069 ( 
.A(n_2434),
.Y(n_3069)
);

NOR2xp67_ASAP7_75t_L g3070 ( 
.A(n_2678),
.B(n_89),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2544),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_2539),
.B(n_1611),
.Y(n_3072)
);

BUFx6f_ASAP7_75t_L g3073 ( 
.A(n_2486),
.Y(n_3073)
);

NAND2xp33_ASAP7_75t_L g3074 ( 
.A(n_2486),
.B(n_1631),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2544),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_L g3076 ( 
.A(n_2694),
.B(n_1614),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2371),
.Y(n_3077)
);

NOR3xp33_ASAP7_75t_L g3078 ( 
.A(n_2667),
.B(n_1372),
.C(n_1371),
.Y(n_3078)
);

AOI221xp5_ASAP7_75t_L g3079 ( 
.A1(n_2610),
.A2(n_2665),
.B1(n_2434),
.B2(n_2663),
.C(n_2466),
.Y(n_3079)
);

OR2x2_ASAP7_75t_SL g3080 ( 
.A(n_2698),
.B(n_1378),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_SL g3081 ( 
.A(n_2686),
.B(n_1617),
.Y(n_3081)
);

NOR3xp33_ASAP7_75t_L g3082 ( 
.A(n_2686),
.B(n_1383),
.C(n_1381),
.Y(n_3082)
);

INVxp67_ASAP7_75t_L g3083 ( 
.A(n_2440),
.Y(n_3083)
);

NOR2xp33_ASAP7_75t_L g3084 ( 
.A(n_2518),
.B(n_1618),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2701),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2518),
.B(n_1619),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2408),
.B(n_1625),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2409),
.B(n_1628),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2565),
.Y(n_3089)
);

NOR3xp33_ASAP7_75t_L g3090 ( 
.A(n_2590),
.B(n_1681),
.C(n_1388),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_SL g3091 ( 
.A(n_2617),
.B(n_1629),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2565),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2409),
.B(n_2617),
.Y(n_3093)
);

NOR2xp67_ASAP7_75t_L g3094 ( 
.A(n_2617),
.B(n_2626),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2704),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2626),
.B(n_1634),
.Y(n_3096)
);

INVxp67_ASAP7_75t_SL g3097 ( 
.A(n_2486),
.Y(n_3097)
);

INVxp67_ASAP7_75t_L g3098 ( 
.A(n_2482),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_SL g3099 ( 
.A(n_2626),
.B(n_2711),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2590),
.B(n_1636),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2705),
.Y(n_3101)
);

INVxp67_ASAP7_75t_L g3102 ( 
.A(n_2482),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_SL g3103 ( 
.A(n_2711),
.B(n_1637),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2577),
.B(n_1639),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2577),
.B(n_1640),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_L g3106 ( 
.A(n_2671),
.B(n_1641),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2615),
.B(n_1644),
.Y(n_3107)
);

BUFx6f_ASAP7_75t_SL g3108 ( 
.A(n_2553),
.Y(n_3108)
);

NOR2xp67_ASAP7_75t_L g3109 ( 
.A(n_2615),
.B(n_89),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2629),
.B(n_1645),
.Y(n_3110)
);

A2O1A1Ixp33_ASAP7_75t_L g3111 ( 
.A1(n_2687),
.A2(n_1318),
.B(n_1321),
.C(n_1292),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2629),
.Y(n_3112)
);

NOR3xp33_ASAP7_75t_L g3113 ( 
.A(n_2586),
.B(n_1390),
.C(n_1385),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2555),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2709),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2559),
.B(n_1648),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2710),
.Y(n_3117)
);

NAND2x1p5_ASAP7_75t_L g3118 ( 
.A(n_2734),
.B(n_2740),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2567),
.Y(n_3119)
);

NOR3xp33_ASAP7_75t_L g3120 ( 
.A(n_2681),
.B(n_1397),
.C(n_1395),
.Y(n_3120)
);

BUFx6f_ASAP7_75t_L g3121 ( 
.A(n_2385),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2566),
.B(n_1649),
.Y(n_3122)
);

NOR2xp33_ASAP7_75t_L g3123 ( 
.A(n_2645),
.B(n_1658),
.Y(n_3123)
);

NOR2xp67_ASAP7_75t_L g3124 ( 
.A(n_2405),
.B(n_89),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_SL g3125 ( 
.A(n_2734),
.B(n_1660),
.Y(n_3125)
);

NOR2xp33_ASAP7_75t_L g3126 ( 
.A(n_2406),
.B(n_1661),
.Y(n_3126)
);

NAND3xp33_ASAP7_75t_L g3127 ( 
.A(n_2639),
.B(n_1287),
.C(n_1282),
.Y(n_3127)
);

NAND2xp33_ASAP7_75t_L g3128 ( 
.A(n_2712),
.B(n_1662),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_SL g3129 ( 
.A(n_2740),
.B(n_1663),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2579),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2714),
.B(n_1666),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2580),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2719),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2598),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2721),
.B(n_1667),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2722),
.B(n_1668),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2414),
.B(n_1674),
.Y(n_3137)
);

OR2x6_ASAP7_75t_L g3138 ( 
.A(n_2728),
.B(n_1350),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_2741),
.B(n_1675),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2416),
.B(n_1676),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2741),
.B(n_2730),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2427),
.B(n_2739),
.Y(n_3142)
);

HB1xp67_ASAP7_75t_L g3143 ( 
.A(n_2685),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2746),
.B(n_1677),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2532),
.B(n_1678),
.Y(n_3145)
);

NOR3xp33_ASAP7_75t_L g3146 ( 
.A(n_2681),
.B(n_1419),
.C(n_1398),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2436),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2602),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2534),
.B(n_2537),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_SL g3150 ( 
.A(n_2379),
.B(n_1679),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_R g3151 ( 
.A(n_2682),
.B(n_1683),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2540),
.B(n_1686),
.Y(n_3152)
);

NOR2xp33_ASAP7_75t_L g3153 ( 
.A(n_2682),
.B(n_1687),
.Y(n_3153)
);

OR2x6_ASAP7_75t_L g3154 ( 
.A(n_2380),
.B(n_1350),
.Y(n_3154)
);

INVx3_ASAP7_75t_L g3155 ( 
.A(n_2656),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2384),
.B(n_1689),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2606),
.Y(n_3157)
);

BUFx3_ASAP7_75t_L g3158 ( 
.A(n_2612),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_SL g3159 ( 
.A(n_2397),
.B(n_1690),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_SL g3160 ( 
.A(n_2403),
.B(n_1691),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2404),
.B(n_1692),
.Y(n_3161)
);

NAND3xp33_ASAP7_75t_L g3162 ( 
.A(n_2437),
.B(n_1287),
.C(n_1282),
.Y(n_3162)
);

NAND2xp33_ASAP7_75t_L g3163 ( 
.A(n_2656),
.B(n_1701),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2613),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2438),
.B(n_1693),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2623),
.B(n_1698),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2441),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2627),
.Y(n_3168)
);

BUFx6f_ASAP7_75t_L g3169 ( 
.A(n_2656),
.Y(n_3169)
);

A2O1A1Ixp33_ASAP7_75t_L g3170 ( 
.A1(n_2635),
.A2(n_1409),
.B(n_1429),
.C(n_1408),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2445),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2638),
.B(n_1702),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2651),
.B(n_1421),
.Y(n_3173)
);

INVx2_ASAP7_75t_SL g3174 ( 
.A(n_2652),
.Y(n_3174)
);

AOI221xp5_ASAP7_75t_L g3175 ( 
.A1(n_2661),
.A2(n_1427),
.B1(n_1447),
.B2(n_1444),
.C(n_1430),
.Y(n_3175)
);

INVx3_ASAP7_75t_L g3176 ( 
.A(n_2446),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2449),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2452),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2453),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2662),
.B(n_1460),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2670),
.B(n_1466),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2457),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2674),
.Y(n_3183)
);

AND2x2_ASAP7_75t_L g3184 ( 
.A(n_2675),
.B(n_1469),
.Y(n_3184)
);

NOR2xp33_ASAP7_75t_L g3185 ( 
.A(n_2679),
.B(n_1471),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2460),
.Y(n_3186)
);

INVxp67_ASAP7_75t_SL g3187 ( 
.A(n_2461),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2676),
.B(n_1474),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_2515),
.Y(n_3189)
);

INVx2_ASAP7_75t_SL g3190 ( 
.A(n_2552),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2554),
.B(n_1475),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2412),
.B(n_1479),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_SL g3193 ( 
.A(n_2568),
.B(n_1339),
.Y(n_3193)
);

INVxp67_ASAP7_75t_L g3194 ( 
.A(n_2725),
.Y(n_3194)
);

BUFx6f_ASAP7_75t_L g3195 ( 
.A(n_2368),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2447),
.Y(n_3196)
);

A2O1A1Ixp33_ASAP7_75t_L g3197 ( 
.A1(n_2506),
.A2(n_1409),
.B(n_1429),
.C(n_1408),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_SL g3198 ( 
.A(n_2568),
.B(n_1405),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2412),
.B(n_1490),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2367),
.B(n_1504),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2447),
.Y(n_3201)
);

BUFx6f_ASAP7_75t_L g3202 ( 
.A(n_2368),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_L g3203 ( 
.A(n_2407),
.B(n_1509),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2367),
.B(n_1511),
.Y(n_3204)
);

INVx4_ASAP7_75t_L g3205 ( 
.A(n_2395),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2374),
.Y(n_3206)
);

NOR3xp33_ASAP7_75t_L g3207 ( 
.A(n_2631),
.B(n_1664),
.C(n_1657),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2447),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2367),
.B(n_1519),
.Y(n_3209)
);

NOR2xp67_ASAP7_75t_L g3210 ( 
.A(n_2376),
.B(n_90),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2374),
.Y(n_3211)
);

BUFx5_ASAP7_75t_L g3212 ( 
.A(n_2374),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2367),
.B(n_1527),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2367),
.B(n_1535),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2447),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2412),
.B(n_1538),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2412),
.B(n_1551),
.Y(n_3217)
);

NOR2xp67_ASAP7_75t_L g3218 ( 
.A(n_2376),
.B(n_90),
.Y(n_3218)
);

INVxp67_ASAP7_75t_L g3219 ( 
.A(n_2725),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2412),
.B(n_1558),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2447),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2412),
.B(n_1560),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_2407),
.B(n_1569),
.Y(n_3223)
);

BUFx5_ASAP7_75t_L g3224 ( 
.A(n_2374),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2374),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_SL g3226 ( 
.A(n_2568),
.B(n_1405),
.Y(n_3226)
);

AND2x2_ASAP7_75t_L g3227 ( 
.A(n_2723),
.B(n_1581),
.Y(n_3227)
);

INVx2_ASAP7_75t_SL g3228 ( 
.A(n_2391),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_2374),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2412),
.B(n_1583),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2374),
.Y(n_3231)
);

NOR2xp33_ASAP7_75t_L g3232 ( 
.A(n_2407),
.B(n_1596),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2374),
.Y(n_3233)
);

NOR2xp33_ASAP7_75t_L g3234 ( 
.A(n_2407),
.B(n_1599),
.Y(n_3234)
);

AO221x1_ASAP7_75t_L g3235 ( 
.A1(n_2383),
.A2(n_1308),
.B1(n_1359),
.B2(n_1287),
.C(n_1282),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2447),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_SL g3237 ( 
.A(n_2568),
.B(n_1405),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2374),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2412),
.B(n_1602),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2447),
.Y(n_3240)
);

BUFx6f_ASAP7_75t_L g3241 ( 
.A(n_2368),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_SL g3242 ( 
.A(n_2568),
.B(n_1497),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_2407),
.B(n_1603),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2447),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_SL g3245 ( 
.A(n_2568),
.B(n_1497),
.Y(n_3245)
);

NOR2xp67_ASAP7_75t_L g3246 ( 
.A(n_2376),
.B(n_91),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2447),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_2412),
.B(n_1616),
.Y(n_3248)
);

INVx2_ASAP7_75t_SL g3249 ( 
.A(n_2391),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_SL g3250 ( 
.A(n_2568),
.B(n_1497),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_SL g3251 ( 
.A(n_2459),
.B(n_1497),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2447),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_2447),
.Y(n_3253)
);

INVx2_ASAP7_75t_SL g3254 ( 
.A(n_2391),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_2723),
.B(n_1623),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_2374),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_2412),
.B(n_1624),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_SL g3258 ( 
.A(n_2568),
.B(n_1497),
.Y(n_3258)
);

INVx2_ASAP7_75t_SL g3259 ( 
.A(n_2391),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_2447),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_2412),
.B(n_1626),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2447),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2447),
.Y(n_3263)
);

NOR3xp33_ASAP7_75t_L g3264 ( 
.A(n_2631),
.B(n_1632),
.C(n_1630),
.Y(n_3264)
);

NOR2xp33_ASAP7_75t_L g3265 ( 
.A(n_2407),
.B(n_1638),
.Y(n_3265)
);

INVx2_ASAP7_75t_SL g3266 ( 
.A(n_2391),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_2374),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2447),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_SL g3269 ( 
.A(n_2568),
.B(n_1508),
.Y(n_3269)
);

OR2x6_ASAP7_75t_L g3270 ( 
.A(n_2645),
.B(n_1435),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2447),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_2412),
.B(n_1642),
.Y(n_3272)
);

NOR2xp33_ASAP7_75t_L g3273 ( 
.A(n_2407),
.B(n_1647),
.Y(n_3273)
);

INVx2_ASAP7_75t_L g3274 ( 
.A(n_2374),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_2374),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2412),
.B(n_1650),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_SL g3277 ( 
.A(n_2568),
.B(n_1508),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2412),
.B(n_1651),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2447),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_2412),
.B(n_1652),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2412),
.B(n_1653),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_2412),
.B(n_1656),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2412),
.B(n_1670),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_SL g3284 ( 
.A(n_2568),
.B(n_1508),
.Y(n_3284)
);

NAND2xp33_ASAP7_75t_L g3285 ( 
.A(n_2374),
.B(n_1508),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2412),
.B(n_1671),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2447),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_2412),
.B(n_1673),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2374),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2412),
.B(n_1680),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_2374),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_2412),
.B(n_1508),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_2374),
.Y(n_3293)
);

NOR2xp33_ASAP7_75t_SL g3294 ( 
.A(n_2459),
.B(n_1508),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_2374),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2447),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2447),
.Y(n_3297)
);

BUFx6f_ASAP7_75t_SL g3298 ( 
.A(n_2391),
.Y(n_3298)
);

AND2x6_ASAP7_75t_SL g3299 ( 
.A(n_2411),
.B(n_0),
.Y(n_3299)
);

NAND3xp33_ASAP7_75t_L g3300 ( 
.A(n_2526),
.B(n_1359),
.C(n_1308),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2447),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_2412),
.B(n_1508),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_2568),
.B(n_1572),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_2374),
.Y(n_3304)
);

NOR2xp33_ASAP7_75t_L g3305 ( 
.A(n_2407),
.B(n_1435),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_2407),
.B(n_1442),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2367),
.B(n_1572),
.Y(n_3307)
);

NOR3xp33_ASAP7_75t_L g3308 ( 
.A(n_2631),
.B(n_1446),
.C(n_1442),
.Y(n_3308)
);

NOR2xp33_ASAP7_75t_L g3309 ( 
.A(n_2407),
.B(n_1446),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_2374),
.Y(n_3310)
);

INVxp33_ASAP7_75t_L g3311 ( 
.A(n_2468),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_2374),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_SL g3313 ( 
.A(n_2568),
.B(n_1572),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_2374),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_2374),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_2412),
.B(n_1572),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2447),
.Y(n_3317)
);

OAI22xp5_ASAP7_75t_L g3318 ( 
.A1(n_2374),
.A2(n_1480),
.B1(n_1491),
.B2(n_1461),
.Y(n_3318)
);

BUFx6f_ASAP7_75t_SL g3319 ( 
.A(n_2391),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_SL g3320 ( 
.A(n_2568),
.B(n_1572),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_2374),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_2412),
.B(n_1572),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2412),
.B(n_1572),
.Y(n_3323)
);

OR2x6_ASAP7_75t_L g3324 ( 
.A(n_2645),
.B(n_1461),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_L g3325 ( 
.A(n_2407),
.B(n_1480),
.Y(n_3325)
);

HB1xp67_ASAP7_75t_L g3326 ( 
.A(n_2454),
.Y(n_3326)
);

AOI221xp5_ASAP7_75t_L g3327 ( 
.A1(n_2417),
.A2(n_1563),
.B1(n_1586),
.B2(n_1546),
.C(n_1491),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_SL g3328 ( 
.A(n_2568),
.B(n_1633),
.Y(n_3328)
);

INVxp33_ASAP7_75t_L g3329 ( 
.A(n_2468),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_2374),
.Y(n_3330)
);

NOR2xp33_ASAP7_75t_L g3331 ( 
.A(n_2407),
.B(n_1546),
.Y(n_3331)
);

CKINVDCx5p33_ASAP7_75t_R g3332 ( 
.A(n_2504),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2412),
.B(n_1633),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_2412),
.B(n_1633),
.Y(n_3334)
);

BUFx3_ASAP7_75t_L g3335 ( 
.A(n_2394),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2447),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_2412),
.B(n_1633),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_2412),
.B(n_1633),
.Y(n_3338)
);

INVx2_ASAP7_75t_SL g3339 ( 
.A(n_2391),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2447),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_2447),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_SL g3342 ( 
.A(n_2568),
.B(n_1633),
.Y(n_3342)
);

INVx2_ASAP7_75t_SL g3343 ( 
.A(n_2391),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_2374),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_L g3345 ( 
.A(n_2407),
.B(n_1563),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_2374),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2447),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_2412),
.B(n_1633),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_SL g3349 ( 
.A(n_2568),
.B(n_1654),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_2412),
.B(n_1586),
.Y(n_3350)
);

NOR2xp67_ASAP7_75t_L g3351 ( 
.A(n_2376),
.B(n_92),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_2412),
.B(n_1589),
.Y(n_3352)
);

NAND2xp33_ASAP7_75t_L g3353 ( 
.A(n_2374),
.B(n_1308),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2447),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_2374),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_2568),
.B(n_1654),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_SL g3357 ( 
.A(n_2568),
.B(n_1684),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_2407),
.B(n_1589),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_2412),
.B(n_1684),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_2412),
.B(n_1697),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_2447),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_2447),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2447),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_2374),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_2568),
.B(n_1697),
.Y(n_3365)
);

NOR3xp33_ASAP7_75t_L g3366 ( 
.A(n_2631),
.B(n_1700),
.C(n_85),
.Y(n_3366)
);

INVx2_ASAP7_75t_SL g3367 ( 
.A(n_2391),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_2412),
.B(n_1700),
.Y(n_3368)
);

NAND3xp33_ASAP7_75t_L g3369 ( 
.A(n_2526),
.B(n_1359),
.C(n_1308),
.Y(n_3369)
);

AO221x1_ASAP7_75t_L g3370 ( 
.A1(n_2383),
.A2(n_1443),
.B1(n_1459),
.B2(n_1439),
.C(n_1359),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_2407),
.B(n_84),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_2367),
.B(n_1439),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_2367),
.B(n_1439),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_2374),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_2367),
.B(n_1439),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_2367),
.B(n_1443),
.Y(n_3376)
);

NOR2xp33_ASAP7_75t_L g3377 ( 
.A(n_2407),
.B(n_84),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_2374),
.Y(n_3378)
);

NOR2xp33_ASAP7_75t_L g3379 ( 
.A(n_2407),
.B(n_85),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_2407),
.A2(n_1459),
.B1(n_1477),
.B2(n_1443),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2447),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_SL g3382 ( 
.A(n_2568),
.B(n_1443),
.Y(n_3382)
);

INVx8_ASAP7_75t_L g3383 ( 
.A(n_2411),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2447),
.Y(n_3384)
);

NOR2xp33_ASAP7_75t_L g3385 ( 
.A(n_2407),
.B(n_85),
.Y(n_3385)
);

NOR2xp33_ASAP7_75t_L g3386 ( 
.A(n_2407),
.B(n_86),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2447),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_2568),
.B(n_1459),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_2447),
.Y(n_3389)
);

NOR2xp67_ASAP7_75t_L g3390 ( 
.A(n_2376),
.B(n_94),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_2766),
.Y(n_3391)
);

NAND2x1p5_ASAP7_75t_L g3392 ( 
.A(n_2751),
.B(n_1459),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2770),
.Y(n_3393)
);

AO22x2_ASAP7_75t_L g3394 ( 
.A1(n_3318),
.A2(n_87),
.B1(n_88),
.B2(n_86),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_2756),
.B(n_86),
.Y(n_3395)
);

BUFx2_ASAP7_75t_L g3396 ( 
.A(n_2965),
.Y(n_3396)
);

NAND2x1p5_ASAP7_75t_L g3397 ( 
.A(n_2751),
.B(n_1477),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2843),
.Y(n_3398)
);

INVxp67_ASAP7_75t_L g3399 ( 
.A(n_3326),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_2805),
.B(n_2814),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_2776),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3227),
.B(n_87),
.Y(n_3402)
);

OAI22xp5_ASAP7_75t_L g3403 ( 
.A1(n_2860),
.A2(n_1579),
.B1(n_1621),
.B2(n_1477),
.Y(n_3403)
);

OAI221xp5_ASAP7_75t_L g3404 ( 
.A1(n_2842),
.A2(n_1621),
.B1(n_1635),
.B2(n_1579),
.C(n_1477),
.Y(n_3404)
);

NAND3xp33_ASAP7_75t_SL g3405 ( 
.A(n_3151),
.B(n_1),
.C(n_2),
.Y(n_3405)
);

NAND2x1p5_ASAP7_75t_L g3406 ( 
.A(n_3021),
.B(n_1579),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2848),
.Y(n_3407)
);

AOI22xp5_ASAP7_75t_L g3408 ( 
.A1(n_2808),
.A2(n_1621),
.B1(n_1635),
.B2(n_1579),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_2898),
.Y(n_3409)
);

INVx3_ASAP7_75t_L g3410 ( 
.A(n_2967),
.Y(n_3410)
);

HB1xp67_ASAP7_75t_L g3411 ( 
.A(n_3270),
.Y(n_3411)
);

INVx2_ASAP7_75t_SL g3412 ( 
.A(n_2967),
.Y(n_3412)
);

AOI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_2812),
.A2(n_1635),
.B1(n_1669),
.B2(n_1621),
.Y(n_3413)
);

INVx3_ASAP7_75t_L g3414 ( 
.A(n_2967),
.Y(n_3414)
);

NAND2x1p5_ASAP7_75t_L g3415 ( 
.A(n_3021),
.B(n_1635),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2749),
.Y(n_3416)
);

NAND2x1p5_ASAP7_75t_L g3417 ( 
.A(n_3066),
.B(n_1669),
.Y(n_3417)
);

NOR2xp33_ASAP7_75t_L g3418 ( 
.A(n_2754),
.B(n_87),
.Y(n_3418)
);

AO22x2_ASAP7_75t_L g3419 ( 
.A1(n_3318),
.A2(n_91),
.B1(n_92),
.B2(n_88),
.Y(n_3419)
);

A2O1A1Ixp33_ASAP7_75t_L g3420 ( 
.A1(n_3371),
.A2(n_1669),
.B(n_3),
.C(n_1),
.Y(n_3420)
);

AOI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_2767),
.A2(n_1669),
.B1(n_92),
.B2(n_93),
.Y(n_3421)
);

NAND2x1p5_ASAP7_75t_L g3422 ( 
.A(n_3066),
.B(n_91),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_2755),
.Y(n_3423)
);

NAND2x1p5_ASAP7_75t_L g3424 ( 
.A(n_3023),
.B(n_93),
.Y(n_3424)
);

NOR2xp33_ASAP7_75t_L g3425 ( 
.A(n_3311),
.B(n_94),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3255),
.B(n_94),
.Y(n_3426)
);

BUFx6f_ASAP7_75t_L g3427 ( 
.A(n_2786),
.Y(n_3427)
);

NAND3xp33_ASAP7_75t_SL g3428 ( 
.A(n_2798),
.B(n_2821),
.C(n_3366),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2768),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3196),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3206),
.Y(n_3431)
);

OAI221xp5_ASAP7_75t_L g3432 ( 
.A1(n_3203),
.A2(n_3232),
.B1(n_3243),
.B2(n_3234),
.C(n_3223),
.Y(n_3432)
);

HB1xp67_ASAP7_75t_L g3433 ( 
.A(n_3270),
.Y(n_3433)
);

AO22x2_ASAP7_75t_L g3434 ( 
.A1(n_2949),
.A2(n_96),
.B1(n_97),
.B2(n_95),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3201),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3208),
.Y(n_3436)
);

AOI22xp5_ASAP7_75t_L g3437 ( 
.A1(n_2931),
.A2(n_96),
.B1(n_97),
.B2(n_95),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3215),
.Y(n_3438)
);

AO22x2_ASAP7_75t_L g3439 ( 
.A1(n_2761),
.A2(n_97),
.B1(n_98),
.B2(n_95),
.Y(n_3439)
);

INVx3_ASAP7_75t_L g3440 ( 
.A(n_3108),
.Y(n_3440)
);

BUFx8_ASAP7_75t_L g3441 ( 
.A(n_3108),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3221),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3236),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_SL g3444 ( 
.A(n_3008),
.B(n_98),
.Y(n_3444)
);

AOI22xp5_ASAP7_75t_L g3445 ( 
.A1(n_2817),
.A2(n_99),
.B1(n_100),
.B2(n_98),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3211),
.Y(n_3446)
);

INVx3_ASAP7_75t_L g3447 ( 
.A(n_2849),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3240),
.Y(n_3448)
);

AO22x2_ASAP7_75t_L g3449 ( 
.A1(n_3194),
.A2(n_100),
.B1(n_101),
.B2(n_99),
.Y(n_3449)
);

NAND2x1p5_ASAP7_75t_L g3450 ( 
.A(n_2921),
.B(n_99),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_R g3451 ( 
.A(n_2804),
.B(n_2),
.Y(n_3451)
);

BUFx6f_ASAP7_75t_SL g3452 ( 
.A(n_2915),
.Y(n_3452)
);

AO22x2_ASAP7_75t_L g3453 ( 
.A1(n_3219),
.A2(n_102),
.B1(n_103),
.B2(n_101),
.Y(n_3453)
);

INVx3_ASAP7_75t_L g3454 ( 
.A(n_2849),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3244),
.Y(n_3455)
);

AO22x2_ASAP7_75t_L g3456 ( 
.A1(n_2870),
.A2(n_104),
.B1(n_105),
.B2(n_103),
.Y(n_3456)
);

OAI221xp5_ASAP7_75t_L g3457 ( 
.A1(n_3265),
.A2(n_3273),
.B1(n_3078),
.B2(n_2826),
.C(n_3082),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3225),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3247),
.Y(n_3459)
);

CKINVDCx20_ASAP7_75t_R g3460 ( 
.A(n_3332),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3252),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3229),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_3329),
.B(n_104),
.Y(n_3463)
);

INVxp67_ASAP7_75t_L g3464 ( 
.A(n_2772),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3253),
.Y(n_3465)
);

AO22x2_ASAP7_75t_L g3466 ( 
.A1(n_2824),
.A2(n_107),
.B1(n_108),
.B2(n_106),
.Y(n_3466)
);

OAI221xp5_ASAP7_75t_L g3467 ( 
.A1(n_3207),
.A2(n_108),
.B1(n_109),
.B2(n_107),
.C(n_106),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3260),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_2760),
.B(n_106),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3262),
.Y(n_3470)
);

AND2x4_ASAP7_75t_L g3471 ( 
.A(n_2915),
.B(n_107),
.Y(n_3471)
);

AO22x2_ASAP7_75t_L g3472 ( 
.A1(n_2828),
.A2(n_109),
.B1(n_110),
.B2(n_108),
.Y(n_3472)
);

OAI221xp5_ASAP7_75t_L g3473 ( 
.A1(n_3264),
.A2(n_112),
.B1(n_113),
.B2(n_111),
.C(n_110),
.Y(n_3473)
);

AOI22xp5_ASAP7_75t_L g3474 ( 
.A1(n_3025),
.A2(n_112),
.B1(n_113),
.B2(n_111),
.Y(n_3474)
);

INVxp67_ASAP7_75t_L g3475 ( 
.A(n_2939),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3263),
.Y(n_3476)
);

AO22x2_ASAP7_75t_L g3477 ( 
.A1(n_2834),
.A2(n_114),
.B1(n_115),
.B2(n_113),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3268),
.Y(n_3478)
);

INVxp67_ASAP7_75t_L g3479 ( 
.A(n_3270),
.Y(n_3479)
);

INVxp67_ASAP7_75t_L g3480 ( 
.A(n_3324),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3231),
.Y(n_3481)
);

CKINVDCx20_ASAP7_75t_R g3482 ( 
.A(n_2835),
.Y(n_3482)
);

AND2x6_ASAP7_75t_L g3483 ( 
.A(n_2765),
.B(n_114),
.Y(n_3483)
);

AND2x4_ASAP7_75t_L g3484 ( 
.A(n_2915),
.B(n_115),
.Y(n_3484)
);

NAND2x1p5_ASAP7_75t_L g3485 ( 
.A(n_3094),
.B(n_115),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3271),
.Y(n_3486)
);

AO22x2_ASAP7_75t_L g3487 ( 
.A1(n_2840),
.A2(n_117),
.B1(n_118),
.B2(n_116),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_2866),
.B(n_116),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3279),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3287),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3296),
.Y(n_3491)
);

AO22x2_ASAP7_75t_L g3492 ( 
.A1(n_2859),
.A2(n_118),
.B1(n_119),
.B2(n_117),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3297),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3301),
.Y(n_3494)
);

AO22x2_ASAP7_75t_L g3495 ( 
.A1(n_2864),
.A2(n_118),
.B1(n_119),
.B2(n_117),
.Y(n_3495)
);

BUFx6f_ASAP7_75t_SL g3496 ( 
.A(n_3324),
.Y(n_3496)
);

AO22x2_ASAP7_75t_L g3497 ( 
.A1(n_2867),
.A2(n_120),
.B1(n_121),
.B2(n_119),
.Y(n_3497)
);

AO22x2_ASAP7_75t_L g3498 ( 
.A1(n_2868),
.A2(n_121),
.B1(n_122),
.B2(n_120),
.Y(n_3498)
);

AND2x4_ASAP7_75t_L g3499 ( 
.A(n_3324),
.B(n_122),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3233),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3238),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3317),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3336),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3340),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_2927),
.B(n_122),
.Y(n_3505)
);

AO22x2_ASAP7_75t_L g3506 ( 
.A1(n_2883),
.A2(n_124),
.B1(n_125),
.B2(n_123),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3256),
.Y(n_3507)
);

AOI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3377),
.A2(n_124),
.B1(n_125),
.B2(n_123),
.Y(n_3508)
);

BUFx12f_ASAP7_75t_L g3509 ( 
.A(n_3036),
.Y(n_3509)
);

AO22x2_ASAP7_75t_L g3510 ( 
.A1(n_2778),
.A2(n_126),
.B1(n_127),
.B2(n_124),
.Y(n_3510)
);

NAND2x1p5_ASAP7_75t_L g3511 ( 
.A(n_3205),
.B(n_2792),
.Y(n_3511)
);

NAND2x1p5_ASAP7_75t_L g3512 ( 
.A(n_3205),
.B(n_126),
.Y(n_3512)
);

OAI221xp5_ASAP7_75t_L g3513 ( 
.A1(n_2809),
.A2(n_128),
.B1(n_129),
.B2(n_127),
.C(n_126),
.Y(n_3513)
);

AND2x4_ASAP7_75t_L g3514 ( 
.A(n_2926),
.B(n_127),
.Y(n_3514)
);

NAND3x1_ASAP7_75t_L g3515 ( 
.A(n_3079),
.B(n_1063),
.C(n_1062),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3341),
.Y(n_3516)
);

OAI221xp5_ASAP7_75t_L g3517 ( 
.A1(n_3305),
.A2(n_130),
.B1(n_131),
.B2(n_129),
.C(n_128),
.Y(n_3517)
);

AO22x2_ASAP7_75t_L g3518 ( 
.A1(n_2787),
.A2(n_130),
.B1(n_131),
.B2(n_128),
.Y(n_3518)
);

NAND3xp33_ASAP7_75t_SL g3519 ( 
.A(n_3327),
.B(n_1),
.C(n_2),
.Y(n_3519)
);

INVx3_ASAP7_75t_L g3520 ( 
.A(n_2906),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3267),
.Y(n_3521)
);

NAND2x1_ASAP7_75t_L g3522 ( 
.A(n_3274),
.B(n_131),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_2899),
.B(n_2957),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3347),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_2927),
.B(n_132),
.Y(n_3525)
);

AO22x2_ASAP7_75t_L g3526 ( 
.A1(n_2790),
.A2(n_133),
.B1(n_134),
.B2(n_132),
.Y(n_3526)
);

NAND2x1p5_ASAP7_75t_L g3527 ( 
.A(n_3335),
.B(n_133),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_2917),
.B(n_134),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3354),
.Y(n_3529)
);

AO22x2_ASAP7_75t_L g3530 ( 
.A1(n_2813),
.A2(n_135),
.B1(n_136),
.B2(n_134),
.Y(n_3530)
);

AO22x1_ASAP7_75t_L g3531 ( 
.A1(n_2815),
.A2(n_1070),
.B1(n_1071),
.B2(n_1069),
.Y(n_3531)
);

AND2x4_ASAP7_75t_L g3532 ( 
.A(n_2852),
.B(n_135),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3275),
.Y(n_3533)
);

AO22x2_ASAP7_75t_L g3534 ( 
.A1(n_2837),
.A2(n_136),
.B1(n_137),
.B2(n_135),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3289),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3361),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3362),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3363),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3381),
.Y(n_3539)
);

AOI22xp5_ASAP7_75t_L g3540 ( 
.A1(n_3379),
.A2(n_3386),
.B1(n_3385),
.B2(n_2779),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3384),
.Y(n_3541)
);

AND2x4_ASAP7_75t_L g3542 ( 
.A(n_2971),
.B(n_137),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3387),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3389),
.Y(n_3544)
);

AND2x4_ASAP7_75t_L g3545 ( 
.A(n_3228),
.B(n_138),
.Y(n_3545)
);

NOR2xp67_ASAP7_75t_L g3546 ( 
.A(n_3098),
.B(n_138),
.Y(n_3546)
);

AND2x4_ASAP7_75t_L g3547 ( 
.A(n_3249),
.B(n_139),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_2853),
.Y(n_3548)
);

AO22x2_ASAP7_75t_L g3549 ( 
.A1(n_2851),
.A2(n_140),
.B1(n_141),
.B2(n_139),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_2928),
.B(n_2938),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3291),
.Y(n_3551)
);

OAI221xp5_ASAP7_75t_L g3552 ( 
.A1(n_3306),
.A2(n_141),
.B1(n_142),
.B2(n_140),
.C(n_139),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_2871),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3293),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_2819),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3295),
.Y(n_3556)
);

AOI22xp5_ASAP7_75t_L g3557 ( 
.A1(n_2963),
.A2(n_142),
.B1(n_143),
.B2(n_141),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_2823),
.Y(n_3558)
);

CKINVDCx20_ASAP7_75t_R g3559 ( 
.A(n_2987),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_2830),
.Y(n_3560)
);

INVx2_ASAP7_75t_SL g3561 ( 
.A(n_3383),
.Y(n_3561)
);

NAND2x1p5_ASAP7_75t_L g3562 ( 
.A(n_3254),
.B(n_142),
.Y(n_3562)
);

AO22x2_ASAP7_75t_L g3563 ( 
.A1(n_2777),
.A2(n_144),
.B1(n_145),
.B2(n_143),
.Y(n_3563)
);

BUFx6f_ASAP7_75t_SL g3564 ( 
.A(n_3259),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_2836),
.Y(n_3565)
);

INVx4_ASAP7_75t_L g3566 ( 
.A(n_2906),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_2928),
.B(n_144),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_2839),
.Y(n_3568)
);

OAI221xp5_ASAP7_75t_L g3569 ( 
.A1(n_3309),
.A2(n_147),
.B1(n_148),
.B2(n_146),
.C(n_145),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_SL g3570 ( 
.A(n_3008),
.B(n_145),
.Y(n_3570)
);

NAND2x1p5_ASAP7_75t_L g3571 ( 
.A(n_3266),
.B(n_146),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_2875),
.Y(n_3572)
);

OAI22xp5_ASAP7_75t_SL g3573 ( 
.A1(n_3080),
.A2(n_2879),
.B1(n_2935),
.B2(n_2781),
.Y(n_3573)
);

AO22x2_ASAP7_75t_L g3574 ( 
.A1(n_2784),
.A2(n_147),
.B1(n_148),
.B2(n_146),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_2876),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_2884),
.Y(n_3576)
);

INVxp67_ASAP7_75t_L g3577 ( 
.A(n_2912),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_2889),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_2890),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_2896),
.Y(n_3580)
);

INVxp67_ASAP7_75t_L g3581 ( 
.A(n_2829),
.Y(n_3581)
);

AO22x2_ASAP7_75t_L g3582 ( 
.A1(n_2789),
.A2(n_149),
.B1(n_150),
.B2(n_148),
.Y(n_3582)
);

CKINVDCx20_ASAP7_75t_R g3583 ( 
.A(n_3143),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_2902),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_2913),
.Y(n_3585)
);

AND2x4_ASAP7_75t_L g3586 ( 
.A(n_3339),
.B(n_149),
.Y(n_3586)
);

OR2x6_ASAP7_75t_L g3587 ( 
.A(n_3383),
.B(n_150),
.Y(n_3587)
);

OAI221xp5_ASAP7_75t_L g3588 ( 
.A1(n_3325),
.A2(n_152),
.B1(n_153),
.B2(n_151),
.C(n_150),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_2916),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_2944),
.Y(n_3590)
);

INVxp67_ASAP7_75t_L g3591 ( 
.A(n_2937),
.Y(n_3591)
);

NAND2x1p5_ASAP7_75t_L g3592 ( 
.A(n_3343),
.B(n_3367),
.Y(n_3592)
);

AO22x2_ASAP7_75t_L g3593 ( 
.A1(n_2791),
.A2(n_152),
.B1(n_154),
.B2(n_151),
.Y(n_3593)
);

CKINVDCx20_ASAP7_75t_R g3594 ( 
.A(n_3383),
.Y(n_3594)
);

AOI22xp33_ASAP7_75t_L g3595 ( 
.A1(n_3090),
.A2(n_152),
.B1(n_154),
.B2(n_151),
.Y(n_3595)
);

BUFx8_ASAP7_75t_L g3596 ( 
.A(n_3298),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_2873),
.B(n_154),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_2922),
.Y(n_3598)
);

NAND2x1p5_ASAP7_75t_L g3599 ( 
.A(n_2765),
.B(n_155),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_2938),
.B(n_155),
.Y(n_3600)
);

OAI221xp5_ASAP7_75t_L g3601 ( 
.A1(n_3331),
.A2(n_157),
.B1(n_158),
.B2(n_156),
.C(n_155),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_2929),
.Y(n_3602)
);

HB1xp67_ASAP7_75t_L g3603 ( 
.A(n_2880),
.Y(n_3603)
);

AO22x2_ASAP7_75t_L g3604 ( 
.A1(n_2795),
.A2(n_157),
.B1(n_158),
.B2(n_156),
.Y(n_3604)
);

OR2x2_ASAP7_75t_SL g3605 ( 
.A(n_3069),
.B(n_157),
.Y(n_3605)
);

OAI221xp5_ASAP7_75t_L g3606 ( 
.A1(n_3345),
.A2(n_161),
.B1(n_162),
.B2(n_160),
.C(n_159),
.Y(n_3606)
);

NOR2xp33_ASAP7_75t_L g3607 ( 
.A(n_3052),
.B(n_2969),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_2930),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3006),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3013),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_2802),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3304),
.Y(n_3612)
);

NAND2x1p5_ASAP7_75t_L g3613 ( 
.A(n_2825),
.B(n_159),
.Y(n_3613)
);

INVx2_ASAP7_75t_L g3614 ( 
.A(n_3310),
.Y(n_3614)
);

NAND2x1p5_ASAP7_75t_L g3615 ( 
.A(n_2825),
.B(n_3032),
.Y(n_3615)
);

AO22x2_ASAP7_75t_L g3616 ( 
.A1(n_3312),
.A2(n_160),
.B1(n_161),
.B2(n_159),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_2954),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_2955),
.Y(n_3618)
);

INVx2_ASAP7_75t_SL g3619 ( 
.A(n_2858),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_2986),
.Y(n_3620)
);

NAND2x1p5_ASAP7_75t_L g3621 ( 
.A(n_3298),
.B(n_161),
.Y(n_3621)
);

CKINVDCx16_ASAP7_75t_R g3622 ( 
.A(n_3319),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_2985),
.B(n_162),
.Y(n_3623)
);

AND2x6_ASAP7_75t_L g3624 ( 
.A(n_3314),
.B(n_163),
.Y(n_3624)
);

OAI22xp5_ASAP7_75t_SL g3625 ( 
.A1(n_3299),
.A2(n_164),
.B1(n_165),
.B2(n_163),
.Y(n_3625)
);

AND2x2_ASAP7_75t_L g3626 ( 
.A(n_2980),
.B(n_163),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_2996),
.Y(n_3627)
);

NAND2x1p5_ASAP7_75t_L g3628 ( 
.A(n_3319),
.B(n_165),
.Y(n_3628)
);

AND2x2_ASAP7_75t_L g3629 ( 
.A(n_3358),
.B(n_165),
.Y(n_3629)
);

OAI221xp5_ASAP7_75t_L g3630 ( 
.A1(n_2759),
.A2(n_168),
.B1(n_169),
.B2(n_167),
.C(n_166),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3000),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3003),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3011),
.Y(n_3633)
);

AO22x2_ASAP7_75t_L g3634 ( 
.A1(n_3315),
.A2(n_168),
.B1(n_169),
.B2(n_167),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3012),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3016),
.Y(n_3636)
);

CKINVDCx5p33_ASAP7_75t_R g3637 ( 
.A(n_2816),
.Y(n_3637)
);

CKINVDCx5p33_ASAP7_75t_R g3638 ( 
.A(n_2984),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_2983),
.B(n_2989),
.Y(n_3639)
);

AO22x2_ASAP7_75t_L g3640 ( 
.A1(n_3321),
.A2(n_3330),
.B1(n_3346),
.B2(n_3344),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3355),
.Y(n_3641)
);

AO22x2_ASAP7_75t_L g3642 ( 
.A1(n_3364),
.A2(n_170),
.B1(n_171),
.B2(n_168),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3184),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3173),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3374),
.Y(n_3645)
);

AO22x2_ASAP7_75t_L g3646 ( 
.A1(n_3378),
.A2(n_2801),
.B1(n_2895),
.B2(n_2983),
.Y(n_3646)
);

BUFx3_ASAP7_75t_L g3647 ( 
.A(n_2822),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3173),
.Y(n_3648)
);

AND2x4_ASAP7_75t_L g3649 ( 
.A(n_3102),
.B(n_170),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_2940),
.Y(n_3650)
);

NAND3x1_ASAP7_75t_L g3651 ( 
.A(n_3072),
.B(n_1074),
.C(n_1073),
.Y(n_3651)
);

AND2x4_ASAP7_75t_L g3652 ( 
.A(n_2968),
.B(n_170),
.Y(n_3652)
);

BUFx8_ASAP7_75t_L g3653 ( 
.A(n_2822),
.Y(n_3653)
);

OR2x2_ASAP7_75t_L g3654 ( 
.A(n_2966),
.B(n_2972),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_2942),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3212),
.Y(n_3656)
);

INVx3_ASAP7_75t_L g3657 ( 
.A(n_3158),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_2999),
.B(n_172),
.Y(n_3658)
);

OR2x6_ASAP7_75t_L g3659 ( 
.A(n_3083),
.B(n_172),
.Y(n_3659)
);

NOR2xp67_ASAP7_75t_L g3660 ( 
.A(n_3123),
.B(n_173),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_2811),
.B(n_173),
.Y(n_3661)
);

AND2x2_ASAP7_75t_L g3662 ( 
.A(n_2998),
.B(n_173),
.Y(n_3662)
);

AND2x4_ASAP7_75t_L g3663 ( 
.A(n_2832),
.B(n_174),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_SL g3664 ( 
.A(n_3008),
.B(n_174),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3004),
.B(n_174),
.Y(n_3665)
);

NAND2x1p5_ASAP7_75t_L g3666 ( 
.A(n_3070),
.B(n_3055),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_2947),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_SL g3668 ( 
.A(n_3008),
.B(n_175),
.Y(n_3668)
);

CKINVDCx5p33_ASAP7_75t_R g3669 ( 
.A(n_3106),
.Y(n_3669)
);

INVx4_ASAP7_75t_L g3670 ( 
.A(n_3008),
.Y(n_3670)
);

AO22x2_ASAP7_75t_L g3671 ( 
.A1(n_2874),
.A2(n_176),
.B1(n_177),
.B2(n_175),
.Y(n_3671)
);

NOR2xp33_ASAP7_75t_L g3672 ( 
.A(n_2862),
.B(n_2793),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_2952),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_2953),
.Y(n_3674)
);

BUFx2_ASAP7_75t_L g3675 ( 
.A(n_3154),
.Y(n_3675)
);

A2O1A1Ixp33_ASAP7_75t_L g3676 ( 
.A1(n_3020),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3212),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_2979),
.Y(n_3678)
);

AND2x4_ASAP7_75t_L g3679 ( 
.A(n_2970),
.B(n_175),
.Y(n_3679)
);

BUFx2_ASAP7_75t_L g3680 ( 
.A(n_3154),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_L g3681 ( 
.A1(n_2936),
.A2(n_177),
.B1(n_178),
.B2(n_176),
.Y(n_3681)
);

AO22x2_ASAP7_75t_L g3682 ( 
.A1(n_2959),
.A2(n_2958),
.B1(n_3146),
.B2(n_3120),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3048),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3181),
.Y(n_3684)
);

INVxp33_ASAP7_75t_SL g3685 ( 
.A(n_2758),
.Y(n_3685)
);

OAI221xp5_ASAP7_75t_L g3686 ( 
.A1(n_2981),
.A2(n_3057),
.B1(n_2752),
.B2(n_2753),
.C(n_2897),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3019),
.B(n_177),
.Y(n_3687)
);

CKINVDCx5p33_ASAP7_75t_R g3688 ( 
.A(n_2941),
.Y(n_3688)
);

NOR2xp67_ASAP7_75t_L g3689 ( 
.A(n_3001),
.B(n_178),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3188),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3002),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_2762),
.B(n_178),
.Y(n_3692)
);

AO22x2_ASAP7_75t_L g3693 ( 
.A1(n_3014),
.A2(n_180),
.B1(n_182),
.B2(n_179),
.Y(n_3693)
);

INVx4_ASAP7_75t_L g3694 ( 
.A(n_3154),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_2844),
.B(n_179),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3212),
.Y(n_3696)
);

CKINVDCx20_ASAP7_75t_R g3697 ( 
.A(n_2799),
.Y(n_3697)
);

NAND2x1p5_ASAP7_75t_L g3698 ( 
.A(n_3081),
.B(n_2748),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3200),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3200),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3204),
.Y(n_3701)
);

INVxp67_ASAP7_75t_L g3702 ( 
.A(n_2945),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_2762),
.B(n_179),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3204),
.Y(n_3704)
);

CKINVDCx5p33_ASAP7_75t_R g3705 ( 
.A(n_3122),
.Y(n_3705)
);

AO22x2_ASAP7_75t_L g3706 ( 
.A1(n_2763),
.A2(n_182),
.B1(n_183),
.B2(n_180),
.Y(n_3706)
);

OR2x2_ASAP7_75t_SL g3707 ( 
.A(n_3116),
.B(n_180),
.Y(n_3707)
);

HB1xp67_ASAP7_75t_L g3708 ( 
.A(n_3035),
.Y(n_3708)
);

CKINVDCx20_ASAP7_75t_R g3709 ( 
.A(n_2807),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_2847),
.B(n_182),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3209),
.Y(n_3711)
);

NAND2x1p5_ASAP7_75t_L g3712 ( 
.A(n_2748),
.B(n_183),
.Y(n_3712)
);

INVx2_ASAP7_75t_SL g3713 ( 
.A(n_2977),
.Y(n_3713)
);

INVx3_ASAP7_75t_L g3714 ( 
.A(n_3017),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3209),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3213),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3213),
.Y(n_3717)
);

AO22x2_ASAP7_75t_L g3718 ( 
.A1(n_2763),
.A2(n_184),
.B1(n_185),
.B2(n_183),
.Y(n_3718)
);

AO22x2_ASAP7_75t_L g3719 ( 
.A1(n_2774),
.A2(n_185),
.B1(n_186),
.B2(n_184),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3214),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_2774),
.B(n_184),
.Y(n_3721)
);

AO22x2_ASAP7_75t_L g3722 ( 
.A1(n_2775),
.A2(n_186),
.B1(n_187),
.B2(n_185),
.Y(n_3722)
);

OR2x6_ASAP7_75t_L g3723 ( 
.A(n_2764),
.B(n_186),
.Y(n_3723)
);

AO22x2_ASAP7_75t_L g3724 ( 
.A1(n_2775),
.A2(n_188),
.B1(n_189),
.B2(n_187),
.Y(n_3724)
);

NAND2x1p5_ASAP7_75t_L g3725 ( 
.A(n_2748),
.B(n_188),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3212),
.Y(n_3726)
);

AOI22xp5_ASAP7_75t_L g3727 ( 
.A1(n_2818),
.A2(n_190),
.B1(n_191),
.B2(n_189),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_2783),
.B(n_189),
.Y(n_3728)
);

HB1xp67_ASAP7_75t_L g3729 ( 
.A(n_3138),
.Y(n_3729)
);

AND2x2_ASAP7_75t_L g3730 ( 
.A(n_2905),
.B(n_190),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3214),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3372),
.Y(n_3732)
);

OAI22xp5_ASAP7_75t_L g3733 ( 
.A1(n_3138),
.A2(n_191),
.B1(n_192),
.B2(n_190),
.Y(n_3733)
);

AO22x2_ASAP7_75t_L g3734 ( 
.A1(n_2783),
.A2(n_192),
.B1(n_193),
.B2(n_191),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3372),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_2918),
.B(n_193),
.Y(n_3736)
);

AOI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_2856),
.A2(n_194),
.B1(n_195),
.B2(n_193),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3373),
.Y(n_3738)
);

AND2x4_ASAP7_75t_L g3739 ( 
.A(n_2992),
.B(n_194),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3373),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3192),
.B(n_194),
.Y(n_3741)
);

AO22x2_ASAP7_75t_L g3742 ( 
.A1(n_3308),
.A2(n_2956),
.B1(n_2950),
.B2(n_3382),
.Y(n_3742)
);

OAI221xp5_ASAP7_75t_L g3743 ( 
.A1(n_3199),
.A2(n_197),
.B1(n_198),
.B2(n_196),
.C(n_195),
.Y(n_3743)
);

BUFx6f_ASAP7_75t_SL g3744 ( 
.A(n_3033),
.Y(n_3744)
);

NAND2xp33_ASAP7_75t_L g3745 ( 
.A(n_2990),
.B(n_195),
.Y(n_3745)
);

AO22x2_ASAP7_75t_L g3746 ( 
.A1(n_3388),
.A2(n_197),
.B1(n_198),
.B2(n_196),
.Y(n_3746)
);

HB1xp67_ASAP7_75t_L g3747 ( 
.A(n_3138),
.Y(n_3747)
);

BUFx2_ASAP7_75t_L g3748 ( 
.A(n_3212),
.Y(n_3748)
);

INVxp67_ASAP7_75t_L g3749 ( 
.A(n_2861),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3375),
.Y(n_3750)
);

AOI22xp5_ASAP7_75t_L g3751 ( 
.A1(n_3153),
.A2(n_197),
.B1(n_199),
.B2(n_196),
.Y(n_3751)
);

A2O1A1Ixp33_ASAP7_75t_L g3752 ( 
.A1(n_3353),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3224),
.Y(n_3753)
);

OAI221xp5_ASAP7_75t_L g3754 ( 
.A1(n_3216),
.A2(n_201),
.B1(n_202),
.B2(n_200),
.C(n_199),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3375),
.Y(n_3755)
);

INVxp67_ASAP7_75t_L g3756 ( 
.A(n_3084),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3217),
.B(n_199),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3376),
.Y(n_3758)
);

AND2x2_ASAP7_75t_L g3759 ( 
.A(n_2865),
.B(n_200),
.Y(n_3759)
);

OR2x6_ASAP7_75t_L g3760 ( 
.A(n_2769),
.B(n_201),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3376),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3030),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_2946),
.B(n_201),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3045),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_3224),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_2951),
.B(n_202),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3307),
.Y(n_3767)
);

AO22x2_ASAP7_75t_L g3768 ( 
.A1(n_2882),
.A2(n_203),
.B1(n_204),
.B2(n_202),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3224),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3224),
.Y(n_3770)
);

HB1xp67_ASAP7_75t_L g3771 ( 
.A(n_3124),
.Y(n_3771)
);

INVxp67_ASAP7_75t_L g3772 ( 
.A(n_2961),
.Y(n_3772)
);

AO22x2_ASAP7_75t_L g3773 ( 
.A1(n_3113),
.A2(n_204),
.B1(n_205),
.B2(n_203),
.Y(n_3773)
);

AO22x2_ASAP7_75t_L g3774 ( 
.A1(n_3034),
.A2(n_205),
.B1(n_206),
.B2(n_204),
.Y(n_3774)
);

AOI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_3058),
.A2(n_3076),
.B1(n_2964),
.B2(n_2907),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3307),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3224),
.Y(n_3777)
);

CKINVDCx5p33_ASAP7_75t_R g3778 ( 
.A(n_2806),
.Y(n_3778)
);

NAND2x1p5_ASAP7_75t_L g3779 ( 
.A(n_2750),
.B(n_205),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3220),
.B(n_206),
.Y(n_3780)
);

AO22x2_ASAP7_75t_L g3781 ( 
.A1(n_3065),
.A2(n_208),
.B1(n_209),
.B2(n_207),
.Y(n_3781)
);

AO22x2_ASAP7_75t_L g3782 ( 
.A1(n_3067),
.A2(n_208),
.B1(n_209),
.B2(n_207),
.Y(n_3782)
);

CKINVDCx5p33_ASAP7_75t_R g3783 ( 
.A(n_2886),
.Y(n_3783)
);

BUFx8_ASAP7_75t_L g3784 ( 
.A(n_3027),
.Y(n_3784)
);

AOI22xp5_ASAP7_75t_L g3785 ( 
.A1(n_2900),
.A2(n_211),
.B1(n_212),
.B2(n_210),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3114),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_2903),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3119),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3130),
.Y(n_3789)
);

BUFx8_ASAP7_75t_L g3790 ( 
.A(n_3026),
.Y(n_3790)
);

AO22x2_ASAP7_75t_L g3791 ( 
.A1(n_3071),
.A2(n_211),
.B1(n_212),
.B2(n_210),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_2909),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3132),
.Y(n_3793)
);

CKINVDCx20_ASAP7_75t_R g3794 ( 
.A(n_2788),
.Y(n_3794)
);

INVx2_ASAP7_75t_L g3795 ( 
.A(n_2933),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3134),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_2943),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3148),
.Y(n_3798)
);

BUFx4f_ASAP7_75t_L g3799 ( 
.A(n_3044),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3157),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3164),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3168),
.Y(n_3802)
);

NAND3xp33_ASAP7_75t_L g3803 ( 
.A(n_3380),
.B(n_213),
.C(n_212),
.Y(n_3803)
);

AO22x2_ASAP7_75t_L g3804 ( 
.A1(n_3075),
.A2(n_214),
.B1(n_215),
.B2(n_213),
.Y(n_3804)
);

AO22x2_ASAP7_75t_L g3805 ( 
.A1(n_3089),
.A2(n_215),
.B1(n_216),
.B2(n_214),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3183),
.Y(n_3806)
);

AO22x2_ASAP7_75t_L g3807 ( 
.A1(n_3092),
.A2(n_215),
.B1(n_216),
.B2(n_214),
.Y(n_3807)
);

INVx2_ASAP7_75t_L g3808 ( 
.A(n_2800),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3170),
.Y(n_3809)
);

NAND3xp33_ASAP7_75t_SL g3810 ( 
.A(n_2758),
.B(n_3),
.C(n_4),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3180),
.Y(n_3811)
);

AO22x2_ASAP7_75t_L g3812 ( 
.A1(n_3063),
.A2(n_218),
.B1(n_219),
.B2(n_217),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3222),
.B(n_217),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3185),
.Y(n_3814)
);

AND2x4_ASAP7_75t_L g3815 ( 
.A(n_2974),
.B(n_217),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3230),
.B(n_218),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_2800),
.Y(n_3817)
);

AOI22xp5_ASAP7_75t_L g3818 ( 
.A1(n_2910),
.A2(n_219),
.B1(n_220),
.B2(n_218),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_2831),
.Y(n_3819)
);

BUFx2_ASAP7_75t_L g3820 ( 
.A(n_3096),
.Y(n_3820)
);

INVx3_ASAP7_75t_L g3821 ( 
.A(n_3174),
.Y(n_3821)
);

AOI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_2911),
.A2(n_220),
.B1(n_221),
.B2(n_219),
.Y(n_3822)
);

BUFx3_ASAP7_75t_L g3823 ( 
.A(n_3093),
.Y(n_3823)
);

BUFx2_ASAP7_75t_L g3824 ( 
.A(n_3086),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_2833),
.Y(n_3825)
);

AND2x4_ASAP7_75t_L g3826 ( 
.A(n_2773),
.B(n_220),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3239),
.B(n_221),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3248),
.B(n_3257),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3109),
.Y(n_3829)
);

NOR2xp33_ASAP7_75t_L g3830 ( 
.A(n_3054),
.B(n_221),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_SL g3831 ( 
.A(n_2990),
.B(n_222),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_2797),
.Y(n_3832)
);

AOI22xp33_ASAP7_75t_L g3833 ( 
.A1(n_2982),
.A2(n_223),
.B1(n_224),
.B2(n_222),
.Y(n_3833)
);

AOI22xp5_ASAP7_75t_L g3834 ( 
.A1(n_2863),
.A2(n_224),
.B1(n_225),
.B2(n_223),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3197),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3037),
.B(n_223),
.Y(n_3836)
);

AO22x2_ASAP7_75t_L g3837 ( 
.A1(n_3166),
.A2(n_225),
.B1(n_226),
.B2(n_224),
.Y(n_3837)
);

AO22x2_ASAP7_75t_L g3838 ( 
.A1(n_3166),
.A2(n_228),
.B1(n_229),
.B2(n_227),
.Y(n_3838)
);

CKINVDCx5p33_ASAP7_75t_R g3839 ( 
.A(n_2855),
.Y(n_3839)
);

OR2x2_ASAP7_75t_SL g3840 ( 
.A(n_2978),
.B(n_227),
.Y(n_3840)
);

OAI22xp5_ASAP7_75t_SL g3841 ( 
.A1(n_3031),
.A2(n_228),
.B1(n_229),
.B2(n_227),
.Y(n_3841)
);

BUFx2_ASAP7_75t_L g3842 ( 
.A(n_3061),
.Y(n_3842)
);

AO22x2_ASAP7_75t_L g3843 ( 
.A1(n_3172),
.A2(n_229),
.B1(n_230),
.B2(n_228),
.Y(n_3843)
);

AO22x2_ASAP7_75t_L g3844 ( 
.A1(n_3172),
.A2(n_3356),
.B1(n_3357),
.B2(n_3349),
.Y(n_3844)
);

CKINVDCx20_ASAP7_75t_R g3845 ( 
.A(n_2782),
.Y(n_3845)
);

AO22x2_ASAP7_75t_L g3846 ( 
.A1(n_3365),
.A2(n_231),
.B1(n_232),
.B2(n_230),
.Y(n_3846)
);

AO22x2_ASAP7_75t_L g3847 ( 
.A1(n_3091),
.A2(n_232),
.B1(n_233),
.B2(n_230),
.Y(n_3847)
);

NOR2xp33_ASAP7_75t_L g3848 ( 
.A(n_2948),
.B(n_233),
.Y(n_3848)
);

AO22x2_ASAP7_75t_L g3849 ( 
.A1(n_3137),
.A2(n_3140),
.B1(n_3152),
.B2(n_3145),
.Y(n_3849)
);

NAND2x1p5_ASAP7_75t_L g3850 ( 
.A(n_2750),
.B(n_233),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3049),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_2975),
.Y(n_3852)
);

AO22x2_ASAP7_75t_L g3853 ( 
.A1(n_3137),
.A2(n_235),
.B1(n_236),
.B2(n_234),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3087),
.Y(n_3854)
);

AO22x2_ASAP7_75t_L g3855 ( 
.A1(n_3140),
.A2(n_235),
.B1(n_236),
.B2(n_234),
.Y(n_3855)
);

AO22x2_ASAP7_75t_L g3856 ( 
.A1(n_3145),
.A2(n_237),
.B1(n_238),
.B2(n_234),
.Y(n_3856)
);

INVxp67_ASAP7_75t_L g3857 ( 
.A(n_3056),
.Y(n_3857)
);

CKINVDCx5p33_ASAP7_75t_R g3858 ( 
.A(n_3064),
.Y(n_3858)
);

INVx3_ASAP7_75t_L g3859 ( 
.A(n_3061),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3088),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_3050),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_2794),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3022),
.B(n_2810),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3039),
.Y(n_3864)
);

BUFx3_ASAP7_75t_L g3865 ( 
.A(n_3112),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3041),
.Y(n_3866)
);

AND2x4_ASAP7_75t_L g3867 ( 
.A(n_2757),
.B(n_237),
.Y(n_3867)
);

NAND2x1p5_ASAP7_75t_L g3868 ( 
.A(n_2750),
.B(n_237),
.Y(n_3868)
);

NAND2x1p5_ASAP7_75t_L g3869 ( 
.A(n_2894),
.B(n_238),
.Y(n_3869)
);

A2O1A1Ixp33_ASAP7_75t_L g3870 ( 
.A1(n_3062),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_3870)
);

NAND2xp33_ASAP7_75t_L g3871 ( 
.A(n_2990),
.B(n_239),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3077),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3085),
.Y(n_3873)
);

AO22x2_ASAP7_75t_L g3874 ( 
.A1(n_3152),
.A2(n_240),
.B1(n_241),
.B2(n_239),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3095),
.Y(n_3875)
);

AO22x2_ASAP7_75t_L g3876 ( 
.A1(n_2920),
.A2(n_241),
.B1(n_242),
.B2(n_240),
.Y(n_3876)
);

BUFx8_ASAP7_75t_L g3877 ( 
.A(n_2990),
.Y(n_3877)
);

NAND2x1p5_ASAP7_75t_L g3878 ( 
.A(n_2894),
.B(n_240),
.Y(n_3878)
);

INVxp67_ASAP7_75t_L g3879 ( 
.A(n_2893),
.Y(n_3879)
);

AND2x4_ASAP7_75t_L g3880 ( 
.A(n_2771),
.B(n_242),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_2850),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_2872),
.Y(n_3882)
);

AND2x4_ASAP7_75t_L g3883 ( 
.A(n_3038),
.B(n_242),
.Y(n_3883)
);

AO22x2_ASAP7_75t_L g3884 ( 
.A1(n_2820),
.A2(n_244),
.B1(n_245),
.B2(n_243),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3101),
.Y(n_3885)
);

INVx3_ASAP7_75t_L g3886 ( 
.A(n_3118),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_2881),
.Y(n_3887)
);

CKINVDCx20_ASAP7_75t_R g3888 ( 
.A(n_2995),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_2885),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3261),
.B(n_243),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3104),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3105),
.Y(n_3892)
);

BUFx2_ASAP7_75t_L g3893 ( 
.A(n_3118),
.Y(n_3893)
);

BUFx3_ASAP7_75t_L g3894 ( 
.A(n_2894),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3107),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3110),
.Y(n_3896)
);

AO22x2_ASAP7_75t_L g3897 ( 
.A1(n_2838),
.A2(n_245),
.B1(n_246),
.B2(n_244),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3115),
.Y(n_3898)
);

OAI221xp5_ASAP7_75t_L g3899 ( 
.A1(n_3272),
.A2(n_246),
.B1(n_247),
.B2(n_245),
.C(n_244),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3350),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3276),
.B(n_3278),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3280),
.B(n_247),
.Y(n_3902)
);

NAND2x1p5_ASAP7_75t_L g3903 ( 
.A(n_2908),
.B(n_248),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_3117),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3352),
.Y(n_3905)
);

AO22x2_ASAP7_75t_L g3906 ( 
.A1(n_2841),
.A2(n_249),
.B1(n_250),
.B2(n_248),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3359),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3133),
.Y(n_3908)
);

BUFx6f_ASAP7_75t_L g3909 ( 
.A(n_2908),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3360),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3368),
.Y(n_3911)
);

HB1xp67_ASAP7_75t_L g3912 ( 
.A(n_3210),
.Y(n_3912)
);

AO22x2_ASAP7_75t_L g3913 ( 
.A1(n_2845),
.A2(n_250),
.B1(n_251),
.B2(n_249),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3191),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3281),
.Y(n_3915)
);

AO22x2_ASAP7_75t_L g3916 ( 
.A1(n_2846),
.A2(n_250),
.B1(n_251),
.B2(n_249),
.Y(n_3916)
);

AOI22xp5_ASAP7_75t_L g3917 ( 
.A1(n_2988),
.A2(n_253),
.B1(n_254),
.B2(n_252),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3282),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_L g3919 ( 
.A(n_2869),
.B(n_252),
.Y(n_3919)
);

CKINVDCx20_ASAP7_75t_R g3920 ( 
.A(n_2997),
.Y(n_3920)
);

AO22x2_ASAP7_75t_L g3921 ( 
.A1(n_2803),
.A2(n_253),
.B1(n_254),
.B2(n_252),
.Y(n_3921)
);

NAND2x1p5_ASAP7_75t_L g3922 ( 
.A(n_2908),
.B(n_2925),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_2991),
.B(n_253),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3283),
.B(n_256),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_3009),
.B(n_256),
.Y(n_3925)
);

INVxp67_ASAP7_75t_L g3926 ( 
.A(n_3218),
.Y(n_3926)
);

BUFx2_ASAP7_75t_L g3927 ( 
.A(n_3100),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3286),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3288),
.B(n_256),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3290),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3156),
.Y(n_3931)
);

AOI22xp5_ASAP7_75t_L g3932 ( 
.A1(n_3128),
.A2(n_258),
.B1(n_259),
.B2(n_257),
.Y(n_3932)
);

INVx3_ASAP7_75t_L g3933 ( 
.A(n_2990),
.Y(n_3933)
);

INVx2_ASAP7_75t_SL g3934 ( 
.A(n_3040),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3175),
.B(n_257),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3156),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3161),
.Y(n_3937)
);

AND2x4_ASAP7_75t_L g3938 ( 
.A(n_3007),
.B(n_257),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3161),
.Y(n_3939)
);

INVxp67_ASAP7_75t_L g3940 ( 
.A(n_3246),
.Y(n_3940)
);

AND2x6_ASAP7_75t_L g3941 ( 
.A(n_2925),
.B(n_258),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3144),
.Y(n_3942)
);

AOI22xp5_ASAP7_75t_L g3943 ( 
.A1(n_2888),
.A2(n_260),
.B1(n_261),
.B2(n_259),
.Y(n_3943)
);

AO22x2_ASAP7_75t_L g3944 ( 
.A1(n_3144),
.A2(n_260),
.B1(n_261),
.B2(n_259),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3351),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3390),
.Y(n_3946)
);

AO22x2_ASAP7_75t_L g3947 ( 
.A1(n_3235),
.A2(n_263),
.B1(n_264),
.B2(n_262),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3010),
.B(n_262),
.Y(n_3948)
);

NAND2x1p5_ASAP7_75t_L g3949 ( 
.A(n_2925),
.B(n_262),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_2919),
.B(n_263),
.Y(n_3950)
);

OAI221xp5_ASAP7_75t_L g3951 ( 
.A1(n_2923),
.A2(n_265),
.B1(n_266),
.B2(n_264),
.C(n_263),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3111),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3131),
.Y(n_3953)
);

AO22x2_ASAP7_75t_L g3954 ( 
.A1(n_3370),
.A2(n_266),
.B1(n_267),
.B2(n_265),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3745),
.A2(n_2857),
.B(n_3285),
.Y(n_3955)
);

HB1xp67_ASAP7_75t_L g3956 ( 
.A(n_3708),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_L g3957 ( 
.A(n_3915),
.B(n_2973),
.Y(n_3957)
);

INVx2_ASAP7_75t_SL g3958 ( 
.A(n_3441),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_SL g3959 ( 
.A(n_3685),
.B(n_3294),
.Y(n_3959)
);

BUFx8_ASAP7_75t_L g3960 ( 
.A(n_3452),
.Y(n_3960)
);

NOR2xp33_ASAP7_75t_L g3961 ( 
.A(n_3428),
.B(n_2914),
.Y(n_3961)
);

AOI21xp5_ASAP7_75t_L g3962 ( 
.A1(n_3871),
.A2(n_2892),
.B(n_2993),
.Y(n_3962)
);

NOR2xp67_ASAP7_75t_L g3963 ( 
.A(n_3509),
.B(n_3046),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_3808),
.A2(n_3005),
.B(n_2993),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_SL g3965 ( 
.A(n_3392),
.B(n_3251),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3918),
.B(n_2932),
.Y(n_3966)
);

BUFx2_ASAP7_75t_L g3967 ( 
.A(n_3653),
.Y(n_3967)
);

O2A1O1Ixp33_ASAP7_75t_L g3968 ( 
.A1(n_3432),
.A2(n_2960),
.B(n_2904),
.C(n_2901),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3928),
.B(n_2891),
.Y(n_3969)
);

AOI22xp5_ASAP7_75t_L g3970 ( 
.A1(n_3457),
.A2(n_3689),
.B1(n_3682),
.B2(n_3540),
.Y(n_3970)
);

AOI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_3817),
.A2(n_3005),
.B(n_2993),
.Y(n_3971)
);

INVx4_ASAP7_75t_L g3972 ( 
.A(n_3941),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3646),
.A2(n_3047),
.B(n_3005),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3646),
.A2(n_3735),
.B(n_3732),
.Y(n_3974)
);

AOI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3738),
.A2(n_3750),
.B(n_3740),
.Y(n_3975)
);

AOI22x1_ASAP7_75t_L g3976 ( 
.A1(n_3406),
.A2(n_3167),
.B1(n_3171),
.B2(n_3147),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_SL g3977 ( 
.A(n_3397),
.B(n_3251),
.Y(n_3977)
);

AOI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_3755),
.A2(n_3073),
.B(n_3047),
.Y(n_3978)
);

INVx2_ASAP7_75t_SL g3979 ( 
.A(n_3596),
.Y(n_3979)
);

A2O1A1Ixp33_ASAP7_75t_L g3980 ( 
.A1(n_3395),
.A2(n_3292),
.B(n_3316),
.C(n_3302),
.Y(n_3980)
);

NOR3xp33_ASAP7_75t_L g3981 ( 
.A(n_3405),
.B(n_2878),
.C(n_2877),
.Y(n_3981)
);

AOI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3758),
.A2(n_3073),
.B(n_3047),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3761),
.A2(n_3195),
.B(n_3073),
.Y(n_3983)
);

AOI21xp5_ASAP7_75t_L g3984 ( 
.A1(n_3640),
.A2(n_3202),
.B(n_3195),
.Y(n_3984)
);

NOR3xp33_ASAP7_75t_L g3985 ( 
.A(n_3686),
.B(n_3024),
.C(n_2934),
.Y(n_3985)
);

HB1xp67_ASAP7_75t_L g3986 ( 
.A(n_3647),
.Y(n_3986)
);

AOI21xp5_ASAP7_75t_L g3987 ( 
.A1(n_3640),
.A2(n_3202),
.B(n_3195),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3930),
.B(n_2976),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3391),
.Y(n_3989)
);

INVx2_ASAP7_75t_L g3990 ( 
.A(n_3401),
.Y(n_3990)
);

O2A1O1Ixp33_ASAP7_75t_L g3991 ( 
.A1(n_3828),
.A2(n_3015),
.B(n_3042),
.C(n_3051),
.Y(n_3991)
);

BUFx2_ASAP7_75t_L g3992 ( 
.A(n_3511),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3400),
.B(n_3126),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3431),
.Y(n_3994)
);

BUFx6f_ASAP7_75t_L g3995 ( 
.A(n_3909),
.Y(n_3995)
);

AOI21xp5_ASAP7_75t_L g3996 ( 
.A1(n_3849),
.A2(n_3241),
.B(n_3202),
.Y(n_3996)
);

OAI21xp5_ASAP7_75t_L g3997 ( 
.A1(n_3901),
.A2(n_3550),
.B(n_3519),
.Y(n_3997)
);

OR2x2_ASAP7_75t_L g3998 ( 
.A(n_3590),
.B(n_3617),
.Y(n_3998)
);

AOI21x1_ASAP7_75t_L g3999 ( 
.A1(n_3748),
.A2(n_3849),
.B(n_3947),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_3639),
.B(n_3053),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_L g4001 ( 
.A(n_3863),
.B(n_3862),
.Y(n_4001)
);

BUFx6f_ASAP7_75t_L g4002 ( 
.A(n_3909),
.Y(n_4002)
);

BUFx2_ASAP7_75t_L g4003 ( 
.A(n_3594),
.Y(n_4003)
);

O2A1O1Ixp33_ASAP7_75t_L g4004 ( 
.A1(n_3420),
.A2(n_3323),
.B(n_3333),
.C(n_3322),
.Y(n_4004)
);

INVx1_ASAP7_75t_SL g4005 ( 
.A(n_3396),
.Y(n_4005)
);

INVx3_ASAP7_75t_L g4006 ( 
.A(n_3670),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3691),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3528),
.B(n_265),
.Y(n_4008)
);

AOI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3699),
.A2(n_3241),
.B(n_3149),
.Y(n_4009)
);

AOI21xp5_ASAP7_75t_L g4010 ( 
.A1(n_3700),
.A2(n_3241),
.B(n_3149),
.Y(n_4010)
);

A2O1A1Ixp33_ASAP7_75t_L g4011 ( 
.A1(n_3943),
.A2(n_3337),
.B(n_3338),
.C(n_3334),
.Y(n_4011)
);

AOI21xp5_ASAP7_75t_L g4012 ( 
.A1(n_3701),
.A2(n_3097),
.B(n_3294),
.Y(n_4012)
);

NOR2xp33_ASAP7_75t_L g4013 ( 
.A(n_3756),
.B(n_3103),
.Y(n_4013)
);

INVx5_ASAP7_75t_L g4014 ( 
.A(n_3941),
.Y(n_4014)
);

NOR3xp33_ASAP7_75t_L g4015 ( 
.A(n_3625),
.B(n_3129),
.C(n_3125),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3704),
.A2(n_3142),
.B(n_3028),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_SL g4017 ( 
.A(n_3694),
.B(n_3059),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3393),
.Y(n_4018)
);

AOI21x1_ASAP7_75t_L g4019 ( 
.A1(n_3954),
.A2(n_3300),
.B(n_2994),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3597),
.B(n_267),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_3711),
.A2(n_3142),
.B(n_3028),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3446),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3715),
.A2(n_3369),
.B(n_3300),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3881),
.B(n_3348),
.Y(n_4024)
);

O2A1O1Ixp33_ASAP7_75t_L g4025 ( 
.A1(n_3857),
.A2(n_3193),
.B(n_3226),
.C(n_3198),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_L g4026 ( 
.A(n_3882),
.B(n_3139),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3398),
.Y(n_4027)
);

AOI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_3716),
.A2(n_3369),
.B(n_2994),
.Y(n_4028)
);

NOR2xp33_ASAP7_75t_L g4029 ( 
.A(n_3879),
.B(n_3150),
.Y(n_4029)
);

AOI21xp5_ASAP7_75t_L g4030 ( 
.A1(n_3717),
.A2(n_3190),
.B(n_2854),
.Y(n_4030)
);

BUFx6f_ASAP7_75t_L g4031 ( 
.A(n_3894),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3887),
.B(n_3135),
.Y(n_4032)
);

AOI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3682),
.A2(n_3163),
.B1(n_3242),
.B2(n_3237),
.Y(n_4033)
);

AOI21xp5_ASAP7_75t_L g4034 ( 
.A1(n_3720),
.A2(n_3141),
.B(n_3060),
.Y(n_4034)
);

HB1xp67_ASAP7_75t_L g4035 ( 
.A(n_3464),
.Y(n_4035)
);

AOI21xp5_ASAP7_75t_L g4036 ( 
.A1(n_3731),
.A2(n_3648),
.B(n_3644),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3889),
.B(n_3819),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3458),
.Y(n_4038)
);

AOI21xp5_ASAP7_75t_L g4039 ( 
.A1(n_3832),
.A2(n_3074),
.B(n_3018),
.Y(n_4039)
);

OAI21xp5_ASAP7_75t_L g4040 ( 
.A1(n_3404),
.A2(n_3043),
.B(n_3127),
.Y(n_4040)
);

OAI22xp5_ASAP7_75t_L g4041 ( 
.A1(n_3840),
.A2(n_3043),
.B1(n_3127),
.B2(n_3136),
.Y(n_4041)
);

AOI21xp5_ASAP7_75t_L g4042 ( 
.A1(n_3835),
.A2(n_3189),
.B(n_2796),
.Y(n_4042)
);

AOI21xp5_ASAP7_75t_L g4043 ( 
.A1(n_3852),
.A2(n_3952),
.B(n_3809),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3407),
.Y(n_4044)
);

AOI21xp5_ASAP7_75t_L g4045 ( 
.A1(n_3767),
.A2(n_2780),
.B(n_2785),
.Y(n_4045)
);

AOI21xp5_ASAP7_75t_L g4046 ( 
.A1(n_3776),
.A2(n_3162),
.B(n_3169),
.Y(n_4046)
);

INVx3_ASAP7_75t_L g4047 ( 
.A(n_3877),
.Y(n_4047)
);

NOR2xp33_ASAP7_75t_L g4048 ( 
.A(n_3581),
.B(n_3159),
.Y(n_4048)
);

OAI22xp5_ASAP7_75t_L g4049 ( 
.A1(n_3707),
.A2(n_3162),
.B1(n_3160),
.B2(n_3165),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3825),
.B(n_3245),
.Y(n_4050)
);

NAND2x1p5_ASAP7_75t_L g4051 ( 
.A(n_3410),
.B(n_3099),
.Y(n_4051)
);

AOI21xp5_ASAP7_75t_L g4052 ( 
.A1(n_3656),
.A2(n_3169),
.B(n_3029),
.Y(n_4052)
);

CKINVDCx10_ASAP7_75t_R g4053 ( 
.A(n_3622),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3811),
.B(n_3250),
.Y(n_4054)
);

HB1xp67_ASAP7_75t_L g4055 ( 
.A(n_3399),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_L g4056 ( 
.A(n_3475),
.B(n_3258),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3409),
.Y(n_4057)
);

OAI22xp5_ASAP7_75t_L g4058 ( 
.A1(n_3587),
.A2(n_3187),
.B1(n_3277),
.B2(n_3269),
.Y(n_4058)
);

AOI22xp5_ASAP7_75t_L g4059 ( 
.A1(n_3607),
.A2(n_3303),
.B1(n_3313),
.B2(n_3284),
.Y(n_4059)
);

INVx4_ASAP7_75t_L g4060 ( 
.A(n_3941),
.Y(n_4060)
);

AO22x1_ASAP7_75t_L g4061 ( 
.A1(n_3624),
.A2(n_3155),
.B1(n_3169),
.B2(n_3176),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_SL g4062 ( 
.A(n_3573),
.B(n_3059),
.Y(n_4062)
);

BUFx12f_ASAP7_75t_L g4063 ( 
.A(n_3566),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3814),
.B(n_3320),
.Y(n_4064)
);

INVx11_ASAP7_75t_L g4065 ( 
.A(n_3784),
.Y(n_4065)
);

AOI21x1_ASAP7_75t_L g4066 ( 
.A1(n_3947),
.A2(n_3029),
.B(n_3328),
.Y(n_4066)
);

OAI21xp5_ASAP7_75t_L g4067 ( 
.A1(n_3803),
.A2(n_3342),
.B(n_3178),
.Y(n_4067)
);

BUFx2_ASAP7_75t_L g4068 ( 
.A(n_3592),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3643),
.B(n_3177),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3416),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3654),
.B(n_3179),
.Y(n_4071)
);

OAI22xp5_ASAP7_75t_L g4072 ( 
.A1(n_3587),
.A2(n_3155),
.B1(n_3186),
.B2(n_3182),
.Y(n_4072)
);

NOR2xp33_ASAP7_75t_L g4073 ( 
.A(n_3591),
.B(n_3702),
.Y(n_4073)
);

AOI21xp5_ASAP7_75t_L g4074 ( 
.A1(n_3677),
.A2(n_3121),
.B(n_3176),
.Y(n_4074)
);

AND2x2_ASAP7_75t_L g4075 ( 
.A(n_3626),
.B(n_267),
.Y(n_4075)
);

AOI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_3696),
.A2(n_3121),
.B(n_3068),
.Y(n_4076)
);

OAI21xp5_ASAP7_75t_L g4077 ( 
.A1(n_3741),
.A2(n_2887),
.B(n_2827),
.Y(n_4077)
);

OAI22xp5_ASAP7_75t_L g4078 ( 
.A1(n_3605),
.A2(n_3121),
.B1(n_2887),
.B2(n_2924),
.Y(n_4078)
);

OAI22xp5_ASAP7_75t_L g4079 ( 
.A1(n_3659),
.A2(n_2887),
.B1(n_2924),
.B2(n_2827),
.Y(n_4079)
);

AOI21xp5_ASAP7_75t_L g4080 ( 
.A1(n_3726),
.A2(n_3068),
.B(n_3059),
.Y(n_4080)
);

AOI21xp5_ASAP7_75t_L g4081 ( 
.A1(n_3753),
.A2(n_3068),
.B(n_3059),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3772),
.B(n_268),
.Y(n_4082)
);

NOR2xp33_ASAP7_75t_L g4083 ( 
.A(n_3749),
.B(n_268),
.Y(n_4083)
);

AOI21xp5_ASAP7_75t_L g4084 ( 
.A1(n_3765),
.A2(n_3068),
.B(n_3059),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3931),
.B(n_268),
.Y(n_4085)
);

BUFx2_ASAP7_75t_L g4086 ( 
.A(n_3615),
.Y(n_4086)
);

AOI21xp5_ASAP7_75t_L g4087 ( 
.A1(n_3769),
.A2(n_3068),
.B(n_2887),
.Y(n_4087)
);

INVxp67_ASAP7_75t_L g4088 ( 
.A(n_3659),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_SL g4089 ( 
.A(n_3415),
.B(n_2962),
.Y(n_4089)
);

O2A1O1Ixp33_ASAP7_75t_L g4090 ( 
.A1(n_3935),
.A2(n_270),
.B(n_271),
.C(n_269),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3423),
.Y(n_4091)
);

AOI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_3770),
.A2(n_2887),
.B(n_2827),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3936),
.B(n_3937),
.Y(n_4093)
);

INVxp67_ASAP7_75t_L g4094 ( 
.A(n_3662),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3429),
.Y(n_4095)
);

O2A1O1Ixp33_ASAP7_75t_L g4096 ( 
.A1(n_3676),
.A2(n_270),
.B(n_271),
.C(n_269),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3939),
.B(n_269),
.Y(n_4097)
);

A2O1A1Ixp33_ASAP7_75t_L g4098 ( 
.A1(n_3660),
.A2(n_2924),
.B(n_2962),
.C(n_2827),
.Y(n_4098)
);

NOR2xp33_ASAP7_75t_L g4099 ( 
.A(n_3858),
.B(n_270),
.Y(n_4099)
);

INVx2_ASAP7_75t_L g4100 ( 
.A(n_3462),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_3942),
.B(n_271),
.Y(n_4101)
);

NAND2x1p5_ASAP7_75t_L g4102 ( 
.A(n_3414),
.B(n_2827),
.Y(n_4102)
);

INVx4_ASAP7_75t_L g4103 ( 
.A(n_3496),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3864),
.B(n_3866),
.Y(n_4104)
);

AOI21xp5_ASAP7_75t_L g4105 ( 
.A1(n_3777),
.A2(n_2962),
.B(n_2924),
.Y(n_4105)
);

NAND2x1p5_ASAP7_75t_L g4106 ( 
.A(n_3412),
.B(n_2924),
.Y(n_4106)
);

AOI21xp5_ASAP7_75t_L g4107 ( 
.A1(n_3444),
.A2(n_2962),
.B(n_273),
.Y(n_4107)
);

OAI21x1_ASAP7_75t_L g4108 ( 
.A1(n_3933),
.A2(n_2962),
.B(n_273),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3430),
.B(n_3435),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_3436),
.B(n_272),
.Y(n_4110)
);

AO21x1_ASAP7_75t_L g4111 ( 
.A1(n_3570),
.A2(n_273),
.B(n_272),
.Y(n_4111)
);

AOI21xp5_ASAP7_75t_L g4112 ( 
.A1(n_3664),
.A2(n_274),
.B(n_272),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3438),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3442),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3443),
.B(n_274),
.Y(n_4115)
);

NOR2xp67_ASAP7_75t_L g4116 ( 
.A(n_3440),
.B(n_3561),
.Y(n_4116)
);

OAI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_3723),
.A2(n_275),
.B1(n_276),
.B2(n_274),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3448),
.B(n_275),
.Y(n_4118)
);

AOI21xp5_ASAP7_75t_L g4119 ( 
.A1(n_3668),
.A2(n_276),
.B(n_275),
.Y(n_4119)
);

AOI21xp5_ASAP7_75t_L g4120 ( 
.A1(n_3844),
.A2(n_3469),
.B(n_3831),
.Y(n_4120)
);

BUFx6f_ASAP7_75t_L g4121 ( 
.A(n_3922),
.Y(n_4121)
);

A2O1A1Ixp33_ASAP7_75t_L g4122 ( 
.A1(n_3752),
.A2(n_278),
.B(n_279),
.C(n_277),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_SL g4123 ( 
.A(n_3417),
.B(n_277),
.Y(n_4123)
);

INVxp67_ASAP7_75t_L g4124 ( 
.A(n_3499),
.Y(n_4124)
);

CKINVDCx10_ASAP7_75t_R g4125 ( 
.A(n_3564),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_3455),
.B(n_278),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3488),
.B(n_1070),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_L g4128 ( 
.A1(n_3723),
.A2(n_279),
.B1(n_280),
.B2(n_278),
.Y(n_4128)
);

NOR2xp67_ASAP7_75t_L g4129 ( 
.A(n_3447),
.B(n_279),
.Y(n_4129)
);

OAI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_3757),
.A2(n_281),
.B(n_280),
.Y(n_4130)
);

AOI21xp5_ASAP7_75t_L g4131 ( 
.A1(n_3844),
.A2(n_281),
.B(n_280),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_3459),
.B(n_282),
.Y(n_4132)
);

O2A1O1Ixp33_ASAP7_75t_SL g4133 ( 
.A1(n_3810),
.A2(n_1059),
.B(n_1060),
.C(n_1058),
.Y(n_4133)
);

AND2x4_ASAP7_75t_L g4134 ( 
.A(n_3886),
.B(n_282),
.Y(n_4134)
);

AOI21xp5_ASAP7_75t_L g4135 ( 
.A1(n_3742),
.A2(n_3829),
.B(n_3403),
.Y(n_4135)
);

AOI22xp5_ASAP7_75t_L g4136 ( 
.A1(n_3775),
.A2(n_283),
.B1(n_285),
.B2(n_282),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_3461),
.B(n_283),
.Y(n_4137)
);

NAND3xp33_ASAP7_75t_SL g4138 ( 
.A(n_3451),
.B(n_5),
.C(n_6),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3465),
.B(n_285),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_3481),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3468),
.Y(n_4141)
);

AOI21xp5_ASAP7_75t_L g4142 ( 
.A1(n_3742),
.A2(n_287),
.B(n_286),
.Y(n_4142)
);

BUFx6f_ASAP7_75t_L g4143 ( 
.A(n_3427),
.Y(n_4143)
);

AOI22xp5_ASAP7_75t_L g4144 ( 
.A1(n_3794),
.A2(n_287),
.B1(n_288),
.B2(n_286),
.Y(n_4144)
);

BUFx6f_ASAP7_75t_L g4145 ( 
.A(n_3427),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3470),
.Y(n_4146)
);

OAI22xp5_ASAP7_75t_L g4147 ( 
.A1(n_3760),
.A2(n_287),
.B1(n_288),
.B2(n_286),
.Y(n_4147)
);

NAND2x1p5_ASAP7_75t_L g4148 ( 
.A(n_3454),
.B(n_291),
.Y(n_4148)
);

AOI21xp5_ASAP7_75t_L g4149 ( 
.A1(n_3954),
.A2(n_289),
.B(n_288),
.Y(n_4149)
);

AOI21xp5_ASAP7_75t_L g4150 ( 
.A1(n_3900),
.A2(n_290),
.B(n_289),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_3675),
.B(n_290),
.Y(n_4151)
);

AOI21xp5_ASAP7_75t_L g4152 ( 
.A1(n_3905),
.A2(n_291),
.B(n_290),
.Y(n_4152)
);

A2O1A1Ixp33_ASAP7_75t_L g4153 ( 
.A1(n_3421),
.A2(n_293),
.B(n_294),
.C(n_292),
.Y(n_4153)
);

AOI21xp5_ASAP7_75t_L g4154 ( 
.A1(n_3907),
.A2(n_293),
.B(n_292),
.Y(n_4154)
);

INVx3_ASAP7_75t_L g4155 ( 
.A(n_3483),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_3476),
.B(n_292),
.Y(n_4156)
);

INVx3_ASAP7_75t_L g4157 ( 
.A(n_3483),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3478),
.B(n_295),
.Y(n_4158)
);

NOR2xp33_ASAP7_75t_L g4159 ( 
.A(n_3479),
.B(n_295),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_3500),
.Y(n_4160)
);

AOI21xp5_ASAP7_75t_L g4161 ( 
.A1(n_3910),
.A2(n_296),
.B(n_295),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_3501),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3486),
.B(n_296),
.Y(n_4163)
);

NAND2x1_ASAP7_75t_L g4164 ( 
.A(n_3624),
.B(n_297),
.Y(n_4164)
);

INVx1_ASAP7_75t_SL g4165 ( 
.A(n_3482),
.Y(n_4165)
);

AOI21xp5_ASAP7_75t_L g4166 ( 
.A1(n_3911),
.A2(n_3680),
.B(n_3521),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3489),
.Y(n_4167)
);

OAI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_3760),
.A2(n_298),
.B1(n_299),
.B2(n_297),
.Y(n_4168)
);

A2O1A1Ixp33_ASAP7_75t_L g4169 ( 
.A1(n_3932),
.A2(n_298),
.B(n_300),
.C(n_297),
.Y(n_4169)
);

NOR2xp33_ASAP7_75t_L g4170 ( 
.A(n_3480),
.B(n_298),
.Y(n_4170)
);

CKINVDCx5p33_ASAP7_75t_R g4171 ( 
.A(n_3460),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3490),
.Y(n_4172)
);

BUFx6f_ASAP7_75t_L g4173 ( 
.A(n_3823),
.Y(n_4173)
);

AOI21xp5_ASAP7_75t_L g4174 ( 
.A1(n_3507),
.A2(n_301),
.B(n_300),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_3491),
.Y(n_4175)
);

AOI21xp5_ASAP7_75t_L g4176 ( 
.A1(n_3533),
.A2(n_301),
.B(n_300),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_3493),
.B(n_301),
.Y(n_4177)
);

O2A1O1Ixp5_ASAP7_75t_L g4178 ( 
.A1(n_3945),
.A2(n_304),
.B(n_305),
.C(n_303),
.Y(n_4178)
);

AOI21xp5_ASAP7_75t_L g4179 ( 
.A1(n_3535),
.A2(n_305),
.B(n_303),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_3759),
.B(n_1065),
.Y(n_4180)
);

OAI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_3394),
.A2(n_307),
.B1(n_308),
.B2(n_306),
.Y(n_4181)
);

NOR2xp67_ASAP7_75t_L g4182 ( 
.A(n_3520),
.B(n_306),
.Y(n_4182)
);

AOI21xp5_ASAP7_75t_L g4183 ( 
.A1(n_3551),
.A2(n_307),
.B(n_306),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3494),
.B(n_307),
.Y(n_4184)
);

AOI21xp5_ASAP7_75t_L g4185 ( 
.A1(n_3554),
.A2(n_309),
.B(n_308),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_3556),
.A2(n_309),
.B(n_308),
.Y(n_4186)
);

O2A1O1Ixp33_ASAP7_75t_L g4187 ( 
.A1(n_3950),
.A2(n_310),
.B(n_311),
.C(n_309),
.Y(n_4187)
);

O2A1O1Ixp33_ASAP7_75t_L g4188 ( 
.A1(n_3517),
.A2(n_312),
.B(n_313),
.C(n_311),
.Y(n_4188)
);

O2A1O1Ixp33_ASAP7_75t_L g4189 ( 
.A1(n_3552),
.A2(n_312),
.B(n_313),
.C(n_311),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_3502),
.B(n_314),
.Y(n_4190)
);

CKINVDCx20_ASAP7_75t_R g4191 ( 
.A(n_3559),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3503),
.Y(n_4192)
);

AOI21xp5_ASAP7_75t_L g4193 ( 
.A1(n_3612),
.A2(n_315),
.B(n_314),
.Y(n_4193)
);

NOR2xp33_ASAP7_75t_R g4194 ( 
.A(n_3637),
.B(n_315),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_3504),
.B(n_315),
.Y(n_4195)
);

NOR2xp33_ASAP7_75t_L g4196 ( 
.A(n_3927),
.B(n_316),
.Y(n_4196)
);

NOR2xp33_ASAP7_75t_L g4197 ( 
.A(n_3411),
.B(n_316),
.Y(n_4197)
);

AND2x4_ASAP7_75t_L g4198 ( 
.A(n_3893),
.B(n_316),
.Y(n_4198)
);

OAI221xp5_ASAP7_75t_L g4199 ( 
.A1(n_3824),
.A2(n_319),
.B1(n_320),
.B2(n_318),
.C(n_317),
.Y(n_4199)
);

OAI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_3394),
.A2(n_3419),
.B1(n_3557),
.B2(n_3445),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_3516),
.B(n_317),
.Y(n_4201)
);

OR2x2_ASAP7_75t_L g4202 ( 
.A(n_3618),
.B(n_3620),
.Y(n_4202)
);

NAND3xp33_ASAP7_75t_L g4203 ( 
.A(n_3830),
.B(n_1061),
.C(n_1060),
.Y(n_4203)
);

AOI21xp5_ASAP7_75t_L g4204 ( 
.A1(n_3614),
.A2(n_318),
.B(n_317),
.Y(n_4204)
);

O2A1O1Ixp33_ASAP7_75t_L g4205 ( 
.A1(n_3569),
.A2(n_320),
.B(n_321),
.C(n_319),
.Y(n_4205)
);

NAND3xp33_ASAP7_75t_SL g4206 ( 
.A(n_3450),
.B(n_3628),
.C(n_3621),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_3629),
.B(n_1063),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_SL g4208 ( 
.A(n_3546),
.B(n_319),
.Y(n_4208)
);

A2O1A1Ixp33_ASAP7_75t_L g4209 ( 
.A1(n_3870),
.A2(n_322),
.B(n_323),
.C(n_321),
.Y(n_4209)
);

A2O1A1Ixp33_ASAP7_75t_L g4210 ( 
.A1(n_3919),
.A2(n_3848),
.B(n_3951),
.C(n_3751),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_3524),
.B(n_321),
.Y(n_4211)
);

HB1xp67_ASAP7_75t_L g4212 ( 
.A(n_3433),
.Y(n_4212)
);

OAI22xp5_ASAP7_75t_L g4213 ( 
.A1(n_3419),
.A2(n_323),
.B1(n_324),
.B2(n_322),
.Y(n_4213)
);

AOI21x1_ASAP7_75t_L g4214 ( 
.A1(n_3912),
.A2(n_323),
.B(n_322),
.Y(n_4214)
);

NOR2xp33_ASAP7_75t_L g4215 ( 
.A(n_3583),
.B(n_324),
.Y(n_4215)
);

OAI21x1_ASAP7_75t_L g4216 ( 
.A1(n_3522),
.A2(n_327),
.B(n_326),
.Y(n_4216)
);

NOR2x1_ASAP7_75t_R g4217 ( 
.A(n_3471),
.B(n_327),
.Y(n_4217)
);

AOI22xp5_ASAP7_75t_L g4218 ( 
.A1(n_3624),
.A2(n_329),
.B1(n_330),
.B2(n_328),
.Y(n_4218)
);

AOI21xp5_ASAP7_75t_L g4219 ( 
.A1(n_3641),
.A2(n_329),
.B(n_328),
.Y(n_4219)
);

NOR2xp33_ASAP7_75t_L g4220 ( 
.A(n_3709),
.B(n_330),
.Y(n_4220)
);

AOI21xp5_ASAP7_75t_L g4221 ( 
.A1(n_3645),
.A2(n_332),
.B(n_331),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_3529),
.B(n_331),
.Y(n_4222)
);

AOI21xp5_ASAP7_75t_L g4223 ( 
.A1(n_3692),
.A2(n_333),
.B(n_332),
.Y(n_4223)
);

AOI21xp5_ASAP7_75t_L g4224 ( 
.A1(n_3703),
.A2(n_333),
.B(n_332),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3536),
.Y(n_4225)
);

AOI21xp5_ASAP7_75t_L g4226 ( 
.A1(n_3721),
.A2(n_335),
.B(n_334),
.Y(n_4226)
);

AOI21xp5_ASAP7_75t_L g4227 ( 
.A1(n_3728),
.A2(n_335),
.B(n_334),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_3505),
.A2(n_335),
.B(n_334),
.Y(n_4228)
);

AOI21xp5_ASAP7_75t_L g4229 ( 
.A1(n_3525),
.A2(n_337),
.B(n_336),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_3537),
.B(n_336),
.Y(n_4230)
);

AND2x2_ASAP7_75t_L g4231 ( 
.A(n_3627),
.B(n_1063),
.Y(n_4231)
);

AOI21xp5_ASAP7_75t_L g4232 ( 
.A1(n_3567),
.A2(n_338),
.B(n_337),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_3631),
.B(n_1066),
.Y(n_4233)
);

AOI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_3600),
.A2(n_340),
.B(n_339),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_3538),
.B(n_3539),
.Y(n_4235)
);

BUFx3_ASAP7_75t_L g4236 ( 
.A(n_3657),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_3632),
.Y(n_4237)
);

AOI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_3914),
.A2(n_3747),
.B(n_3729),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_3684),
.A2(n_341),
.B(n_339),
.Y(n_4239)
);

OAI22xp5_ASAP7_75t_L g4240 ( 
.A1(n_3437),
.A2(n_343),
.B1(n_344),
.B2(n_342),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_3541),
.B(n_342),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_3841),
.A2(n_343),
.B1(n_344),
.B2(n_342),
.Y(n_4242)
);

AOI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_3690),
.A2(n_344),
.B(n_343),
.Y(n_4243)
);

CKINVDCx8_ASAP7_75t_R g4244 ( 
.A(n_3483),
.Y(n_4244)
);

NOR2xp33_ASAP7_75t_L g4245 ( 
.A(n_3778),
.B(n_345),
.Y(n_4245)
);

BUFx6f_ASAP7_75t_L g4246 ( 
.A(n_3865),
.Y(n_4246)
);

OAI22xp5_ASAP7_75t_L g4247 ( 
.A1(n_3512),
.A2(n_346),
.B1(n_347),
.B2(n_345),
.Y(n_4247)
);

BUFx6f_ASAP7_75t_L g4248 ( 
.A(n_3842),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_3543),
.Y(n_4249)
);

AOI21x1_ASAP7_75t_L g4250 ( 
.A1(n_3812),
.A2(n_346),
.B(n_345),
.Y(n_4250)
);

AOI21xp5_ASAP7_75t_L g4251 ( 
.A1(n_3812),
.A2(n_347),
.B(n_346),
.Y(n_4251)
);

AOI22xp33_ASAP7_75t_L g4252 ( 
.A1(n_3661),
.A2(n_348),
.B1(n_349),
.B2(n_347),
.Y(n_4252)
);

AOI21xp5_ASAP7_75t_L g4253 ( 
.A1(n_3780),
.A2(n_349),
.B(n_348),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_3544),
.B(n_3548),
.Y(n_4254)
);

OAI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_3813),
.A2(n_351),
.B(n_350),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_3633),
.Y(n_4256)
);

OAI22xp5_ASAP7_75t_L g4257 ( 
.A1(n_3508),
.A2(n_3449),
.B1(n_3453),
.B2(n_3439),
.Y(n_4257)
);

AOI21x1_ASAP7_75t_L g4258 ( 
.A1(n_3946),
.A2(n_351),
.B(n_350),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_3553),
.Y(n_4259)
);

NAND2x1p5_ASAP7_75t_L g4260 ( 
.A(n_3484),
.B(n_354),
.Y(n_4260)
);

CKINVDCx10_ASAP7_75t_R g4261 ( 
.A(n_3744),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3555),
.B(n_350),
.Y(n_4262)
);

NOR2xp33_ASAP7_75t_L g4263 ( 
.A(n_3523),
.B(n_352),
.Y(n_4263)
);

NAND3xp33_ASAP7_75t_L g4264 ( 
.A(n_3413),
.B(n_1065),
.C(n_1064),
.Y(n_4264)
);

AND2x4_ASAP7_75t_L g4265 ( 
.A(n_3635),
.B(n_353),
.Y(n_4265)
);

OAI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_3816),
.A2(n_354),
.B(n_353),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_3558),
.Y(n_4267)
);

INVx8_ASAP7_75t_L g4268 ( 
.A(n_3514),
.Y(n_4268)
);

OAI22xp5_ASAP7_75t_L g4269 ( 
.A1(n_3439),
.A2(n_354),
.B1(n_355),
.B2(n_353),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_3560),
.B(n_355),
.Y(n_4270)
);

AOI21xp5_ASAP7_75t_L g4271 ( 
.A1(n_3827),
.A2(n_3902),
.B(n_3890),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_3565),
.B(n_355),
.Y(n_4272)
);

OR2x2_ASAP7_75t_L g4273 ( 
.A(n_3636),
.B(n_356),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_3568),
.Y(n_4274)
);

INVx5_ASAP7_75t_L g4275 ( 
.A(n_3821),
.Y(n_4275)
);

AOI21xp5_ASAP7_75t_L g4276 ( 
.A1(n_3924),
.A2(n_357),
.B(n_356),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_L g4277 ( 
.A(n_3598),
.B(n_356),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_3799),
.B(n_358),
.Y(n_4278)
);

AOI21xp5_ASAP7_75t_L g4279 ( 
.A1(n_3929),
.A2(n_3792),
.B(n_3787),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_SL g4280 ( 
.A(n_3712),
.B(n_358),
.Y(n_4280)
);

INVx3_ASAP7_75t_L g4281 ( 
.A(n_3714),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_3602),
.Y(n_4282)
);

AOI21xp5_ASAP7_75t_L g4283 ( 
.A1(n_3795),
.A2(n_359),
.B(n_358),
.Y(n_4283)
);

AOI21xp5_ASAP7_75t_L g4284 ( 
.A1(n_3797),
.A2(n_360),
.B(n_359),
.Y(n_4284)
);

INVx2_ASAP7_75t_SL g4285 ( 
.A(n_3638),
.Y(n_4285)
);

AOI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_3851),
.A2(n_360),
.B(n_359),
.Y(n_4286)
);

AOI21xp5_ASAP7_75t_L g4287 ( 
.A1(n_3861),
.A2(n_361),
.B(n_360),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_3872),
.A2(n_362),
.B(n_361),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_3608),
.B(n_362),
.Y(n_4289)
);

BUFx6f_ASAP7_75t_L g4290 ( 
.A(n_3725),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_3609),
.Y(n_4291)
);

OAI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_3948),
.A2(n_364),
.B(n_363),
.Y(n_4292)
);

O2A1O1Ixp33_ASAP7_75t_L g4293 ( 
.A1(n_3588),
.A2(n_364),
.B(n_365),
.C(n_363),
.Y(n_4293)
);

HB1xp67_ASAP7_75t_L g4294 ( 
.A(n_3762),
.Y(n_4294)
);

A2O1A1Ixp33_ASAP7_75t_L g4295 ( 
.A1(n_3630),
.A2(n_3754),
.B(n_3899),
.C(n_3743),
.Y(n_4295)
);

NOR2xp67_ASAP7_75t_L g4296 ( 
.A(n_3688),
.B(n_364),
.Y(n_4296)
);

OAI22xp5_ASAP7_75t_L g4297 ( 
.A1(n_3449),
.A2(n_366),
.B1(n_367),
.B2(n_365),
.Y(n_4297)
);

AND2x4_ASAP7_75t_L g4298 ( 
.A(n_3610),
.B(n_3611),
.Y(n_4298)
);

OAI21xp5_ASAP7_75t_L g4299 ( 
.A1(n_3408),
.A2(n_366),
.B(n_365),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_SL g4300 ( 
.A(n_3779),
.B(n_366),
.Y(n_4300)
);

NOR2xp33_ASAP7_75t_SL g4301 ( 
.A(n_3888),
.B(n_367),
.Y(n_4301)
);

OAI21xp5_ASAP7_75t_L g4302 ( 
.A1(n_3623),
.A2(n_368),
.B(n_367),
.Y(n_4302)
);

INVx2_ASAP7_75t_SL g4303 ( 
.A(n_3527),
.Y(n_4303)
);

INVx3_ASAP7_75t_L g4304 ( 
.A(n_3698),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_3572),
.Y(n_4305)
);

OAI21xp5_ASAP7_75t_L g4306 ( 
.A1(n_3687),
.A2(n_3658),
.B(n_3665),
.Y(n_4306)
);

HB1xp67_ASAP7_75t_L g4307 ( 
.A(n_3764),
.Y(n_4307)
);

OAI22xp5_ASAP7_75t_L g4308 ( 
.A1(n_3453),
.A2(n_369),
.B1(n_370),
.B2(n_368),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_SL g4309 ( 
.A(n_3850),
.B(n_3868),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_3873),
.A2(n_369),
.B(n_368),
.Y(n_4310)
);

AOI21xp5_ASAP7_75t_L g4311 ( 
.A1(n_3875),
.A2(n_371),
.B(n_370),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3575),
.Y(n_4312)
);

OAI21xp5_ASAP7_75t_L g4313 ( 
.A1(n_3402),
.A2(n_3426),
.B(n_3836),
.Y(n_4313)
);

AOI21xp5_ASAP7_75t_L g4314 ( 
.A1(n_3885),
.A2(n_372),
.B(n_370),
.Y(n_4314)
);

BUFx6f_ASAP7_75t_L g4315 ( 
.A(n_3869),
.Y(n_4315)
);

OAI22xp5_ASAP7_75t_L g4316 ( 
.A1(n_3599),
.A2(n_373),
.B1(n_374),
.B2(n_372),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_3891),
.B(n_372),
.Y(n_4317)
);

AND2x2_ASAP7_75t_L g4318 ( 
.A(n_3695),
.B(n_1068),
.Y(n_4318)
);

AOI21xp5_ASAP7_75t_L g4319 ( 
.A1(n_3898),
.A2(n_374),
.B(n_373),
.Y(n_4319)
);

AOI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_3904),
.A2(n_374),
.B(n_373),
.Y(n_4320)
);

AOI21xp5_ASAP7_75t_L g4321 ( 
.A1(n_3908),
.A2(n_376),
.B(n_375),
.Y(n_4321)
);

INVxp67_ASAP7_75t_L g4322 ( 
.A(n_3815),
.Y(n_4322)
);

OAI21x1_ASAP7_75t_L g4323 ( 
.A1(n_3878),
.A2(n_376),
.B(n_375),
.Y(n_4323)
);

HB1xp67_ASAP7_75t_L g4324 ( 
.A(n_3613),
.Y(n_4324)
);

AND2x2_ASAP7_75t_L g4325 ( 
.A(n_3710),
.B(n_3730),
.Y(n_4325)
);

AOI21xp5_ASAP7_75t_L g4326 ( 
.A1(n_3953),
.A2(n_376),
.B(n_375),
.Y(n_4326)
);

A2O1A1Ixp33_ASAP7_75t_L g4327 ( 
.A1(n_3834),
.A2(n_378),
.B(n_379),
.C(n_377),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_3576),
.Y(n_4328)
);

AOI21x1_ASAP7_75t_L g4329 ( 
.A1(n_3771),
.A2(n_378),
.B(n_377),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_3892),
.B(n_379),
.Y(n_4330)
);

INVx3_ASAP7_75t_L g4331 ( 
.A(n_3903),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_3736),
.B(n_1057),
.Y(n_4332)
);

AND2x2_ASAP7_75t_SL g4333 ( 
.A(n_3532),
.B(n_379),
.Y(n_4333)
);

INVx2_ASAP7_75t_SL g4334 ( 
.A(n_3424),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_3895),
.B(n_3896),
.Y(n_4335)
);

NOR2xp33_ASAP7_75t_L g4336 ( 
.A(n_3920),
.B(n_380),
.Y(n_4336)
);

A2O1A1Ixp33_ASAP7_75t_L g4337 ( 
.A1(n_3785),
.A2(n_382),
.B(n_383),
.C(n_381),
.Y(n_4337)
);

OAI21xp33_ASAP7_75t_L g4338 ( 
.A1(n_3706),
.A2(n_6),
.B(n_7),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_3854),
.B(n_381),
.Y(n_4339)
);

OAI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_3923),
.A2(n_383),
.B(n_382),
.Y(n_4340)
);

O2A1O1Ixp33_ASAP7_75t_L g4341 ( 
.A1(n_3601),
.A2(n_383),
.B(n_384),
.C(n_382),
.Y(n_4341)
);

AOI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_3786),
.A2(n_385),
.B(n_384),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_3578),
.Y(n_4343)
);

AOI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_3788),
.A2(n_386),
.B(n_385),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_3860),
.B(n_385),
.Y(n_4345)
);

AND2x6_ASAP7_75t_L g4346 ( 
.A(n_3678),
.B(n_389),
.Y(n_4346)
);

NOR2xp33_ASAP7_75t_L g4347 ( 
.A(n_3845),
.B(n_386),
.Y(n_4347)
);

O2A1O1Ixp33_ASAP7_75t_L g4348 ( 
.A1(n_3606),
.A2(n_388),
.B(n_389),
.C(n_387),
.Y(n_4348)
);

AOI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_3789),
.A2(n_3796),
.B(n_3793),
.Y(n_4349)
);

AO21x1_ASAP7_75t_L g4350 ( 
.A1(n_3949),
.A2(n_388),
.B(n_387),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_3763),
.B(n_388),
.Y(n_4351)
);

AOI21x1_ASAP7_75t_L g4352 ( 
.A1(n_3434),
.A2(n_390),
.B(n_389),
.Y(n_4352)
);

NOR2xp33_ASAP7_75t_L g4353 ( 
.A(n_3697),
.B(n_390),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_3474),
.A2(n_391),
.B1(n_392),
.B2(n_390),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_SL g4355 ( 
.A(n_3666),
.B(n_391),
.Y(n_4355)
);

AOI22x1_ASAP7_75t_L g4356 ( 
.A1(n_3706),
.A2(n_392),
.B1(n_393),
.B2(n_391),
.Y(n_4356)
);

NOR2xp33_ASAP7_75t_L g4357 ( 
.A(n_3839),
.B(n_392),
.Y(n_4357)
);

AOI21xp5_ASAP7_75t_L g4358 ( 
.A1(n_3798),
.A2(n_3801),
.B(n_3800),
.Y(n_4358)
);

AND2x2_ASAP7_75t_SL g4359 ( 
.A(n_3542),
.B(n_393),
.Y(n_4359)
);

AOI21xp5_ASAP7_75t_L g4360 ( 
.A1(n_3802),
.A2(n_394),
.B(n_393),
.Y(n_4360)
);

NOR2xp33_ASAP7_75t_SL g4361 ( 
.A(n_3669),
.B(n_394),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_3579),
.Y(n_4362)
);

AOI21xp5_ASAP7_75t_L g4363 ( 
.A1(n_3806),
.A2(n_396),
.B(n_394),
.Y(n_4363)
);

INVx4_ASAP7_75t_L g4364 ( 
.A(n_3485),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_3766),
.B(n_396),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_3650),
.B(n_396),
.Y(n_4366)
);

INVx2_ASAP7_75t_SL g4367 ( 
.A(n_3790),
.Y(n_4367)
);

NAND2xp5_ASAP7_75t_L g4368 ( 
.A(n_3655),
.B(n_3667),
.Y(n_4368)
);

AND2x4_ASAP7_75t_L g4369 ( 
.A(n_3580),
.B(n_397),
.Y(n_4369)
);

NOR2xp33_ASAP7_75t_L g4370 ( 
.A(n_3705),
.B(n_3577),
.Y(n_4370)
);

OAI21xp5_ASAP7_75t_L g4371 ( 
.A1(n_3925),
.A2(n_3425),
.B(n_3418),
.Y(n_4371)
);

CKINVDCx10_ASAP7_75t_R g4372 ( 
.A(n_3783),
.Y(n_4372)
);

NOR2xp33_ASAP7_75t_L g4373 ( 
.A(n_3672),
.B(n_3820),
.Y(n_4373)
);

AOI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_3584),
.A2(n_398),
.B(n_397),
.Y(n_4374)
);

AND2x2_ASAP7_75t_SL g4375 ( 
.A(n_3545),
.B(n_399),
.Y(n_4375)
);

NOR2x1p5_ASAP7_75t_SL g4376 ( 
.A(n_3673),
.B(n_3674),
.Y(n_4376)
);

AOI21xp5_ASAP7_75t_L g4377 ( 
.A1(n_3585),
.A2(n_3683),
.B(n_3589),
.Y(n_4377)
);

O2A1O1Ixp33_ASAP7_75t_L g4378 ( 
.A1(n_3467),
.A2(n_3473),
.B(n_3940),
.C(n_3926),
.Y(n_4378)
);

NOR2xp67_ASAP7_75t_L g4379 ( 
.A(n_3934),
.B(n_399),
.Y(n_4379)
);

AOI21xp5_ASAP7_75t_L g4380 ( 
.A1(n_3837),
.A2(n_401),
.B(n_400),
.Y(n_4380)
);

OAI21xp5_ASAP7_75t_L g4381 ( 
.A1(n_3463),
.A2(n_401),
.B(n_400),
.Y(n_4381)
);

OAI21xp33_ASAP7_75t_L g4382 ( 
.A1(n_3718),
.A2(n_6),
.B(n_7),
.Y(n_4382)
);

INVx4_ASAP7_75t_L g4383 ( 
.A(n_3422),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_3595),
.B(n_401),
.Y(n_4384)
);

AOI22xp5_ASAP7_75t_L g4385 ( 
.A1(n_3739),
.A2(n_403),
.B1(n_404),
.B2(n_402),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_3434),
.Y(n_4386)
);

OAI221xp5_ASAP7_75t_L g4387 ( 
.A1(n_3681),
.A2(n_405),
.B1(n_406),
.B2(n_403),
.C(n_402),
.Y(n_4387)
);

INVxp67_ASAP7_75t_L g4388 ( 
.A(n_3547),
.Y(n_4388)
);

BUFx8_ASAP7_75t_L g4389 ( 
.A(n_3649),
.Y(n_4389)
);

OAI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_3818),
.A2(n_405),
.B(n_402),
.Y(n_4390)
);

AOI22xp5_ASAP7_75t_L g4391 ( 
.A1(n_3867),
.A2(n_406),
.B1(n_407),
.B2(n_405),
.Y(n_4391)
);

A2O1A1Ixp33_ASAP7_75t_L g4392 ( 
.A1(n_3822),
.A2(n_408),
.B(n_409),
.C(n_407),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_3944),
.Y(n_4393)
);

NOR2xp33_ASAP7_75t_L g4394 ( 
.A(n_3619),
.B(n_408),
.Y(n_4394)
);

OAI21xp5_ASAP7_75t_L g4395 ( 
.A1(n_3917),
.A2(n_410),
.B(n_409),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_3603),
.B(n_409),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_3466),
.Y(n_4397)
);

AOI22xp5_ASAP7_75t_L g4398 ( 
.A1(n_3880),
.A2(n_411),
.B1(n_412),
.B2(n_410),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_3679),
.B(n_410),
.Y(n_4399)
);

AOI21xp5_ASAP7_75t_L g4400 ( 
.A1(n_3837),
.A2(n_413),
.B(n_411),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_3713),
.B(n_411),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_SL g4402 ( 
.A(n_3562),
.B(n_3571),
.Y(n_4402)
);

AOI21xp5_ASAP7_75t_L g4403 ( 
.A1(n_3838),
.A2(n_414),
.B(n_413),
.Y(n_4403)
);

OAI321xp33_ASAP7_75t_L g4404 ( 
.A1(n_3513),
.A2(n_9),
.A3(n_11),
.B1(n_7),
.B2(n_8),
.C(n_10),
.Y(n_4404)
);

NOR2xp33_ASAP7_75t_L g4405 ( 
.A(n_3663),
.B(n_413),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_3456),
.B(n_414),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_3456),
.B(n_414),
.Y(n_4407)
);

CKINVDCx10_ASAP7_75t_R g4408 ( 
.A(n_3651),
.Y(n_4408)
);

O2A1O1Ixp33_ASAP7_75t_L g4409 ( 
.A1(n_3733),
.A2(n_416),
.B(n_417),
.C(n_415),
.Y(n_4409)
);

AO21x1_ASAP7_75t_L g4410 ( 
.A1(n_3586),
.A2(n_416),
.B(n_415),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_3727),
.B(n_416),
.Y(n_4411)
);

A2O1A1Ixp33_ASAP7_75t_L g4412 ( 
.A1(n_3737),
.A2(n_419),
.B(n_420),
.C(n_418),
.Y(n_4412)
);

AOI22x1_ASAP7_75t_L g4413 ( 
.A1(n_3718),
.A2(n_419),
.B1(n_420),
.B2(n_418),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_3833),
.B(n_418),
.Y(n_4414)
);

OAI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_3534),
.A2(n_422),
.B1(n_423),
.B2(n_420),
.Y(n_4415)
);

OAI21xp5_ASAP7_75t_L g4416 ( 
.A1(n_3515),
.A2(n_424),
.B(n_423),
.Y(n_4416)
);

BUFx4f_ASAP7_75t_L g4417 ( 
.A(n_3883),
.Y(n_4417)
);

OAI21xp5_ASAP7_75t_L g4418 ( 
.A1(n_3826),
.A2(n_425),
.B(n_423),
.Y(n_4418)
);

O2A1O1Ixp33_ASAP7_75t_L g4419 ( 
.A1(n_3938),
.A2(n_426),
.B(n_427),
.C(n_425),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_L g4420 ( 
.A(n_3773),
.B(n_3719),
.Y(n_4420)
);

AND2x6_ASAP7_75t_L g4421 ( 
.A(n_3859),
.B(n_3466),
.Y(n_4421)
);

NOR2xp33_ASAP7_75t_L g4422 ( 
.A(n_3652),
.B(n_425),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_3944),
.Y(n_4423)
);

AOI33xp33_ASAP7_75t_L g4424 ( 
.A1(n_3534),
.A2(n_9),
.A3(n_11),
.B1(n_7),
.B2(n_8),
.B3(n_10),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_3773),
.B(n_426),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_3472),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_3719),
.B(n_427),
.Y(n_4427)
);

BUFx4f_ASAP7_75t_L g4428 ( 
.A(n_3472),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_3853),
.Y(n_4429)
);

CKINVDCx10_ASAP7_75t_R g4430 ( 
.A(n_3531),
.Y(n_4430)
);

OAI22xp5_ASAP7_75t_L g4431 ( 
.A1(n_3549),
.A2(n_428),
.B1(n_429),
.B2(n_427),
.Y(n_4431)
);

AOI21xp5_ASAP7_75t_L g4432 ( 
.A1(n_3838),
.A2(n_429),
.B(n_428),
.Y(n_4432)
);

CKINVDCx10_ASAP7_75t_R g4433 ( 
.A(n_3549),
.Y(n_4433)
);

AND2x2_ASAP7_75t_SL g4434 ( 
.A(n_3671),
.B(n_3477),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_3722),
.B(n_428),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_3477),
.Y(n_4436)
);

O2A1O1Ixp33_ASAP7_75t_L g4437 ( 
.A1(n_3768),
.A2(n_430),
.B(n_431),
.C(n_429),
.Y(n_4437)
);

AOI21xp5_ASAP7_75t_L g4438 ( 
.A1(n_3843),
.A2(n_431),
.B(n_430),
.Y(n_4438)
);

A2O1A1Ixp33_ASAP7_75t_L g4439 ( 
.A1(n_3722),
.A2(n_431),
.B(n_432),
.C(n_430),
.Y(n_4439)
);

NOR2xp33_ASAP7_75t_L g4440 ( 
.A(n_3768),
.B(n_432),
.Y(n_4440)
);

AOI21xp5_ASAP7_75t_L g4441 ( 
.A1(n_3843),
.A2(n_434),
.B(n_433),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_3724),
.B(n_433),
.Y(n_4442)
);

OAI22xp5_ASAP7_75t_L g4443 ( 
.A1(n_3724),
.A2(n_435),
.B1(n_436),
.B2(n_434),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_3734),
.B(n_434),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_3734),
.B(n_435),
.Y(n_4445)
);

OAI21xp5_ASAP7_75t_L g4446 ( 
.A1(n_3746),
.A2(n_437),
.B(n_436),
.Y(n_4446)
);

INVx2_ASAP7_75t_SL g4447 ( 
.A(n_3921),
.Y(n_4447)
);

OAI22xp5_ASAP7_75t_L g4448 ( 
.A1(n_3921),
.A2(n_437),
.B1(n_438),
.B2(n_436),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_SL g4449 ( 
.A(n_3853),
.B(n_438),
.Y(n_4449)
);

NOR2xp33_ASAP7_75t_L g4450 ( 
.A(n_3855),
.B(n_438),
.Y(n_4450)
);

AOI21xp5_ASAP7_75t_L g4451 ( 
.A1(n_3855),
.A2(n_440),
.B(n_439),
.Y(n_4451)
);

BUFx8_ASAP7_75t_L g4452 ( 
.A(n_3563),
.Y(n_4452)
);

CKINVDCx10_ASAP7_75t_R g4453 ( 
.A(n_3563),
.Y(n_4453)
);

AOI21x1_ASAP7_75t_L g4454 ( 
.A1(n_3876),
.A2(n_441),
.B(n_439),
.Y(n_4454)
);

NOR2x1_ASAP7_75t_L g4455 ( 
.A(n_3487),
.B(n_439),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_L g4456 ( 
.A(n_3856),
.B(n_441),
.Y(n_4456)
);

NOR2xp33_ASAP7_75t_L g4457 ( 
.A(n_3856),
.B(n_441),
.Y(n_4457)
);

INVx2_ASAP7_75t_L g4458 ( 
.A(n_3874),
.Y(n_4458)
);

NOR2xp33_ASAP7_75t_L g4459 ( 
.A(n_3874),
.B(n_442),
.Y(n_4459)
);

AOI21xp5_ASAP7_75t_L g4460 ( 
.A1(n_3671),
.A2(n_443),
.B(n_442),
.Y(n_4460)
);

AOI21xp5_ASAP7_75t_L g4461 ( 
.A1(n_3746),
.A2(n_443),
.B(n_442),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_SL g4462 ( 
.A(n_3876),
.B(n_443),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_SL g4463 ( 
.A(n_3487),
.B(n_444),
.Y(n_4463)
);

AOI21xp5_ASAP7_75t_L g4464 ( 
.A1(n_3492),
.A2(n_445),
.B(n_444),
.Y(n_4464)
);

OAI21xp5_ASAP7_75t_L g4465 ( 
.A1(n_3846),
.A2(n_446),
.B(n_445),
.Y(n_4465)
);

NOR2xp33_ASAP7_75t_L g4466 ( 
.A(n_3846),
.B(n_446),
.Y(n_4466)
);

AOI21xp5_ASAP7_75t_L g4467 ( 
.A1(n_3492),
.A2(n_447),
.B(n_446),
.Y(n_4467)
);

AOI21xp5_ASAP7_75t_L g4468 ( 
.A1(n_3495),
.A2(n_448),
.B(n_447),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_L g4469 ( 
.A(n_3574),
.B(n_447),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_3574),
.B(n_448),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_SL g4471 ( 
.A(n_3495),
.B(n_449),
.Y(n_4471)
);

NOR2xp33_ASAP7_75t_L g4472 ( 
.A(n_3847),
.B(n_449),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_3582),
.B(n_3593),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_3497),
.Y(n_4474)
);

AOI21xp5_ASAP7_75t_L g4475 ( 
.A1(n_3497),
.A2(n_450),
.B(n_449),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_3582),
.B(n_450),
.Y(n_4476)
);

AOI21x1_ASAP7_75t_L g4477 ( 
.A1(n_3693),
.A2(n_451),
.B(n_450),
.Y(n_4477)
);

AOI21xp5_ASAP7_75t_L g4478 ( 
.A1(n_3498),
.A2(n_452),
.B(n_451),
.Y(n_4478)
);

AOI21xp5_ASAP7_75t_L g4479 ( 
.A1(n_3498),
.A2(n_452),
.B(n_451),
.Y(n_4479)
);

AOI21xp5_ASAP7_75t_L g4480 ( 
.A1(n_3506),
.A2(n_453),
.B(n_452),
.Y(n_4480)
);

OAI22xp5_ASAP7_75t_L g4481 ( 
.A1(n_3847),
.A2(n_454),
.B1(n_455),
.B2(n_453),
.Y(n_4481)
);

AOI21xp5_ASAP7_75t_L g4482 ( 
.A1(n_3506),
.A2(n_454),
.B(n_453),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_3510),
.Y(n_4483)
);

AOI21x1_ASAP7_75t_L g4484 ( 
.A1(n_3693),
.A2(n_455),
.B(n_454),
.Y(n_4484)
);

AOI21xp5_ASAP7_75t_L g4485 ( 
.A1(n_3510),
.A2(n_3526),
.B(n_3518),
.Y(n_4485)
);

NOR2x1_ASAP7_75t_L g4486 ( 
.A(n_3518),
.B(n_457),
.Y(n_4486)
);

O2A1O1Ixp33_ASAP7_75t_L g4487 ( 
.A1(n_3884),
.A2(n_458),
.B(n_459),
.C(n_457),
.Y(n_4487)
);

AOI21xp5_ASAP7_75t_L g4488 ( 
.A1(n_3526),
.A2(n_458),
.B(n_457),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_3593),
.B(n_458),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_3604),
.B(n_459),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_3604),
.B(n_459),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_3530),
.Y(n_4492)
);

AND2x2_ASAP7_75t_L g4493 ( 
.A(n_3781),
.B(n_1057),
.Y(n_4493)
);

BUFx6f_ASAP7_75t_L g4494 ( 
.A(n_3884),
.Y(n_4494)
);

NAND3xp33_ASAP7_75t_L g4495 ( 
.A(n_3897),
.B(n_1058),
.C(n_1057),
.Y(n_4495)
);

AOI21xp5_ASAP7_75t_L g4496 ( 
.A1(n_3530),
.A2(n_461),
.B(n_460),
.Y(n_4496)
);

INVx2_ASAP7_75t_L g4497 ( 
.A(n_3616),
.Y(n_4497)
);

NOR3xp33_ASAP7_75t_L g4498 ( 
.A(n_3897),
.B(n_461),
.C(n_460),
.Y(n_4498)
);

INVx2_ASAP7_75t_L g4499 ( 
.A(n_3616),
.Y(n_4499)
);

AOI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_3634),
.A2(n_463),
.B(n_462),
.Y(n_4500)
);

O2A1O1Ixp33_ASAP7_75t_L g4501 ( 
.A1(n_3906),
.A2(n_463),
.B(n_464),
.C(n_462),
.Y(n_4501)
);

AOI21xp5_ASAP7_75t_L g4502 ( 
.A1(n_3955),
.A2(n_3642),
.B(n_3634),
.Y(n_4502)
);

BUFx6f_ASAP7_75t_L g4503 ( 
.A(n_4173),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4325),
.B(n_3805),
.Y(n_4504)
);

AOI22xp5_ASAP7_75t_L g4505 ( 
.A1(n_3970),
.A2(n_3913),
.B1(n_3916),
.B2(n_3906),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_L g4506 ( 
.A(n_4001),
.B(n_3781),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4007),
.Y(n_4507)
);

O2A1O1Ixp33_ASAP7_75t_L g4508 ( 
.A1(n_4210),
.A2(n_3916),
.B(n_3913),
.C(n_3791),
.Y(n_4508)
);

AOI21xp5_ASAP7_75t_L g4509 ( 
.A1(n_3962),
.A2(n_3642),
.B(n_3782),
.Y(n_4509)
);

NOR2xp33_ASAP7_75t_L g4510 ( 
.A(n_4217),
.B(n_463),
.Y(n_4510)
);

A2O1A1Ixp33_ASAP7_75t_L g4511 ( 
.A1(n_4428),
.A2(n_3782),
.B(n_3804),
.C(n_3791),
.Y(n_4511)
);

O2A1O1Ixp33_ASAP7_75t_L g4512 ( 
.A1(n_4378),
.A2(n_3804),
.B(n_3807),
.C(n_3805),
.Y(n_4512)
);

NOR2xp33_ASAP7_75t_L g4513 ( 
.A(n_4088),
.B(n_464),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4018),
.Y(n_4514)
);

AOI21xp5_ASAP7_75t_L g4515 ( 
.A1(n_3973),
.A2(n_3807),
.B(n_3774),
.Y(n_4515)
);

OR2x6_ASAP7_75t_L g4516 ( 
.A(n_3967),
.B(n_3774),
.Y(n_4516)
);

NOR2xp33_ASAP7_75t_SL g4517 ( 
.A(n_4244),
.B(n_1066),
.Y(n_4517)
);

O2A1O1Ixp33_ASAP7_75t_L g4518 ( 
.A1(n_3968),
.A2(n_466),
.B(n_467),
.C(n_465),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_SL g4519 ( 
.A(n_4014),
.B(n_465),
.Y(n_4519)
);

BUFx6f_ASAP7_75t_L g4520 ( 
.A(n_4173),
.Y(n_4520)
);

INVx4_ASAP7_75t_L g4521 ( 
.A(n_4065),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4008),
.B(n_465),
.Y(n_4522)
);

O2A1O1Ixp33_ASAP7_75t_L g4523 ( 
.A1(n_3985),
.A2(n_467),
.B(n_468),
.C(n_466),
.Y(n_4523)
);

A2O1A1Ixp33_ASAP7_75t_L g4524 ( 
.A1(n_4428),
.A2(n_467),
.B(n_468),
.C(n_466),
.Y(n_4524)
);

AND2x4_ASAP7_75t_L g4525 ( 
.A(n_4155),
.B(n_468),
.Y(n_4525)
);

O2A1O1Ixp33_ASAP7_75t_L g4526 ( 
.A1(n_3991),
.A2(n_470),
.B(n_471),
.C(n_469),
.Y(n_4526)
);

AOI21xp5_ASAP7_75t_L g4527 ( 
.A1(n_3984),
.A2(n_470),
.B(n_469),
.Y(n_4527)
);

NOR2xp33_ASAP7_75t_L g4528 ( 
.A(n_4301),
.B(n_4453),
.Y(n_4528)
);

CKINVDCx5p33_ASAP7_75t_R g4529 ( 
.A(n_4125),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4027),
.Y(n_4530)
);

AOI22xp33_ASAP7_75t_L g4531 ( 
.A1(n_4452),
.A2(n_472),
.B1(n_473),
.B2(n_471),
.Y(n_4531)
);

INVx2_ASAP7_75t_L g4532 ( 
.A(n_3989),
.Y(n_4532)
);

BUFx6f_ASAP7_75t_L g4533 ( 
.A(n_4173),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_SL g4534 ( 
.A(n_4014),
.B(n_471),
.Y(n_4534)
);

AOI21xp5_ASAP7_75t_L g4535 ( 
.A1(n_3987),
.A2(n_473),
.B(n_472),
.Y(n_4535)
);

HB1xp67_ASAP7_75t_L g4536 ( 
.A(n_3956),
.Y(n_4536)
);

NOR2xp33_ASAP7_75t_SL g4537 ( 
.A(n_3972),
.B(n_4060),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_3990),
.Y(n_4538)
);

AOI21xp5_ASAP7_75t_L g4539 ( 
.A1(n_3996),
.A2(n_473),
.B(n_472),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4044),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4093),
.B(n_474),
.Y(n_4541)
);

OAI22x1_ASAP7_75t_L g4542 ( 
.A1(n_3972),
.A2(n_476),
.B1(n_477),
.B2(n_475),
.Y(n_4542)
);

AOI21xp5_ASAP7_75t_L g4543 ( 
.A1(n_4061),
.A2(n_476),
.B(n_475),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_3994),
.Y(n_4544)
);

OAI22xp5_ASAP7_75t_L g4545 ( 
.A1(n_4333),
.A2(n_4375),
.B1(n_4359),
.B2(n_4434),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4037),
.B(n_475),
.Y(n_4546)
);

O2A1O1Ixp33_ASAP7_75t_L g4547 ( 
.A1(n_4138),
.A2(n_477),
.B(n_478),
.C(n_476),
.Y(n_4547)
);

NOR2x1p5_ASAP7_75t_L g4548 ( 
.A(n_4206),
.B(n_477),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4057),
.Y(n_4549)
);

INVx3_ASAP7_75t_L g4550 ( 
.A(n_4364),
.Y(n_4550)
);

A2O1A1Ixp33_ASAP7_75t_L g4551 ( 
.A1(n_4164),
.A2(n_479),
.B(n_480),
.C(n_478),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4070),
.Y(n_4552)
);

OAI21x1_ASAP7_75t_L g4553 ( 
.A1(n_3964),
.A2(n_3971),
.B(n_4046),
.Y(n_4553)
);

AOI21xp5_ASAP7_75t_L g4554 ( 
.A1(n_4098),
.A2(n_3977),
.B(n_3965),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4022),
.Y(n_4555)
);

OAI22xp5_ASAP7_75t_L g4556 ( 
.A1(n_4060),
.A2(n_479),
.B1(n_481),
.B2(n_478),
.Y(n_4556)
);

CKINVDCx6p67_ASAP7_75t_R g4557 ( 
.A(n_4053),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4038),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4335),
.B(n_481),
.Y(n_4559)
);

OAI22xp5_ASAP7_75t_L g4560 ( 
.A1(n_4417),
.A2(n_482),
.B1(n_483),
.B2(n_481),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_4091),
.Y(n_4561)
);

BUFx2_ASAP7_75t_L g4562 ( 
.A(n_4246),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4095),
.Y(n_4563)
);

OAI22xp5_ASAP7_75t_SL g4564 ( 
.A1(n_4191),
.A2(n_483),
.B1(n_484),
.B2(n_482),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_4079),
.A2(n_483),
.B(n_482),
.Y(n_4565)
);

INVx3_ASAP7_75t_L g4566 ( 
.A(n_4364),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4100),
.Y(n_4567)
);

AOI21xp5_ASAP7_75t_L g4568 ( 
.A1(n_4023),
.A2(n_485),
.B(n_484),
.Y(n_4568)
);

AOI21xp5_ASAP7_75t_L g4569 ( 
.A1(n_4028),
.A2(n_485),
.B(n_484),
.Y(n_4569)
);

NOR2xp33_ASAP7_75t_L g4570 ( 
.A(n_4433),
.B(n_485),
.Y(n_4570)
);

O2A1O1Ixp33_ASAP7_75t_L g4571 ( 
.A1(n_4439),
.A2(n_488),
.B(n_489),
.C(n_487),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_L g4572 ( 
.A(n_4104),
.B(n_487),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_L g4573 ( 
.A(n_4113),
.B(n_487),
.Y(n_4573)
);

NOR2xp33_ASAP7_75t_L g4574 ( 
.A(n_4361),
.B(n_488),
.Y(n_4574)
);

BUFx3_ASAP7_75t_L g4575 ( 
.A(n_4143),
.Y(n_4575)
);

BUFx6f_ASAP7_75t_L g4576 ( 
.A(n_4246),
.Y(n_4576)
);

AOI21xp5_ASAP7_75t_L g4577 ( 
.A1(n_4040),
.A2(n_489),
.B(n_488),
.Y(n_4577)
);

AOI21xp5_ASAP7_75t_L g4578 ( 
.A1(n_3974),
.A2(n_490),
.B(n_489),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_4114),
.B(n_491),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4141),
.Y(n_4580)
);

INVx2_ASAP7_75t_L g4581 ( 
.A(n_4140),
.Y(n_4581)
);

O2A1O1Ixp5_ASAP7_75t_L g4582 ( 
.A1(n_4089),
.A2(n_492),
.B(n_493),
.C(n_491),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4146),
.B(n_492),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4167),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4172),
.B(n_493),
.Y(n_4585)
);

NOR2xp33_ASAP7_75t_L g4586 ( 
.A(n_4005),
.B(n_493),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4175),
.B(n_494),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4192),
.Y(n_4588)
);

AOI21xp5_ASAP7_75t_L g4589 ( 
.A1(n_4030),
.A2(n_495),
.B(n_494),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_4225),
.B(n_4249),
.Y(n_4590)
);

AND2x2_ASAP7_75t_L g4591 ( 
.A(n_4020),
.B(n_495),
.Y(n_4591)
);

NOR2xp33_ASAP7_75t_L g4592 ( 
.A(n_3961),
.B(n_495),
.Y(n_4592)
);

O2A1O1Ixp33_ASAP7_75t_L g4593 ( 
.A1(n_3997),
.A2(n_497),
.B(n_498),
.C(n_496),
.Y(n_4593)
);

AOI21xp5_ASAP7_75t_L g4594 ( 
.A1(n_4012),
.A2(n_497),
.B(n_496),
.Y(n_4594)
);

NOR3xp33_ASAP7_75t_L g4595 ( 
.A(n_4402),
.B(n_4407),
.C(n_4406),
.Y(n_4595)
);

AOI21xp5_ASAP7_75t_L g4596 ( 
.A1(n_4077),
.A2(n_499),
.B(n_498),
.Y(n_4596)
);

AO21x1_ASAP7_75t_L g4597 ( 
.A1(n_4485),
.A2(n_499),
.B(n_498),
.Y(n_4597)
);

NOR2xp67_ASAP7_75t_L g4598 ( 
.A(n_4014),
.B(n_504),
.Y(n_4598)
);

O2A1O1Ixp5_ASAP7_75t_L g4599 ( 
.A1(n_4123),
.A2(n_500),
.B(n_501),
.C(n_499),
.Y(n_4599)
);

INVx3_ASAP7_75t_L g4600 ( 
.A(n_4047),
.Y(n_4600)
);

O2A1O1Ixp33_ASAP7_75t_L g4601 ( 
.A1(n_4278),
.A2(n_501),
.B(n_502),
.C(n_500),
.Y(n_4601)
);

NOR3xp33_ASAP7_75t_SL g4602 ( 
.A(n_4171),
.B(n_503),
.C(n_502),
.Y(n_4602)
);

AOI21xp5_ASAP7_75t_L g4603 ( 
.A1(n_4120),
.A2(n_504),
.B(n_503),
.Y(n_4603)
);

NAND2xp5_ASAP7_75t_SL g4604 ( 
.A(n_4155),
.B(n_504),
.Y(n_4604)
);

A2O1A1Ixp33_ASAP7_75t_L g4605 ( 
.A1(n_4338),
.A2(n_506),
.B(n_507),
.C(n_505),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_SL g4606 ( 
.A(n_4157),
.B(n_506),
.Y(n_4606)
);

NOR2xp67_ASAP7_75t_L g4607 ( 
.A(n_4047),
.B(n_513),
.Y(n_4607)
);

INVx1_ASAP7_75t_SL g4608 ( 
.A(n_4068),
.Y(n_4608)
);

OAI22xp5_ASAP7_75t_L g4609 ( 
.A1(n_4417),
.A2(n_508),
.B1(n_509),
.B2(n_507),
.Y(n_4609)
);

AOI21xp5_ASAP7_75t_L g4610 ( 
.A1(n_4045),
.A2(n_508),
.B(n_507),
.Y(n_4610)
);

AOI22xp33_ASAP7_75t_L g4611 ( 
.A1(n_4452),
.A2(n_511),
.B1(n_512),
.B2(n_509),
.Y(n_4611)
);

INVx1_ASAP7_75t_SL g4612 ( 
.A(n_4143),
.Y(n_4612)
);

AOI21xp5_ASAP7_75t_L g4613 ( 
.A1(n_3975),
.A2(n_512),
.B(n_511),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_SL g4614 ( 
.A(n_4157),
.B(n_511),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_L g4615 ( 
.A(n_4259),
.B(n_513),
.Y(n_4615)
);

OAI22xp5_ASAP7_75t_L g4616 ( 
.A1(n_4218),
.A2(n_4379),
.B1(n_4242),
.B2(n_4257),
.Y(n_4616)
);

A2O1A1Ixp33_ASAP7_75t_SL g4617 ( 
.A1(n_4450),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_4267),
.B(n_4274),
.Y(n_4618)
);

OAI21xp5_ASAP7_75t_L g4619 ( 
.A1(n_4149),
.A2(n_4271),
.B(n_4251),
.Y(n_4619)
);

AOI21xp5_ASAP7_75t_L g4620 ( 
.A1(n_4052),
.A2(n_514),
.B(n_513),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_4282),
.B(n_514),
.Y(n_4621)
);

O2A1O1Ixp33_ASAP7_75t_L g4622 ( 
.A1(n_4208),
.A2(n_515),
.B(n_516),
.C(n_514),
.Y(n_4622)
);

INVx2_ASAP7_75t_SL g4623 ( 
.A(n_4143),
.Y(n_4623)
);

NOR2xp33_ASAP7_75t_SL g4624 ( 
.A(n_3960),
.B(n_1069),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4291),
.Y(n_4625)
);

NOR2xp33_ASAP7_75t_L g4626 ( 
.A(n_4383),
.B(n_515),
.Y(n_4626)
);

A2O1A1Ixp33_ASAP7_75t_SL g4627 ( 
.A1(n_4457),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4075),
.B(n_515),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4160),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4305),
.B(n_517),
.Y(n_4630)
);

A2O1A1Ixp33_ASAP7_75t_L g4631 ( 
.A1(n_4382),
.A2(n_518),
.B(n_519),
.C(n_517),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4127),
.B(n_519),
.Y(n_4632)
);

BUFx4f_ASAP7_75t_L g4633 ( 
.A(n_3958),
.Y(n_4633)
);

AOI21xp5_ASAP7_75t_L g4634 ( 
.A1(n_3976),
.A2(n_520),
.B(n_519),
.Y(n_4634)
);

INVx1_ASAP7_75t_SL g4635 ( 
.A(n_4145),
.Y(n_4635)
);

O2A1O1Ixp33_ASAP7_75t_L g4636 ( 
.A1(n_3981),
.A2(n_521),
.B(n_522),
.C(n_520),
.Y(n_4636)
);

OAI22xp5_ASAP7_75t_L g4637 ( 
.A1(n_4418),
.A2(n_521),
.B1(n_522),
.B2(n_520),
.Y(n_4637)
);

BUFx6f_ASAP7_75t_L g4638 ( 
.A(n_4246),
.Y(n_4638)
);

INVx3_ASAP7_75t_L g4639 ( 
.A(n_4383),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4312),
.B(n_521),
.Y(n_4640)
);

NAND2xp5_ASAP7_75t_L g4641 ( 
.A(n_4343),
.B(n_522),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_4362),
.B(n_523),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_3998),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4328),
.B(n_523),
.Y(n_4644)
);

INVx3_ASAP7_75t_SL g4645 ( 
.A(n_3979),
.Y(n_4645)
);

NOR2xp33_ASAP7_75t_L g4646 ( 
.A(n_4124),
.B(n_523),
.Y(n_4646)
);

OAI21x1_ASAP7_75t_L g4647 ( 
.A1(n_3978),
.A2(n_525),
.B(n_524),
.Y(n_4647)
);

BUFx6f_ASAP7_75t_L g4648 ( 
.A(n_4145),
.Y(n_4648)
);

O2A1O1Ixp5_ASAP7_75t_L g4649 ( 
.A1(n_4462),
.A2(n_3959),
.B(n_4449),
.C(n_4062),
.Y(n_4649)
);

A2O1A1Ixp33_ASAP7_75t_SL g4650 ( 
.A1(n_4459),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4298),
.B(n_524),
.Y(n_4651)
);

NAND2xp5_ASAP7_75t_SL g4652 ( 
.A(n_4494),
.B(n_524),
.Y(n_4652)
);

AOI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_4041),
.A2(n_527),
.B(n_525),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4298),
.B(n_525),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_4109),
.B(n_527),
.Y(n_4655)
);

BUFx3_ASAP7_75t_L g4656 ( 
.A(n_4145),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4202),
.Y(n_4657)
);

O2A1O1Ixp33_ASAP7_75t_L g4658 ( 
.A1(n_4117),
.A2(n_528),
.B(n_529),
.C(n_527),
.Y(n_4658)
);

INVx2_ASAP7_75t_L g4659 ( 
.A(n_4162),
.Y(n_4659)
);

OR2x2_ASAP7_75t_L g4660 ( 
.A(n_4294),
.B(n_528),
.Y(n_4660)
);

NAND2xp5_ASAP7_75t_SL g4661 ( 
.A(n_4494),
.B(n_528),
.Y(n_4661)
);

BUFx6f_ASAP7_75t_L g4662 ( 
.A(n_4031),
.Y(n_4662)
);

AND2x2_ASAP7_75t_L g4663 ( 
.A(n_4318),
.B(n_529),
.Y(n_4663)
);

AOI21xp5_ASAP7_75t_L g4664 ( 
.A1(n_3982),
.A2(n_530),
.B(n_529),
.Y(n_4664)
);

OAI22xp5_ASAP7_75t_L g4665 ( 
.A1(n_4295),
.A2(n_531),
.B1(n_532),
.B2(n_530),
.Y(n_4665)
);

AOI21x1_ASAP7_75t_L g4666 ( 
.A1(n_3999),
.A2(n_531),
.B(n_530),
.Y(n_4666)
);

HB1xp67_ASAP7_75t_L g4667 ( 
.A(n_4307),
.Y(n_4667)
);

INVx1_ASAP7_75t_SL g4668 ( 
.A(n_4003),
.Y(n_4668)
);

INVxp67_ASAP7_75t_SL g4669 ( 
.A(n_4474),
.Y(n_4669)
);

O2A1O1Ixp33_ASAP7_75t_L g4670 ( 
.A1(n_4128),
.A2(n_532),
.B(n_533),
.C(n_531),
.Y(n_4670)
);

AOI21xp5_ASAP7_75t_L g4671 ( 
.A1(n_3983),
.A2(n_533),
.B(n_532),
.Y(n_4671)
);

OAI21xp33_ASAP7_75t_SL g4672 ( 
.A1(n_4455),
.A2(n_4486),
.B(n_4471),
.Y(n_4672)
);

BUFx6f_ASAP7_75t_L g4673 ( 
.A(n_4031),
.Y(n_4673)
);

AOI21xp5_ASAP7_75t_L g4674 ( 
.A1(n_4016),
.A2(n_534),
.B(n_533),
.Y(n_4674)
);

CKINVDCx8_ASAP7_75t_R g4675 ( 
.A(n_4372),
.Y(n_4675)
);

NOR2xp67_ASAP7_75t_L g4676 ( 
.A(n_4103),
.B(n_536),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4235),
.B(n_535),
.Y(n_4677)
);

NOR2x1p5_ASAP7_75t_L g4678 ( 
.A(n_4103),
.B(n_535),
.Y(n_4678)
);

INVx2_ASAP7_75t_SL g4679 ( 
.A(n_3960),
.Y(n_4679)
);

OAI21x1_ASAP7_75t_L g4680 ( 
.A1(n_4009),
.A2(n_536),
.B(n_535),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_SL g4681 ( 
.A(n_4494),
.B(n_536),
.Y(n_4681)
);

INVx5_ASAP7_75t_L g4682 ( 
.A(n_4346),
.Y(n_4682)
);

O2A1O1Ixp33_ASAP7_75t_SL g4683 ( 
.A1(n_4463),
.A2(n_4153),
.B(n_4337),
.C(n_4327),
.Y(n_4683)
);

AOI21xp5_ASAP7_75t_L g4684 ( 
.A1(n_4021),
.A2(n_538),
.B(n_537),
.Y(n_4684)
);

BUFx12f_ASAP7_75t_L g4685 ( 
.A(n_4367),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4254),
.B(n_537),
.Y(n_4686)
);

NAND3xp33_ASAP7_75t_L g4687 ( 
.A(n_4498),
.B(n_538),
.C(n_537),
.Y(n_4687)
);

INVxp67_ASAP7_75t_L g4688 ( 
.A(n_4196),
.Y(n_4688)
);

INVx2_ASAP7_75t_L g4689 ( 
.A(n_4237),
.Y(n_4689)
);

INVx2_ASAP7_75t_L g4690 ( 
.A(n_4256),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_4368),
.B(n_538),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_4473),
.B(n_539),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4036),
.B(n_539),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_SL g4694 ( 
.A(n_4006),
.B(n_540),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_SL g4695 ( 
.A(n_4006),
.B(n_540),
.Y(n_4695)
);

BUFx2_ASAP7_75t_L g4696 ( 
.A(n_3992),
.Y(n_4696)
);

AND2x2_ASAP7_75t_L g4697 ( 
.A(n_4332),
.B(n_540),
.Y(n_4697)
);

NAND2xp5_ASAP7_75t_L g4698 ( 
.A(n_4349),
.B(n_541),
.Y(n_4698)
);

AOI21xp5_ASAP7_75t_L g4699 ( 
.A1(n_4092),
.A2(n_542),
.B(n_541),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4376),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_L g4701 ( 
.A(n_4358),
.B(n_541),
.Y(n_4701)
);

O2A1O1Ixp33_ASAP7_75t_L g4702 ( 
.A1(n_4147),
.A2(n_543),
.B(n_544),
.C(n_542),
.Y(n_4702)
);

BUFx6f_ASAP7_75t_L g4703 ( 
.A(n_4031),
.Y(n_4703)
);

NOR2xp33_ASAP7_75t_SL g4704 ( 
.A(n_4063),
.B(n_1065),
.Y(n_4704)
);

NOR2xp33_ASAP7_75t_R g4705 ( 
.A(n_4261),
.B(n_1064),
.Y(n_4705)
);

INVx5_ASAP7_75t_L g4706 ( 
.A(n_4346),
.Y(n_4706)
);

NAND3xp33_ASAP7_75t_L g4707 ( 
.A(n_4356),
.B(n_544),
.C(n_543),
.Y(n_4707)
);

BUFx12f_ASAP7_75t_L g4708 ( 
.A(n_4389),
.Y(n_4708)
);

OAI21x1_ASAP7_75t_L g4709 ( 
.A1(n_4010),
.A2(n_544),
.B(n_543),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4377),
.B(n_545),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4069),
.Y(n_4711)
);

OR2x2_ASAP7_75t_L g4712 ( 
.A(n_4094),
.B(n_545),
.Y(n_4712)
);

INVx2_ASAP7_75t_SL g4713 ( 
.A(n_4268),
.Y(n_4713)
);

OAI21x1_ASAP7_75t_L g4714 ( 
.A1(n_4108),
.A2(n_547),
.B(n_546),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_4231),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4207),
.B(n_546),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_SL g4717 ( 
.A(n_4078),
.B(n_546),
.Y(n_4717)
);

AO32x2_ASAP7_75t_L g4718 ( 
.A1(n_4447),
.A2(n_564),
.A3(n_572),
.B1(n_556),
.B2(n_548),
.Y(n_4718)
);

NOR2xp33_ASAP7_75t_L g4719 ( 
.A(n_4322),
.B(n_547),
.Y(n_4719)
);

O2A1O1Ixp5_ASAP7_75t_L g4720 ( 
.A1(n_4135),
.A2(n_549),
.B(n_550),
.C(n_548),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_SL g4721 ( 
.A(n_4290),
.B(n_549),
.Y(n_4721)
);

INVx2_ASAP7_75t_L g4722 ( 
.A(n_4233),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4273),
.Y(n_4723)
);

NAND2xp5_ASAP7_75t_L g4724 ( 
.A(n_4071),
.B(n_549),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_SL g4725 ( 
.A(n_4290),
.B(n_551),
.Y(n_4725)
);

O2A1O1Ixp33_ASAP7_75t_L g4726 ( 
.A1(n_4168),
.A2(n_553),
.B(n_554),
.C(n_552),
.Y(n_4726)
);

INVx3_ASAP7_75t_L g4727 ( 
.A(n_4236),
.Y(n_4727)
);

AOI21xp5_ASAP7_75t_L g4728 ( 
.A1(n_4105),
.A2(n_553),
.B(n_552),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_SL g4729 ( 
.A(n_4290),
.B(n_552),
.Y(n_4729)
);

A2O1A1Ixp33_ASAP7_75t_L g4730 ( 
.A1(n_4424),
.A2(n_4501),
.B(n_4487),
.C(n_4437),
.Y(n_4730)
);

AOI21xp5_ASAP7_75t_L g4731 ( 
.A1(n_4043),
.A2(n_555),
.B(n_554),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_SL g4732 ( 
.A(n_4315),
.B(n_4072),
.Y(n_4732)
);

NOR2xp33_ASAP7_75t_SL g4733 ( 
.A(n_4268),
.B(n_1060),
.Y(n_4733)
);

AOI22xp33_ASAP7_75t_SL g4734 ( 
.A1(n_4421),
.A2(n_556),
.B1(n_557),
.B2(n_555),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_SL g4735 ( 
.A(n_4315),
.B(n_555),
.Y(n_4735)
);

BUFx8_ASAP7_75t_L g4736 ( 
.A(n_4285),
.Y(n_4736)
);

INVx5_ASAP7_75t_L g4737 ( 
.A(n_4346),
.Y(n_4737)
);

O2A1O1Ixp33_ASAP7_75t_L g4738 ( 
.A1(n_4306),
.A2(n_557),
.B(n_558),
.C(n_556),
.Y(n_4738)
);

NAND2xp5_ASAP7_75t_L g4739 ( 
.A(n_4035),
.B(n_557),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_3995),
.Y(n_4740)
);

AOI21x1_ASAP7_75t_L g4741 ( 
.A1(n_4131),
.A2(n_559),
.B(n_558),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4055),
.B(n_559),
.Y(n_4742)
);

NOR2xp33_ASAP7_75t_L g4743 ( 
.A(n_4357),
.B(n_559),
.Y(n_4743)
);

OAI21xp5_ASAP7_75t_L g4744 ( 
.A1(n_4188),
.A2(n_561),
.B(n_560),
.Y(n_4744)
);

CKINVDCx5p33_ASAP7_75t_R g4745 ( 
.A(n_4389),
.Y(n_4745)
);

AOI21xp5_ASAP7_75t_L g4746 ( 
.A1(n_4087),
.A2(n_561),
.B(n_560),
.Y(n_4746)
);

AOI21xp5_ASAP7_75t_L g4747 ( 
.A1(n_3980),
.A2(n_562),
.B(n_560),
.Y(n_4747)
);

NOR2xp33_ASAP7_75t_R g4748 ( 
.A(n_4430),
.B(n_1072),
.Y(n_4748)
);

INVx2_ASAP7_75t_L g4749 ( 
.A(n_3995),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4265),
.Y(n_4750)
);

AOI21xp5_ASAP7_75t_L g4751 ( 
.A1(n_4080),
.A2(n_563),
.B(n_562),
.Y(n_4751)
);

AND2x4_ASAP7_75t_L g4752 ( 
.A(n_4397),
.B(n_562),
.Y(n_4752)
);

OAI22xp5_ASAP7_75t_L g4753 ( 
.A1(n_4495),
.A2(n_4200),
.B1(n_4260),
.B2(n_4391),
.Y(n_4753)
);

CKINVDCx20_ASAP7_75t_R g4754 ( 
.A(n_4165),
.Y(n_4754)
);

AOI21xp5_ASAP7_75t_L g4755 ( 
.A1(n_4081),
.A2(n_564),
.B(n_563),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_SL g4756 ( 
.A(n_4315),
.B(n_564),
.Y(n_4756)
);

O2A1O1Ixp5_ASAP7_75t_L g4757 ( 
.A1(n_4309),
.A2(n_566),
.B(n_567),
.C(n_565),
.Y(n_4757)
);

BUFx3_ASAP7_75t_L g4758 ( 
.A(n_4086),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4000),
.B(n_565),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4265),
.Y(n_4760)
);

BUFx3_ASAP7_75t_L g4761 ( 
.A(n_4275),
.Y(n_4761)
);

AND2x2_ASAP7_75t_L g4762 ( 
.A(n_4180),
.B(n_566),
.Y(n_4762)
);

NOR2x1_ASAP7_75t_L g4763 ( 
.A(n_4129),
.B(n_566),
.Y(n_4763)
);

O2A1O1Ixp33_ASAP7_75t_L g4764 ( 
.A1(n_4371),
.A2(n_568),
.B(n_569),
.C(n_567),
.Y(n_4764)
);

BUFx3_ASAP7_75t_L g4765 ( 
.A(n_4275),
.Y(n_4765)
);

BUFx6f_ASAP7_75t_L g4766 ( 
.A(n_3995),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_SL g4767 ( 
.A(n_4248),
.B(n_567),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4002),
.Y(n_4768)
);

AOI22xp33_ASAP7_75t_L g4769 ( 
.A1(n_4421),
.A2(n_569),
.B1(n_570),
.B2(n_568),
.Y(n_4769)
);

AOI21x1_ASAP7_75t_L g4770 ( 
.A1(n_4019),
.A2(n_570),
.B(n_568),
.Y(n_4770)
);

AOI22xp33_ASAP7_75t_L g4771 ( 
.A1(n_4421),
.A2(n_571),
.B1(n_572),
.B2(n_570),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4369),
.Y(n_4772)
);

BUFx3_ASAP7_75t_L g4773 ( 
.A(n_4275),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_L g4774 ( 
.A(n_4493),
.B(n_571),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_3966),
.B(n_571),
.Y(n_4775)
);

INVxp67_ASAP7_75t_SL g4776 ( 
.A(n_4497),
.Y(n_4776)
);

AND2x2_ASAP7_75t_L g4777 ( 
.A(n_4369),
.B(n_573),
.Y(n_4777)
);

AO32x2_ASAP7_75t_L g4778 ( 
.A1(n_4269),
.A2(n_590),
.A3(n_598),
.B1(n_582),
.B2(n_574),
.Y(n_4778)
);

A2O1A1Ixp33_ASAP7_75t_L g4779 ( 
.A1(n_4189),
.A2(n_574),
.B(n_575),
.C(n_573),
.Y(n_4779)
);

AOI22xp5_ASAP7_75t_L g4780 ( 
.A1(n_4373),
.A2(n_1067),
.B1(n_1068),
.B2(n_1066),
.Y(n_4780)
);

AOI21xp5_ASAP7_75t_L g4781 ( 
.A1(n_4084),
.A2(n_575),
.B(n_573),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_3988),
.B(n_3957),
.Y(n_4782)
);

INVx2_ASAP7_75t_L g4783 ( 
.A(n_4002),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_SL g4784 ( 
.A(n_4248),
.B(n_576),
.Y(n_4784)
);

O2A1O1Ixp33_ASAP7_75t_L g4785 ( 
.A1(n_4297),
.A2(n_578),
.B(n_579),
.C(n_577),
.Y(n_4785)
);

NOR2xp33_ASAP7_75t_L g4786 ( 
.A(n_3993),
.B(n_577),
.Y(n_4786)
);

AOI22xp5_ASAP7_75t_L g4787 ( 
.A1(n_4346),
.A2(n_1074),
.B1(n_1072),
.B2(n_578),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_L g4788 ( 
.A(n_4313),
.B(n_577),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4420),
.B(n_579),
.Y(n_4789)
);

INVx5_ASAP7_75t_L g4790 ( 
.A(n_4002),
.Y(n_4790)
);

O2A1O1Ixp33_ASAP7_75t_L g4791 ( 
.A1(n_4308),
.A2(n_580),
.B(n_581),
.C(n_579),
.Y(n_4791)
);

OAI22xp5_ASAP7_75t_L g4792 ( 
.A1(n_4398),
.A2(n_581),
.B1(n_582),
.B2(n_580),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4216),
.Y(n_4793)
);

OAI22xp5_ASAP7_75t_L g4794 ( 
.A1(n_4385),
.A2(n_581),
.B1(n_582),
.B2(n_580),
.Y(n_4794)
);

AOI33xp33_ASAP7_75t_L g4795 ( 
.A1(n_4252),
.A2(n_14),
.A3(n_16),
.B1(n_12),
.B2(n_13),
.B3(n_15),
.Y(n_4795)
);

INVxp67_ASAP7_75t_L g4796 ( 
.A(n_4073),
.Y(n_4796)
);

A2O1A1Ixp33_ASAP7_75t_L g4797 ( 
.A1(n_4205),
.A2(n_584),
.B(n_585),
.C(n_583),
.Y(n_4797)
);

AOI21xp5_ASAP7_75t_L g4798 ( 
.A1(n_4279),
.A2(n_584),
.B(n_583),
.Y(n_4798)
);

NAND2x1p5_ASAP7_75t_L g4799 ( 
.A(n_4116),
.B(n_583),
.Y(n_4799)
);

AOI21xp5_ASAP7_75t_L g4800 ( 
.A1(n_4042),
.A2(n_585),
.B(n_584),
.Y(n_4800)
);

BUFx12f_ASAP7_75t_L g4801 ( 
.A(n_4198),
.Y(n_4801)
);

AOI21xp5_ASAP7_75t_L g4802 ( 
.A1(n_4076),
.A2(n_586),
.B(n_585),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_4413),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4032),
.B(n_586),
.Y(n_4804)
);

A2O1A1Ixp33_ASAP7_75t_L g4805 ( 
.A1(n_4293),
.A2(n_587),
.B(n_588),
.C(n_586),
.Y(n_4805)
);

INVx2_ASAP7_75t_L g4806 ( 
.A(n_4352),
.Y(n_4806)
);

BUFx2_ASAP7_75t_L g4807 ( 
.A(n_4248),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_4085),
.B(n_587),
.Y(n_4808)
);

BUFx6f_ASAP7_75t_L g4809 ( 
.A(n_4121),
.Y(n_4809)
);

NOR2xp33_ASAP7_75t_R g4810 ( 
.A(n_4408),
.B(n_1061),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4469),
.Y(n_4811)
);

BUFx6f_ASAP7_75t_L g4812 ( 
.A(n_4121),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_SL g4813 ( 
.A(n_4281),
.B(n_4121),
.Y(n_4813)
);

CKINVDCx8_ASAP7_75t_R g4814 ( 
.A(n_4198),
.Y(n_4814)
);

NAND2x1p5_ASAP7_75t_L g4815 ( 
.A(n_4334),
.B(n_587),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4097),
.B(n_589),
.Y(n_4816)
);

HB1xp67_ASAP7_75t_L g4817 ( 
.A(n_3986),
.Y(n_4817)
);

OAI22xp5_ASAP7_75t_L g4818 ( 
.A1(n_4340),
.A2(n_590),
.B1(n_591),
.B2(n_589),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4470),
.Y(n_4819)
);

BUFx6f_ASAP7_75t_L g4820 ( 
.A(n_4106),
.Y(n_4820)
);

AOI21x1_ASAP7_75t_L g4821 ( 
.A1(n_4250),
.A2(n_590),
.B(n_589),
.Y(n_4821)
);

AND2x4_ASAP7_75t_SL g4822 ( 
.A(n_4324),
.B(n_591),
.Y(n_4822)
);

NAND2x1p5_ASAP7_75t_L g4823 ( 
.A(n_4303),
.B(n_592),
.Y(n_4823)
);

AND2x2_ASAP7_75t_L g4824 ( 
.A(n_4134),
.B(n_592),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4476),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4101),
.B(n_4425),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4212),
.B(n_592),
.Y(n_4827)
);

CKINVDCx16_ASAP7_75t_R g4828 ( 
.A(n_4194),
.Y(n_4828)
);

AOI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_4166),
.A2(n_594),
.B(n_593),
.Y(n_4829)
);

OAI22x1_ASAP7_75t_L g4830 ( 
.A1(n_4215),
.A2(n_594),
.B1(n_595),
.B2(n_593),
.Y(n_4830)
);

NOR3xp33_ASAP7_75t_SL g4831 ( 
.A(n_4199),
.B(n_596),
.C(n_593),
.Y(n_4831)
);

BUFx2_ASAP7_75t_L g4832 ( 
.A(n_4281),
.Y(n_4832)
);

O2A1O1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_4415),
.A2(n_4431),
.B(n_4151),
.C(n_4392),
.Y(n_4833)
);

INVxp67_ASAP7_75t_SL g4834 ( 
.A(n_4499),
.Y(n_4834)
);

INVx2_ASAP7_75t_SL g4835 ( 
.A(n_4134),
.Y(n_4835)
);

BUFx6f_ASAP7_75t_L g4836 ( 
.A(n_4102),
.Y(n_4836)
);

INVx2_ASAP7_75t_L g4837 ( 
.A(n_4258),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_SL g4838 ( 
.A(n_4460),
.B(n_596),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4238),
.B(n_596),
.Y(n_4839)
);

AOI21xp5_ASAP7_75t_L g4840 ( 
.A1(n_4011),
.A2(n_598),
.B(n_597),
.Y(n_4840)
);

AOI21x1_ASAP7_75t_L g4841 ( 
.A1(n_4142),
.A2(n_599),
.B(n_597),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_L g4842 ( 
.A(n_4489),
.B(n_599),
.Y(n_4842)
);

NAND3xp33_ASAP7_75t_L g4843 ( 
.A(n_4440),
.B(n_601),
.C(n_600),
.Y(n_4843)
);

O2A1O1Ixp33_ASAP7_75t_L g4844 ( 
.A1(n_4412),
.A2(n_601),
.B(n_602),
.C(n_600),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4490),
.B(n_600),
.Y(n_4845)
);

A2O1A1Ixp33_ASAP7_75t_L g4846 ( 
.A1(n_4341),
.A2(n_603),
.B(n_604),
.C(n_602),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_L g4847 ( 
.A(n_4491),
.B(n_602),
.Y(n_4847)
);

NAND2xp5_ASAP7_75t_L g4848 ( 
.A(n_4110),
.B(n_603),
.Y(n_4848)
);

CKINVDCx14_ASAP7_75t_R g4849 ( 
.A(n_4220),
.Y(n_4849)
);

NOR2xp33_ASAP7_75t_L g4850 ( 
.A(n_4370),
.B(n_4099),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4386),
.Y(n_4851)
);

INVx4_ASAP7_75t_L g4852 ( 
.A(n_4148),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4426),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4436),
.Y(n_4854)
);

AO21x2_ASAP7_75t_L g4855 ( 
.A1(n_4465),
.A2(n_4446),
.B(n_4400),
.Y(n_4855)
);

HB1xp67_ASAP7_75t_L g4856 ( 
.A(n_4388),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4115),
.B(n_603),
.Y(n_4857)
);

OAI22xp5_ASAP7_75t_L g4858 ( 
.A1(n_4136),
.A2(n_4181),
.B1(n_4213),
.B2(n_4144),
.Y(n_4858)
);

AND2x4_ASAP7_75t_L g4859 ( 
.A(n_4483),
.B(n_604),
.Y(n_4859)
);

BUFx2_ASAP7_75t_L g4860 ( 
.A(n_4421),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_SL g4861 ( 
.A(n_4380),
.B(n_604),
.Y(n_4861)
);

AOI21xp5_ASAP7_75t_L g4862 ( 
.A1(n_4004),
.A2(n_606),
.B(n_605),
.Y(n_4862)
);

O2A1O1Ixp33_ASAP7_75t_L g4863 ( 
.A1(n_4443),
.A2(n_606),
.B(n_607),
.C(n_605),
.Y(n_4863)
);

NAND2xp5_ASAP7_75t_L g4864 ( 
.A(n_4118),
.B(n_606),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4492),
.Y(n_4865)
);

BUFx2_ASAP7_75t_L g4866 ( 
.A(n_4304),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4427),
.Y(n_4867)
);

HB1xp67_ASAP7_75t_L g4868 ( 
.A(n_4393),
.Y(n_4868)
);

AO32x2_ASAP7_75t_L g4869 ( 
.A1(n_4448),
.A2(n_624),
.A3(n_632),
.B1(n_616),
.B2(n_608),
.Y(n_4869)
);

AOI21xp5_ASAP7_75t_L g4870 ( 
.A1(n_4074),
.A2(n_608),
.B(n_607),
.Y(n_4870)
);

BUFx3_ASAP7_75t_L g4871 ( 
.A(n_4304),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4126),
.B(n_609),
.Y(n_4872)
);

NOR2xp33_ASAP7_75t_L g4873 ( 
.A(n_4013),
.B(n_609),
.Y(n_4873)
);

NOR2xp67_ASAP7_75t_L g4874 ( 
.A(n_4296),
.B(n_4403),
.Y(n_4874)
);

AOI21xp5_ASAP7_75t_L g4875 ( 
.A1(n_4039),
.A2(n_610),
.B(n_609),
.Y(n_4875)
);

AND2x2_ASAP7_75t_L g4876 ( 
.A(n_4405),
.B(n_610),
.Y(n_4876)
);

BUFx6f_ASAP7_75t_L g4877 ( 
.A(n_4331),
.Y(n_4877)
);

INVx4_ASAP7_75t_L g4878 ( 
.A(n_4331),
.Y(n_4878)
);

AOI21xp5_ASAP7_75t_L g4879 ( 
.A1(n_4107),
.A2(n_612),
.B(n_611),
.Y(n_4879)
);

BUFx2_ASAP7_75t_L g4880 ( 
.A(n_4051),
.Y(n_4880)
);

CKINVDCx20_ASAP7_75t_R g4881 ( 
.A(n_4347),
.Y(n_4881)
);

NOR2xp33_ASAP7_75t_L g4882 ( 
.A(n_4263),
.B(n_611),
.Y(n_4882)
);

INVx2_ASAP7_75t_L g4883 ( 
.A(n_4454),
.Y(n_4883)
);

AND2x2_ASAP7_75t_L g4884 ( 
.A(n_4197),
.B(n_611),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4435),
.Y(n_4885)
);

OAI22xp5_ASAP7_75t_L g4886 ( 
.A1(n_4395),
.A2(n_4182),
.B1(n_4390),
.B2(n_4381),
.Y(n_4886)
);

A2O1A1Ixp33_ASAP7_75t_L g4887 ( 
.A1(n_4348),
.A2(n_613),
.B(n_614),
.C(n_612),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_SL g4888 ( 
.A(n_4432),
.B(n_612),
.Y(n_4888)
);

BUFx6f_ASAP7_75t_L g4889 ( 
.A(n_4323),
.Y(n_4889)
);

NAND2x1p5_ASAP7_75t_L g4890 ( 
.A(n_3963),
.B(n_613),
.Y(n_4890)
);

BUFx6f_ASAP7_75t_L g4891 ( 
.A(n_4017),
.Y(n_4891)
);

BUFx6f_ASAP7_75t_L g4892 ( 
.A(n_4026),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4132),
.B(n_613),
.Y(n_4893)
);

A2O1A1Ixp33_ASAP7_75t_L g4894 ( 
.A1(n_4419),
.A2(n_615),
.B(n_616),
.C(n_614),
.Y(n_4894)
);

BUFx2_ASAP7_75t_L g4895 ( 
.A(n_4423),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_SL g4896 ( 
.A(n_4438),
.B(n_615),
.Y(n_4896)
);

AOI21xp5_ASAP7_75t_L g4897 ( 
.A1(n_4049),
.A2(n_618),
.B(n_617),
.Y(n_4897)
);

OR2x2_ASAP7_75t_L g4898 ( 
.A(n_4442),
.B(n_617),
.Y(n_4898)
);

INVx3_ASAP7_75t_L g4899 ( 
.A(n_4429),
.Y(n_4899)
);

NOR2xp33_ASAP7_75t_L g4900 ( 
.A(n_4029),
.B(n_617),
.Y(n_4900)
);

AOI21xp5_ASAP7_75t_L g4901 ( 
.A1(n_4133),
.A2(n_619),
.B(n_618),
.Y(n_4901)
);

BUFx6f_ASAP7_75t_L g4902 ( 
.A(n_4066),
.Y(n_4902)
);

AOI21xp5_ASAP7_75t_L g4903 ( 
.A1(n_4034),
.A2(n_619),
.B(n_618),
.Y(n_4903)
);

OAI21xp33_ASAP7_75t_L g4904 ( 
.A1(n_4472),
.A2(n_621),
.B(n_620),
.Y(n_4904)
);

BUFx3_ASAP7_75t_L g4905 ( 
.A(n_4336),
.Y(n_4905)
);

INVxp67_ASAP7_75t_L g4906 ( 
.A(n_4083),
.Y(n_4906)
);

AOI21xp5_ASAP7_75t_L g4907 ( 
.A1(n_4280),
.A2(n_621),
.B(n_620),
.Y(n_4907)
);

CKINVDCx5p33_ASAP7_75t_R g4908 ( 
.A(n_4353),
.Y(n_4908)
);

O2A1O1Ixp33_ASAP7_75t_SL g4909 ( 
.A1(n_4300),
.A2(n_622),
.B(n_623),
.C(n_621),
.Y(n_4909)
);

INVx2_ASAP7_75t_L g4910 ( 
.A(n_4477),
.Y(n_4910)
);

HB1xp67_ASAP7_75t_L g4911 ( 
.A(n_4458),
.Y(n_4911)
);

AOI22xp5_ASAP7_75t_L g4912 ( 
.A1(n_4015),
.A2(n_1068),
.B1(n_1071),
.B2(n_1067),
.Y(n_4912)
);

HB1xp67_ASAP7_75t_L g4913 ( 
.A(n_4401),
.Y(n_4913)
);

O2A1O1Ixp33_ASAP7_75t_L g4914 ( 
.A1(n_4247),
.A2(n_623),
.B(n_624),
.C(n_622),
.Y(n_4914)
);

NAND2xp5_ASAP7_75t_SL g4915 ( 
.A(n_4441),
.B(n_622),
.Y(n_4915)
);

O2A1O1Ixp33_ASAP7_75t_L g4916 ( 
.A1(n_4355),
.A2(n_625),
.B(n_626),
.C(n_624),
.Y(n_4916)
);

NOR2xp33_ASAP7_75t_L g4917 ( 
.A(n_4048),
.B(n_625),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4444),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4445),
.Y(n_4919)
);

AOI21xp5_ASAP7_75t_L g4920 ( 
.A1(n_4024),
.A2(n_626),
.B(n_625),
.Y(n_4920)
);

CKINVDCx14_ASAP7_75t_R g4921 ( 
.A(n_4245),
.Y(n_4921)
);

NOR2xp33_ASAP7_75t_L g4922 ( 
.A(n_4422),
.B(n_626),
.Y(n_4922)
);

BUFx2_ASAP7_75t_L g4923 ( 
.A(n_4456),
.Y(n_4923)
);

OAI22xp5_ASAP7_75t_SL g4924 ( 
.A1(n_4466),
.A2(n_4394),
.B1(n_4170),
.B2(n_4159),
.Y(n_4924)
);

AOI21xp5_ASAP7_75t_L g4925 ( 
.A1(n_4464),
.A2(n_628),
.B(n_627),
.Y(n_4925)
);

BUFx3_ASAP7_75t_L g4926 ( 
.A(n_4399),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4137),
.Y(n_4927)
);

A2O1A1Ixp33_ASAP7_75t_L g4928 ( 
.A1(n_4096),
.A2(n_628),
.B(n_629),
.C(n_627),
.Y(n_4928)
);

A2O1A1Ixp33_ASAP7_75t_SL g4929 ( 
.A1(n_4416),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_4929)
);

AOI21x1_ASAP7_75t_L g4930 ( 
.A1(n_4484),
.A2(n_4468),
.B(n_4467),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4139),
.Y(n_4931)
);

AOI21xp5_ASAP7_75t_L g4932 ( 
.A1(n_4475),
.A2(n_630),
.B(n_629),
.Y(n_4932)
);

NAND2x1_ASAP7_75t_SL g4933 ( 
.A(n_4214),
.B(n_1054),
.Y(n_4933)
);

AND2x2_ASAP7_75t_L g4934 ( 
.A(n_4351),
.B(n_629),
.Y(n_4934)
);

INVx1_ASAP7_75t_SL g4935 ( 
.A(n_4396),
.Y(n_4935)
);

AO21x2_ASAP7_75t_L g4936 ( 
.A1(n_4451),
.A2(n_631),
.B(n_630),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_4156),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_4478),
.A2(n_631),
.B(n_630),
.Y(n_4938)
);

OAI22xp33_ASAP7_75t_L g4939 ( 
.A1(n_4316),
.A2(n_633),
.B1(n_634),
.B2(n_632),
.Y(n_4939)
);

BUFx6f_ASAP7_75t_SL g4940 ( 
.A(n_4410),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_SL g4941 ( 
.A(n_4350),
.B(n_633),
.Y(n_4941)
);

OAI21xp5_ASAP7_75t_L g4942 ( 
.A1(n_4264),
.A2(n_634),
.B(n_633),
.Y(n_4942)
);

A2O1A1Ixp33_ASAP7_75t_L g4943 ( 
.A1(n_4409),
.A2(n_635),
.B(n_636),
.C(n_634),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4158),
.B(n_635),
.Y(n_4944)
);

O2A1O1Ixp33_ASAP7_75t_L g4945 ( 
.A1(n_4481),
.A2(n_636),
.B(n_637),
.C(n_635),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_L g4946 ( 
.A(n_4163),
.B(n_636),
.Y(n_4946)
);

BUFx3_ASAP7_75t_L g4947 ( 
.A(n_4082),
.Y(n_4947)
);

NOR2xp33_ASAP7_75t_L g4948 ( 
.A(n_4365),
.B(n_637),
.Y(n_4948)
);

INVx2_ASAP7_75t_L g4949 ( 
.A(n_4329),
.Y(n_4949)
);

AOI21xp5_ASAP7_75t_L g4950 ( 
.A1(n_4479),
.A2(n_4482),
.B(n_4480),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4643),
.B(n_4177),
.Y(n_4951)
);

INVx2_ASAP7_75t_L g4952 ( 
.A(n_4689),
.Y(n_4952)
);

AO31x2_ASAP7_75t_L g4953 ( 
.A1(n_4806),
.A2(n_4111),
.A3(n_4496),
.B(n_4488),
.Y(n_4953)
);

NAND3xp33_ASAP7_75t_L g4954 ( 
.A(n_4595),
.B(n_4203),
.C(n_4461),
.Y(n_4954)
);

AO32x2_ASAP7_75t_L g4955 ( 
.A1(n_4753),
.A2(n_4240),
.A3(n_4354),
.B1(n_4058),
.B2(n_4500),
.Y(n_4955)
);

NAND3x1_ASAP7_75t_L g4956 ( 
.A(n_4528),
.B(n_4255),
.C(n_4130),
.Y(n_4956)
);

OAI21x1_ASAP7_75t_L g4957 ( 
.A1(n_4553),
.A2(n_4178),
.B(n_4067),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_SL g4958 ( 
.A(n_4682),
.B(n_4292),
.Y(n_4958)
);

NOR4xp25_ASAP7_75t_L g4959 ( 
.A(n_4545),
.B(n_4187),
.C(n_4330),
.D(n_4317),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_SL g4960 ( 
.A(n_4682),
.B(n_4266),
.Y(n_4960)
);

AOI21xp5_ASAP7_75t_L g4961 ( 
.A1(n_4502),
.A2(n_4299),
.B(n_4302),
.Y(n_4961)
);

A2O1A1Ixp33_ASAP7_75t_L g4962 ( 
.A1(n_4508),
.A2(n_4512),
.B(n_4548),
.C(n_4607),
.Y(n_4962)
);

BUFx6f_ASAP7_75t_L g4963 ( 
.A(n_4576),
.Y(n_4963)
);

NAND2xp5_ASAP7_75t_L g4964 ( 
.A(n_4657),
.B(n_4184),
.Y(n_4964)
);

AOI21xp5_ASAP7_75t_L g4965 ( 
.A1(n_4554),
.A2(n_4090),
.B(n_4112),
.Y(n_4965)
);

NAND2x1p5_ASAP7_75t_L g4966 ( 
.A(n_4521),
.B(n_4633),
.Y(n_4966)
);

BUFx2_ASAP7_75t_L g4967 ( 
.A(n_4562),
.Y(n_4967)
);

INVx3_ASAP7_75t_L g4968 ( 
.A(n_4708),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4667),
.Y(n_4969)
);

OAI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4560),
.A2(n_4609),
.B(n_4734),
.Y(n_4970)
);

AO32x2_ASAP7_75t_L g4971 ( 
.A1(n_4564),
.A2(n_4616),
.A3(n_4886),
.B1(n_4924),
.B2(n_4858),
.Y(n_4971)
);

O2A1O1Ixp5_ASAP7_75t_L g4972 ( 
.A1(n_4511),
.A2(n_4224),
.B(n_4226),
.C(n_4223),
.Y(n_4972)
);

OR2x2_ASAP7_75t_L g4973 ( 
.A(n_4536),
.B(n_4339),
.Y(n_4973)
);

AO31x2_ASAP7_75t_L g4974 ( 
.A1(n_4883),
.A2(n_4169),
.A3(n_4209),
.B(n_4122),
.Y(n_4974)
);

INVx3_ASAP7_75t_L g4975 ( 
.A(n_4814),
.Y(n_4975)
);

O2A1O1Ixp5_ASAP7_75t_L g4976 ( 
.A1(n_4515),
.A2(n_4228),
.B(n_4229),
.C(n_4227),
.Y(n_4976)
);

INVx2_ASAP7_75t_L g4977 ( 
.A(n_4690),
.Y(n_4977)
);

BUFx3_ASAP7_75t_L g4978 ( 
.A(n_4736),
.Y(n_4978)
);

NAND3xp33_ASAP7_75t_L g4979 ( 
.A(n_4602),
.B(n_4234),
.C(n_4232),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4723),
.B(n_4190),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4532),
.Y(n_4981)
);

AOI22xp33_ASAP7_75t_L g4982 ( 
.A1(n_4516),
.A2(n_4387),
.B1(n_4411),
.B2(n_4414),
.Y(n_4982)
);

AND2x6_ASAP7_75t_L g4983 ( 
.A(n_4700),
.B(n_4033),
.Y(n_4983)
);

AO32x2_ASAP7_75t_L g4984 ( 
.A1(n_4556),
.A2(n_4404),
.A3(n_4345),
.B1(n_4366),
.B2(n_4211),
.Y(n_4984)
);

INVx2_ASAP7_75t_SL g4985 ( 
.A(n_4727),
.Y(n_4985)
);

NAND2x1_ASAP7_75t_L g4986 ( 
.A(n_4860),
.B(n_4195),
.Y(n_4986)
);

AOI21xp5_ASAP7_75t_L g4987 ( 
.A1(n_4732),
.A2(n_4119),
.B(n_4253),
.Y(n_4987)
);

OA21x2_ASAP7_75t_L g4988 ( 
.A1(n_4649),
.A2(n_4222),
.B(n_4201),
.Y(n_4988)
);

AOI31xp67_ASAP7_75t_L g4989 ( 
.A1(n_4910),
.A2(n_4949),
.A3(n_4837),
.B(n_4803),
.Y(n_4989)
);

O2A1O1Ixp33_ASAP7_75t_L g4990 ( 
.A1(n_4617),
.A2(n_3969),
.B(n_4241),
.C(n_4230),
.Y(n_4990)
);

NAND2xp5_ASAP7_75t_L g4991 ( 
.A(n_4504),
.B(n_4262),
.Y(n_4991)
);

AOI21xp5_ASAP7_75t_L g4992 ( 
.A1(n_4619),
.A2(n_4276),
.B(n_4152),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4711),
.B(n_4270),
.Y(n_4993)
);

AOI221x1_ASAP7_75t_L g4994 ( 
.A1(n_4542),
.A2(n_4830),
.B1(n_4570),
.B2(n_4603),
.C(n_4904),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4506),
.B(n_4272),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4811),
.B(n_4819),
.Y(n_4996)
);

BUFx2_ASAP7_75t_L g4997 ( 
.A(n_4576),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4825),
.B(n_4277),
.Y(n_4998)
);

OA21x2_ASAP7_75t_L g4999 ( 
.A1(n_4509),
.A2(n_4289),
.B(n_4176),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_L g5000 ( 
.A(n_4507),
.B(n_4054),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_SL g5001 ( 
.A(n_4682),
.B(n_4326),
.Y(n_5001)
);

NOR3xp33_ASAP7_75t_L g5002 ( 
.A(n_4592),
.B(n_4056),
.C(n_4384),
.Y(n_5002)
);

NOR2xp33_ASAP7_75t_SL g5003 ( 
.A(n_4828),
.B(n_4239),
.Y(n_5003)
);

AO31x2_ASAP7_75t_L g5004 ( 
.A1(n_4793),
.A2(n_4179),
.A3(n_4183),
.B(n_4174),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_SL g5005 ( 
.A(n_4706),
.B(n_4243),
.Y(n_5005)
);

AOI21xp5_ASAP7_75t_L g5006 ( 
.A1(n_4706),
.A2(n_4154),
.B(n_4150),
.Y(n_5006)
);

BUFx2_ASAP7_75t_L g5007 ( 
.A(n_4576),
.Y(n_5007)
);

O2A1O1Ixp33_ASAP7_75t_SL g5008 ( 
.A1(n_4524),
.A2(n_4161),
.B(n_4344),
.C(n_4342),
.Y(n_5008)
);

OAI21x1_ASAP7_75t_L g5009 ( 
.A1(n_4930),
.A2(n_4186),
.B(n_4185),
.Y(n_5009)
);

OAI21x1_ASAP7_75t_L g5010 ( 
.A1(n_4770),
.A2(n_4666),
.B(n_4714),
.Y(n_5010)
);

NOR2xp67_ASAP7_75t_L g5011 ( 
.A(n_4706),
.B(n_640),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_L g5012 ( 
.A(n_4514),
.B(n_4530),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4540),
.Y(n_5013)
);

OAI21x1_ASAP7_75t_L g5014 ( 
.A1(n_4680),
.A2(n_4204),
.B(n_4193),
.Y(n_5014)
);

OAI22x1_ASAP7_75t_L g5015 ( 
.A1(n_4678),
.A2(n_4059),
.B1(n_4050),
.B2(n_638),
.Y(n_5015)
);

NOR3xp33_ASAP7_75t_SL g5016 ( 
.A(n_4529),
.B(n_4363),
.C(n_4360),
.Y(n_5016)
);

AO31x2_ASAP7_75t_L g5017 ( 
.A1(n_4597),
.A2(n_4221),
.A3(n_4219),
.B(n_4283),
.Y(n_5017)
);

OAI21x1_ASAP7_75t_L g5018 ( 
.A1(n_4709),
.A2(n_4286),
.B(n_4284),
.Y(n_5018)
);

A2O1A1Ixp33_ASAP7_75t_L g5019 ( 
.A1(n_4672),
.A2(n_4374),
.B(n_4287),
.C(n_4310),
.Y(n_5019)
);

OAI21x1_ASAP7_75t_L g5020 ( 
.A1(n_4539),
.A2(n_4311),
.B(n_4288),
.Y(n_5020)
);

OAI21x1_ASAP7_75t_L g5021 ( 
.A1(n_4647),
.A2(n_4319),
.B(n_4314),
.Y(n_5021)
);

AOI21xp5_ASAP7_75t_L g5022 ( 
.A1(n_4737),
.A2(n_4321),
.B(n_4320),
.Y(n_5022)
);

AOI21xp5_ASAP7_75t_L g5023 ( 
.A1(n_4737),
.A2(n_4064),
.B(n_4025),
.Y(n_5023)
);

AND3x4_ASAP7_75t_L g5024 ( 
.A(n_4676),
.B(n_638),
.C(n_637),
.Y(n_5024)
);

BUFx3_ASAP7_75t_L g5025 ( 
.A(n_4685),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4549),
.Y(n_5026)
);

OA21x2_ASAP7_75t_L g5027 ( 
.A1(n_4867),
.A2(n_4918),
.B(n_4885),
.Y(n_5027)
);

AO31x2_ASAP7_75t_L g5028 ( 
.A1(n_4923),
.A2(n_640),
.A3(n_641),
.B(n_639),
.Y(n_5028)
);

AOI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_4737),
.A2(n_640),
.B(n_639),
.Y(n_5029)
);

NOR4xp25_ASAP7_75t_L g5030 ( 
.A(n_4935),
.B(n_642),
.C(n_643),
.D(n_641),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_SL g5031 ( 
.A(n_4537),
.B(n_641),
.Y(n_5031)
);

OR2x2_ASAP7_75t_L g5032 ( 
.A(n_4817),
.B(n_642),
.Y(n_5032)
);

NOR2xp67_ASAP7_75t_SL g5033 ( 
.A(n_4675),
.B(n_643),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_SL g5034 ( 
.A(n_4820),
.B(n_644),
.Y(n_5034)
);

OA22x2_ASAP7_75t_L g5035 ( 
.A1(n_4516),
.A2(n_645),
.B1(n_646),
.B2(n_644),
.Y(n_5035)
);

NAND3xp33_ASAP7_75t_L g5036 ( 
.A(n_4505),
.B(n_646),
.C(n_644),
.Y(n_5036)
);

NOR2xp67_ASAP7_75t_SL g5037 ( 
.A(n_4745),
.B(n_646),
.Y(n_5037)
);

BUFx3_ASAP7_75t_L g5038 ( 
.A(n_4645),
.Y(n_5038)
);

OAI21xp5_ASAP7_75t_L g5039 ( 
.A1(n_4687),
.A2(n_648),
.B(n_647),
.Y(n_5039)
);

OR2x2_ASAP7_75t_L g5040 ( 
.A(n_4552),
.B(n_4561),
.Y(n_5040)
);

OAI21xp5_ASAP7_75t_SL g5041 ( 
.A1(n_4890),
.A2(n_648),
.B(n_647),
.Y(n_5041)
);

CKINVDCx20_ASAP7_75t_R g5042 ( 
.A(n_4557),
.Y(n_5042)
);

AND3x4_ASAP7_75t_L g5043 ( 
.A(n_4763),
.B(n_649),
.C(n_647),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_4563),
.B(n_649),
.Y(n_5044)
);

OAI21x1_ASAP7_75t_SL g5045 ( 
.A1(n_4852),
.A2(n_651),
.B(n_650),
.Y(n_5045)
);

A2O1A1Ixp33_ASAP7_75t_L g5046 ( 
.A1(n_4547),
.A2(n_651),
.B(n_652),
.C(n_650),
.Y(n_5046)
);

BUFx12f_ASAP7_75t_L g5047 ( 
.A(n_4679),
.Y(n_5047)
);

O2A1O1Ixp5_ASAP7_75t_L g5048 ( 
.A1(n_4652),
.A2(n_653),
.B(n_654),
.C(n_651),
.Y(n_5048)
);

O2A1O1Ixp33_ASAP7_75t_SL g5049 ( 
.A1(n_4551),
.A2(n_654),
.B(n_655),
.C(n_653),
.Y(n_5049)
);

INVxp67_ASAP7_75t_SL g5050 ( 
.A(n_4832),
.Y(n_5050)
);

AND2x2_ASAP7_75t_L g5051 ( 
.A(n_4892),
.B(n_14),
.Y(n_5051)
);

BUFx12f_ASAP7_75t_L g5052 ( 
.A(n_4713),
.Y(n_5052)
);

INVx5_ASAP7_75t_L g5053 ( 
.A(n_4550),
.Y(n_5053)
);

BUFx2_ASAP7_75t_L g5054 ( 
.A(n_4638),
.Y(n_5054)
);

INVx2_ASAP7_75t_SL g5055 ( 
.A(n_4758),
.Y(n_5055)
);

AO31x2_ASAP7_75t_L g5056 ( 
.A1(n_4919),
.A2(n_654),
.A3(n_655),
.B(n_653),
.Y(n_5056)
);

NAND3xp33_ASAP7_75t_L g5057 ( 
.A(n_4842),
.B(n_656),
.C(n_655),
.Y(n_5057)
);

AOI21x1_ASAP7_75t_L g5058 ( 
.A1(n_4661),
.A2(n_657),
.B(n_656),
.Y(n_5058)
);

OAI21xp5_ASAP7_75t_L g5059 ( 
.A1(n_4757),
.A2(n_657),
.B(n_656),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_4580),
.Y(n_5060)
);

INVx2_ASAP7_75t_L g5061 ( 
.A(n_4538),
.Y(n_5061)
);

A2O1A1Ixp33_ASAP7_75t_L g5062 ( 
.A1(n_4764),
.A2(n_658),
.B(n_659),
.C(n_657),
.Y(n_5062)
);

BUFx3_ASAP7_75t_L g5063 ( 
.A(n_4696),
.Y(n_5063)
);

AOI21x1_ASAP7_75t_L g5064 ( 
.A1(n_4681),
.A2(n_4598),
.B(n_4821),
.Y(n_5064)
);

OAI21x1_ASAP7_75t_L g5065 ( 
.A1(n_4950),
.A2(n_4749),
.B(n_4740),
.Y(n_5065)
);

OAI21x1_ASAP7_75t_L g5066 ( 
.A1(n_4768),
.A2(n_659),
.B(n_658),
.Y(n_5066)
);

CKINVDCx5p33_ASAP7_75t_R g5067 ( 
.A(n_4705),
.Y(n_5067)
);

INVxp33_ASAP7_75t_L g5068 ( 
.A(n_4748),
.Y(n_5068)
);

OAI21x1_ASAP7_75t_L g5069 ( 
.A1(n_4783),
.A2(n_659),
.B(n_658),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_4584),
.B(n_660),
.Y(n_5070)
);

AOI21xp5_ASAP7_75t_L g5071 ( 
.A1(n_4717),
.A2(n_4813),
.B(n_4683),
.Y(n_5071)
);

OAI21x1_ASAP7_75t_L g5072 ( 
.A1(n_4527),
.A2(n_661),
.B(n_660),
.Y(n_5072)
);

NOR2xp33_ASAP7_75t_SL g5073 ( 
.A(n_4624),
.B(n_660),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4588),
.Y(n_5074)
);

O2A1O1Ixp33_ASAP7_75t_L g5075 ( 
.A1(n_4627),
.A2(n_662),
.B(n_663),
.C(n_661),
.Y(n_5075)
);

INVxp67_ASAP7_75t_SL g5076 ( 
.A(n_4669),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_4625),
.B(n_662),
.Y(n_5077)
);

A2O1A1Ixp33_ASAP7_75t_L g5078 ( 
.A1(n_4733),
.A2(n_665),
.B(n_666),
.C(n_664),
.Y(n_5078)
);

O2A1O1Ixp33_ASAP7_75t_L g5079 ( 
.A1(n_4650),
.A2(n_4847),
.B(n_4845),
.C(n_4929),
.Y(n_5079)
);

INVx2_ASAP7_75t_L g5080 ( 
.A(n_4544),
.Y(n_5080)
);

OAI21x1_ASAP7_75t_L g5081 ( 
.A1(n_4535),
.A2(n_665),
.B(n_664),
.Y(n_5081)
);

INVx2_ASAP7_75t_SL g5082 ( 
.A(n_4639),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_4590),
.Y(n_5083)
);

OA21x2_ASAP7_75t_L g5084 ( 
.A1(n_4776),
.A2(n_665),
.B(n_664),
.Y(n_5084)
);

NAND3xp33_ASAP7_75t_L g5085 ( 
.A(n_4843),
.B(n_667),
.C(n_666),
.Y(n_5085)
);

AOI21xp5_ASAP7_75t_L g5086 ( 
.A1(n_4941),
.A2(n_4840),
.B(n_4747),
.Y(n_5086)
);

AOI21xp5_ASAP7_75t_L g5087 ( 
.A1(n_4862),
.A2(n_667),
.B(n_666),
.Y(n_5087)
);

A2O1A1Ixp33_ASAP7_75t_L g5088 ( 
.A1(n_4914),
.A2(n_668),
.B(n_669),
.C(n_667),
.Y(n_5088)
);

OR2x2_ASAP7_75t_L g5089 ( 
.A(n_4660),
.B(n_668),
.Y(n_5089)
);

AOI21xp5_ASAP7_75t_L g5090 ( 
.A1(n_4707),
.A2(n_670),
.B(n_668),
.Y(n_5090)
);

O2A1O1Ixp33_ASAP7_75t_L g5091 ( 
.A1(n_4788),
.A2(n_671),
.B(n_672),
.C(n_670),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4715),
.B(n_670),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4618),
.Y(n_5093)
);

OAI21x1_ASAP7_75t_L g5094 ( 
.A1(n_4720),
.A2(n_4899),
.B(n_4543),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_L g5095 ( 
.A(n_4722),
.B(n_671),
.Y(n_5095)
);

AOI31xp67_ASAP7_75t_L g5096 ( 
.A1(n_4851),
.A2(n_672),
.A3(n_673),
.B(n_671),
.Y(n_5096)
);

AOI21x1_ASAP7_75t_L g5097 ( 
.A1(n_4874),
.A2(n_674),
.B(n_673),
.Y(n_5097)
);

AOI21xp5_ASAP7_75t_L g5098 ( 
.A1(n_4826),
.A2(n_675),
.B(n_674),
.Y(n_5098)
);

NAND2xp5_ASAP7_75t_L g5099 ( 
.A(n_4927),
.B(n_675),
.Y(n_5099)
);

BUFx6f_ASAP7_75t_L g5100 ( 
.A(n_4638),
.Y(n_5100)
);

AND3x2_ASAP7_75t_L g5101 ( 
.A(n_4704),
.B(n_4517),
.C(n_4510),
.Y(n_5101)
);

BUFx12f_ASAP7_75t_L g5102 ( 
.A(n_4801),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_4555),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_SL g5104 ( 
.A(n_4820),
.B(n_676),
.Y(n_5104)
);

AO31x2_ASAP7_75t_L g5105 ( 
.A1(n_4730),
.A2(n_4807),
.A3(n_4895),
.B(n_4854),
.Y(n_5105)
);

OAI22xp5_ASAP7_75t_L g5106 ( 
.A1(n_4769),
.A2(n_678),
.B1(n_679),
.B2(n_677),
.Y(n_5106)
);

OAI21x1_ASAP7_75t_L g5107 ( 
.A1(n_4568),
.A2(n_678),
.B(n_677),
.Y(n_5107)
);

OAI21x1_ASAP7_75t_L g5108 ( 
.A1(n_4569),
.A2(n_679),
.B(n_678),
.Y(n_5108)
);

NAND2xp5_ASAP7_75t_SL g5109 ( 
.A(n_4820),
.B(n_680),
.Y(n_5109)
);

AOI221x1_ASAP7_75t_L g5110 ( 
.A1(n_4578),
.A2(n_4574),
.B1(n_4653),
.B2(n_4692),
.C(n_4774),
.Y(n_5110)
);

A2O1A1Ixp33_ASAP7_75t_L g5111 ( 
.A1(n_4626),
.A2(n_681),
.B(n_682),
.C(n_680),
.Y(n_5111)
);

NOR2xp67_ASAP7_75t_L g5112 ( 
.A(n_4566),
.B(n_685),
.Y(n_5112)
);

OAI21x1_ASAP7_75t_L g5113 ( 
.A1(n_4589),
.A2(n_682),
.B(n_681),
.Y(n_5113)
);

OAI21xp5_ASAP7_75t_L g5114 ( 
.A1(n_4605),
.A2(n_682),
.B(n_681),
.Y(n_5114)
);

AOI21xp5_ASAP7_75t_L g5115 ( 
.A1(n_4596),
.A2(n_684),
.B(n_683),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4558),
.Y(n_5116)
);

AOI21xp33_ASAP7_75t_L g5117 ( 
.A1(n_4526),
.A2(n_684),
.B(n_683),
.Y(n_5117)
);

AND2x6_ASAP7_75t_L g5118 ( 
.A(n_4525),
.B(n_684),
.Y(n_5118)
);

INVxp67_ASAP7_75t_L g5119 ( 
.A(n_4947),
.Y(n_5119)
);

OAI21x1_ASAP7_75t_L g5120 ( 
.A1(n_4594),
.A2(n_686),
.B(n_685),
.Y(n_5120)
);

AOI21xp5_ASAP7_75t_L g5121 ( 
.A1(n_4565),
.A2(n_686),
.B(n_685),
.Y(n_5121)
);

AOI21xp5_ASAP7_75t_L g5122 ( 
.A1(n_4519),
.A2(n_687),
.B(n_686),
.Y(n_5122)
);

AOI21xp5_ASAP7_75t_L g5123 ( 
.A1(n_4534),
.A2(n_688),
.B(n_687),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_4567),
.Y(n_5124)
);

NAND2xp5_ASAP7_75t_L g5125 ( 
.A(n_4931),
.B(n_687),
.Y(n_5125)
);

OAI21x1_ASAP7_75t_L g5126 ( 
.A1(n_4800),
.A2(n_689),
.B(n_688),
.Y(n_5126)
);

OAI21x1_ASAP7_75t_L g5127 ( 
.A1(n_4741),
.A2(n_690),
.B(n_689),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_4581),
.Y(n_5128)
);

INVxp67_ASAP7_75t_SL g5129 ( 
.A(n_4834),
.Y(n_5129)
);

OAI21x1_ASAP7_75t_L g5130 ( 
.A1(n_4664),
.A2(n_690),
.B(n_689),
.Y(n_5130)
);

NOR2xp33_ASAP7_75t_L g5131 ( 
.A(n_4921),
.B(n_15),
.Y(n_5131)
);

BUFx3_ASAP7_75t_L g5132 ( 
.A(n_4600),
.Y(n_5132)
);

AOI211x1_ASAP7_75t_L g5133 ( 
.A1(n_4739),
.A2(n_691),
.B(n_692),
.C(n_690),
.Y(n_5133)
);

AND2x4_ASAP7_75t_L g5134 ( 
.A(n_4835),
.B(n_691),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_4937),
.B(n_691),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_4629),
.Y(n_5136)
);

NAND2xp5_ASAP7_75t_L g5137 ( 
.A(n_4782),
.B(n_692),
.Y(n_5137)
);

NAND2xp5_ASAP7_75t_L g5138 ( 
.A(n_4892),
.B(n_692),
.Y(n_5138)
);

NAND2x1_ASAP7_75t_L g5139 ( 
.A(n_4525),
.B(n_693),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_4659),
.Y(n_5140)
);

NAND2xp5_ASAP7_75t_L g5141 ( 
.A(n_4853),
.B(n_693),
.Y(n_5141)
);

OR2x2_ASAP7_75t_L g5142 ( 
.A(n_4865),
.B(n_693),
.Y(n_5142)
);

INVx2_ASAP7_75t_L g5143 ( 
.A(n_4638),
.Y(n_5143)
);

AOI21xp5_ASAP7_75t_L g5144 ( 
.A1(n_4861),
.A2(n_695),
.B(n_694),
.Y(n_5144)
);

AO31x2_ASAP7_75t_L g5145 ( 
.A1(n_4634),
.A2(n_4631),
.A3(n_4637),
.B(n_4750),
.Y(n_5145)
);

NAND2xp5_ASAP7_75t_SL g5146 ( 
.A(n_4790),
.B(n_695),
.Y(n_5146)
);

AO22x2_ASAP7_75t_L g5147 ( 
.A1(n_4752),
.A2(n_696),
.B1(n_697),
.B2(n_695),
.Y(n_5147)
);

BUFx2_ASAP7_75t_L g5148 ( 
.A(n_4503),
.Y(n_5148)
);

NAND2x1p5_ASAP7_75t_L g5149 ( 
.A(n_4878),
.B(n_696),
.Y(n_5149)
);

BUFx2_ASAP7_75t_SL g5150 ( 
.A(n_4754),
.Y(n_5150)
);

INVx2_ASAP7_75t_L g5151 ( 
.A(n_4673),
.Y(n_5151)
);

AOI21xp5_ASAP7_75t_L g5152 ( 
.A1(n_4888),
.A2(n_698),
.B(n_697),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_4772),
.B(n_697),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_4868),
.Y(n_5154)
);

AOI21x1_ASAP7_75t_L g5155 ( 
.A1(n_4841),
.A2(n_699),
.B(n_698),
.Y(n_5155)
);

AOI21xp5_ASAP7_75t_L g5156 ( 
.A1(n_4896),
.A2(n_700),
.B(n_698),
.Y(n_5156)
);

OAI21x1_ASAP7_75t_L g5157 ( 
.A1(n_4671),
.A2(n_701),
.B(n_700),
.Y(n_5157)
);

A2O1A1Ixp33_ASAP7_75t_L g5158 ( 
.A1(n_4518),
.A2(n_702),
.B(n_703),
.C(n_701),
.Y(n_5158)
);

OAI21x1_ASAP7_75t_L g5159 ( 
.A1(n_4933),
.A2(n_703),
.B(n_702),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4911),
.Y(n_5160)
);

AND2x2_ASAP7_75t_L g5161 ( 
.A(n_4522),
.B(n_15),
.Y(n_5161)
);

O2A1O1Ixp33_ASAP7_75t_L g5162 ( 
.A1(n_4523),
.A2(n_704),
.B(n_705),
.C(n_702),
.Y(n_5162)
);

INVx1_ASAP7_75t_SL g5163 ( 
.A(n_4608),
.Y(n_5163)
);

OAI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_4897),
.A2(n_705),
.B(n_704),
.Y(n_5164)
);

NOR2x1_ASAP7_75t_SL g5165 ( 
.A(n_4761),
.B(n_704),
.Y(n_5165)
);

OAI21x1_ASAP7_75t_L g5166 ( 
.A1(n_4620),
.A2(n_707),
.B(n_706),
.Y(n_5166)
);

OAI21xp5_ASAP7_75t_L g5167 ( 
.A1(n_4599),
.A2(n_707),
.B(n_706),
.Y(n_5167)
);

AOI21xp5_ASAP7_75t_L g5168 ( 
.A1(n_4915),
.A2(n_709),
.B(n_708),
.Y(n_5168)
);

OAI21x1_ASAP7_75t_L g5169 ( 
.A1(n_4674),
.A2(n_709),
.B(n_708),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_4913),
.B(n_708),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_4789),
.B(n_709),
.Y(n_5171)
);

AND2x2_ASAP7_75t_L g5172 ( 
.A(n_4591),
.B(n_4628),
.Y(n_5172)
);

O2A1O1Ixp33_ASAP7_75t_SL g5173 ( 
.A1(n_4894),
.A2(n_711),
.B(n_712),
.C(n_710),
.Y(n_5173)
);

INVx2_ASAP7_75t_L g5174 ( 
.A(n_4673),
.Y(n_5174)
);

INVx2_ASAP7_75t_L g5175 ( 
.A(n_4673),
.Y(n_5175)
);

INVx2_ASAP7_75t_L g5176 ( 
.A(n_4703),
.Y(n_5176)
);

OA21x2_ASAP7_75t_L g5177 ( 
.A1(n_4839),
.A2(n_711),
.B(n_710),
.Y(n_5177)
);

INVx5_ASAP7_75t_L g5178 ( 
.A(n_4662),
.Y(n_5178)
);

OAI21x1_ASAP7_75t_L g5179 ( 
.A1(n_4684),
.A2(n_711),
.B(n_710),
.Y(n_5179)
);

INVx2_ASAP7_75t_SL g5180 ( 
.A(n_4503),
.Y(n_5180)
);

NOR4xp25_ASAP7_75t_L g5181 ( 
.A(n_4668),
.B(n_714),
.C(n_715),
.D(n_712),
.Y(n_5181)
);

INVx2_ASAP7_75t_L g5182 ( 
.A(n_4703),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_4856),
.Y(n_5183)
);

CKINVDCx5p33_ASAP7_75t_R g5184 ( 
.A(n_4810),
.Y(n_5184)
);

AOI21x1_ASAP7_75t_L g5185 ( 
.A1(n_4604),
.A2(n_716),
.B(n_714),
.Y(n_5185)
);

NOR2x1_ASAP7_75t_SL g5186 ( 
.A(n_4765),
.B(n_714),
.Y(n_5186)
);

AO31x2_ASAP7_75t_L g5187 ( 
.A1(n_4760),
.A2(n_717),
.A3(n_718),
.B(n_716),
.Y(n_5187)
);

AO21x2_ASAP7_75t_L g5188 ( 
.A1(n_4698),
.A2(n_718),
.B(n_717),
.Y(n_5188)
);

AOI21xp5_ASAP7_75t_L g5189 ( 
.A1(n_4838),
.A2(n_720),
.B(n_719),
.Y(n_5189)
);

AND2x2_ASAP7_75t_L g5190 ( 
.A(n_4716),
.B(n_16),
.Y(n_5190)
);

INVx4_ASAP7_75t_SL g5191 ( 
.A(n_4773),
.Y(n_5191)
);

AO21x1_ASAP7_75t_L g5192 ( 
.A1(n_4752),
.A2(n_720),
.B(n_719),
.Y(n_5192)
);

NAND2xp5_ASAP7_75t_L g5193 ( 
.A(n_4859),
.B(n_719),
.Y(n_5193)
);

AND2x2_ASAP7_75t_L g5194 ( 
.A(n_4632),
.B(n_16),
.Y(n_5194)
);

OAI21xp5_ASAP7_75t_L g5195 ( 
.A1(n_4577),
.A2(n_721),
.B(n_720),
.Y(n_5195)
);

OAI21x1_ASAP7_75t_L g5196 ( 
.A1(n_4829),
.A2(n_722),
.B(n_721),
.Y(n_5196)
);

AND2x2_ASAP7_75t_L g5197 ( 
.A(n_4663),
.B(n_16),
.Y(n_5197)
);

O2A1O1Ixp33_ASAP7_75t_SL g5198 ( 
.A1(n_4779),
.A2(n_723),
.B(n_724),
.C(n_722),
.Y(n_5198)
);

OAI21xp5_ASAP7_75t_L g5199 ( 
.A1(n_4582),
.A2(n_724),
.B(n_723),
.Y(n_5199)
);

OAI21x1_ASAP7_75t_L g5200 ( 
.A1(n_4875),
.A2(n_724),
.B(n_723),
.Y(n_5200)
);

NAND2xp5_ASAP7_75t_L g5201 ( 
.A(n_4859),
.B(n_4898),
.Y(n_5201)
);

OAI21xp5_ASAP7_75t_L g5202 ( 
.A1(n_4738),
.A2(n_726),
.B(n_725),
.Y(n_5202)
);

AO21x2_ASAP7_75t_L g5203 ( 
.A1(n_4701),
.A2(n_726),
.B(n_725),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_L g5204 ( 
.A(n_4762),
.B(n_4697),
.Y(n_5204)
);

OAI21x1_ASAP7_75t_L g5205 ( 
.A1(n_4798),
.A2(n_727),
.B(n_726),
.Y(n_5205)
);

NAND2xp5_ASAP7_75t_L g5206 ( 
.A(n_4777),
.B(n_1074),
.Y(n_5206)
);

AOI21xp5_ASAP7_75t_L g5207 ( 
.A1(n_4833),
.A2(n_728),
.B(n_727),
.Y(n_5207)
);

AO32x2_ASAP7_75t_L g5208 ( 
.A1(n_4818),
.A2(n_729),
.A3(n_730),
.B1(n_728),
.B2(n_727),
.Y(n_5208)
);

NAND2xp5_ASAP7_75t_L g5209 ( 
.A(n_4724),
.B(n_4655),
.Y(n_5209)
);

INVx1_ASAP7_75t_SL g5210 ( 
.A(n_4822),
.Y(n_5210)
);

OAI21x1_ASAP7_75t_L g5211 ( 
.A1(n_4610),
.A2(n_729),
.B(n_728),
.Y(n_5211)
);

INVx3_ASAP7_75t_L g5212 ( 
.A(n_4662),
.Y(n_5212)
);

AOI21xp5_ASAP7_75t_L g5213 ( 
.A1(n_4612),
.A2(n_4635),
.B(n_4614),
.Y(n_5213)
);

BUFx2_ASAP7_75t_L g5214 ( 
.A(n_4503),
.Y(n_5214)
);

OR2x6_ASAP7_75t_L g5215 ( 
.A(n_4799),
.B(n_729),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_L g5216 ( 
.A(n_4677),
.B(n_4686),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_4691),
.B(n_1072),
.Y(n_5217)
);

AOI21xp5_ASAP7_75t_L g5218 ( 
.A1(n_4606),
.A2(n_731),
.B(n_730),
.Y(n_5218)
);

OA21x2_ASAP7_75t_L g5219 ( 
.A1(n_4710),
.A2(n_731),
.B(n_730),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_4827),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_4786),
.B(n_732),
.Y(n_5221)
);

INVx1_ASAP7_75t_SL g5222 ( 
.A(n_4520),
.Y(n_5222)
);

CKINVDCx5p33_ASAP7_75t_R g5223 ( 
.A(n_4849),
.Y(n_5223)
);

OAI22x1_ASAP7_75t_L g5224 ( 
.A1(n_4908),
.A2(n_4787),
.B1(n_4850),
.B2(n_4815),
.Y(n_5224)
);

AO31x2_ASAP7_75t_L g5225 ( 
.A1(n_4866),
.A2(n_733),
.A3(n_734),
.B(n_732),
.Y(n_5225)
);

OAI21xp5_ASAP7_75t_L g5226 ( 
.A1(n_4593),
.A2(n_733),
.B(n_732),
.Y(n_5226)
);

OR2x2_ASAP7_75t_L g5227 ( 
.A(n_4712),
.B(n_1071),
.Y(n_5227)
);

AOI21xp5_ASAP7_75t_L g5228 ( 
.A1(n_4909),
.A2(n_734),
.B(n_733),
.Y(n_5228)
);

NOR2xp33_ASAP7_75t_L g5229 ( 
.A(n_4881),
.B(n_17),
.Y(n_5229)
);

INVx2_ASAP7_75t_L g5230 ( 
.A(n_4703),
.Y(n_5230)
);

AOI21xp5_ASAP7_75t_L g5231 ( 
.A1(n_4942),
.A2(n_736),
.B(n_735),
.Y(n_5231)
);

NOR2xp33_ASAP7_75t_SL g5232 ( 
.A(n_4824),
.B(n_735),
.Y(n_5232)
);

AND2x4_ASAP7_75t_L g5233 ( 
.A(n_4575),
.B(n_735),
.Y(n_5233)
);

OAI21xp5_ASAP7_75t_L g5234 ( 
.A1(n_4636),
.A2(n_4920),
.B(n_4912),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_4573),
.Y(n_5235)
);

NOR2x1_ASAP7_75t_SL g5236 ( 
.A(n_4836),
.B(n_736),
.Y(n_5236)
);

CKINVDCx20_ASAP7_75t_R g5237 ( 
.A(n_5042),
.Y(n_5237)
);

INVx3_ASAP7_75t_L g5238 ( 
.A(n_5038),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5040),
.Y(n_5239)
);

AND2x2_ASAP7_75t_L g5240 ( 
.A(n_5172),
.B(n_4969),
.Y(n_5240)
);

AOI22xp33_ASAP7_75t_L g5241 ( 
.A1(n_5043),
.A2(n_4940),
.B1(n_5002),
.B2(n_4970),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_4981),
.Y(n_5242)
);

AOI221xp5_ASAP7_75t_L g5243 ( 
.A1(n_4959),
.A2(n_4882),
.B1(n_4873),
.B2(n_4917),
.C(n_4900),
.Y(n_5243)
);

OAI21x1_ASAP7_75t_L g5244 ( 
.A1(n_4957),
.A2(n_4784),
.B(n_4767),
.Y(n_5244)
);

OAI21x1_ASAP7_75t_L g5245 ( 
.A1(n_5010),
.A2(n_4695),
.B(n_4694),
.Y(n_5245)
);

INVxp67_ASAP7_75t_L g5246 ( 
.A(n_5063),
.Y(n_5246)
);

AOI22xp33_ASAP7_75t_L g5247 ( 
.A1(n_5118),
.A2(n_4905),
.B1(n_4855),
.B2(n_4744),
.Y(n_5247)
);

NAND2xp5_ASAP7_75t_L g5248 ( 
.A(n_4996),
.B(n_4906),
.Y(n_5248)
);

OAI21xp5_ASAP7_75t_L g5249 ( 
.A1(n_5041),
.A2(n_4823),
.B(n_4743),
.Y(n_5249)
);

O2A1O1Ixp33_ASAP7_75t_SL g5250 ( 
.A1(n_4962),
.A2(n_4586),
.B(n_4943),
.C(n_4805),
.Y(n_5250)
);

BUFx3_ASAP7_75t_L g5251 ( 
.A(n_4978),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_5013),
.Y(n_5252)
);

BUFx3_ASAP7_75t_L g5253 ( 
.A(n_4966),
.Y(n_5253)
);

NOR2xp33_ASAP7_75t_L g5254 ( 
.A(n_5068),
.B(n_4796),
.Y(n_5254)
);

AOI22xp5_ASAP7_75t_L g5255 ( 
.A1(n_5024),
.A2(n_4956),
.B1(n_5118),
.B2(n_5003),
.Y(n_5255)
);

INVx1_ASAP7_75t_L g5256 ( 
.A(n_5026),
.Y(n_5256)
);

CKINVDCx20_ASAP7_75t_R g5257 ( 
.A(n_5025),
.Y(n_5257)
);

HB1xp67_ASAP7_75t_L g5258 ( 
.A(n_5076),
.Y(n_5258)
);

OAI21x1_ASAP7_75t_L g5259 ( 
.A1(n_5065),
.A2(n_4728),
.B(n_4699),
.Y(n_5259)
);

OAI21x1_ASAP7_75t_L g5260 ( 
.A1(n_5064),
.A2(n_4802),
.B(n_4901),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_5060),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_5074),
.Y(n_5262)
);

AOI21xp5_ASAP7_75t_L g5263 ( 
.A1(n_4958),
.A2(n_4725),
.B(n_4721),
.Y(n_5263)
);

OAI21x1_ASAP7_75t_L g5264 ( 
.A1(n_5094),
.A2(n_4746),
.B(n_4751),
.Y(n_5264)
);

CKINVDCx5p33_ASAP7_75t_R g5265 ( 
.A(n_5047),
.Y(n_5265)
);

AO21x2_ASAP7_75t_L g5266 ( 
.A1(n_5141),
.A2(n_4742),
.B(n_4654),
.Y(n_5266)
);

OAI21xp5_ASAP7_75t_L g5267 ( 
.A1(n_5181),
.A2(n_5035),
.B(n_5030),
.Y(n_5267)
);

INVxp67_ASAP7_75t_SL g5268 ( 
.A(n_5129),
.Y(n_5268)
);

AND2x4_ASAP7_75t_L g5269 ( 
.A(n_5050),
.B(n_4520),
.Y(n_5269)
);

INVx2_ASAP7_75t_L g5270 ( 
.A(n_5061),
.Y(n_5270)
);

AO21x2_ASAP7_75t_L g5271 ( 
.A1(n_5097),
.A2(n_4651),
.B(n_4583),
.Y(n_5271)
);

INVx1_ASAP7_75t_L g5272 ( 
.A(n_5012),
.Y(n_5272)
);

OA21x2_ASAP7_75t_L g5273 ( 
.A1(n_4994),
.A2(n_5023),
.B(n_4961),
.Y(n_5273)
);

INVx1_ASAP7_75t_SL g5274 ( 
.A(n_5210),
.Y(n_5274)
);

OA21x2_ASAP7_75t_L g5275 ( 
.A1(n_5071),
.A2(n_4693),
.B(n_4585),
.Y(n_5275)
);

AOI21xp33_ASAP7_75t_L g5276 ( 
.A1(n_5079),
.A2(n_5224),
.B(n_5015),
.Y(n_5276)
);

OAI21x1_ASAP7_75t_L g5277 ( 
.A1(n_5009),
.A2(n_4781),
.B(n_4755),
.Y(n_5277)
);

INVx2_ASAP7_75t_L g5278 ( 
.A(n_5080),
.Y(n_5278)
);

BUFx12f_ASAP7_75t_L g5279 ( 
.A(n_5102),
.Y(n_5279)
);

OA21x2_ASAP7_75t_L g5280 ( 
.A1(n_4992),
.A2(n_4587),
.B(n_4579),
.Y(n_5280)
);

OR2x2_ASAP7_75t_L g5281 ( 
.A(n_5154),
.B(n_4926),
.Y(n_5281)
);

OAI21x1_ASAP7_75t_L g5282 ( 
.A1(n_4986),
.A2(n_4903),
.B(n_4925),
.Y(n_5282)
);

HB1xp67_ASAP7_75t_L g5283 ( 
.A(n_4967),
.Y(n_5283)
);

CKINVDCx5p33_ASAP7_75t_R g5284 ( 
.A(n_5067),
.Y(n_5284)
);

CKINVDCx20_ASAP7_75t_R g5285 ( 
.A(n_5223),
.Y(n_5285)
);

OAI21xp5_ASAP7_75t_L g5286 ( 
.A1(n_5112),
.A2(n_4922),
.B(n_4771),
.Y(n_5286)
);

AO21x2_ASAP7_75t_L g5287 ( 
.A1(n_5044),
.A2(n_4621),
.B(n_4615),
.Y(n_5287)
);

NAND2x1p5_ASAP7_75t_L g5288 ( 
.A(n_5053),
.B(n_4790),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_5160),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_L g5290 ( 
.A(n_5083),
.B(n_4688),
.Y(n_5290)
);

AOI22xp33_ASAP7_75t_L g5291 ( 
.A1(n_5118),
.A2(n_4936),
.B1(n_4531),
.B2(n_4611),
.Y(n_5291)
);

OAI221xp5_ASAP7_75t_L g5292 ( 
.A1(n_5073),
.A2(n_4780),
.B1(n_4831),
.B2(n_4948),
.C(n_4513),
.Y(n_5292)
);

NOR2xp33_ASAP7_75t_SL g5293 ( 
.A(n_5184),
.B(n_4876),
.Y(n_5293)
);

INVx2_ASAP7_75t_L g5294 ( 
.A(n_4952),
.Y(n_5294)
);

OR2x2_ASAP7_75t_L g5295 ( 
.A(n_5183),
.B(n_4520),
.Y(n_5295)
);

OAI21x1_ASAP7_75t_SL g5296 ( 
.A1(n_5165),
.A2(n_4571),
.B(n_4785),
.Y(n_5296)
);

INVx1_ASAP7_75t_L g5297 ( 
.A(n_5093),
.Y(n_5297)
);

INVx8_ASAP7_75t_L g5298 ( 
.A(n_5052),
.Y(n_5298)
);

OAI21x1_ASAP7_75t_L g5299 ( 
.A1(n_4960),
.A2(n_5005),
.B(n_5001),
.Y(n_5299)
);

AOI21xp5_ASAP7_75t_SL g5300 ( 
.A1(n_5186),
.A2(n_4791),
.B(n_4945),
.Y(n_5300)
);

OAI21x1_ASAP7_75t_L g5301 ( 
.A1(n_5022),
.A2(n_4938),
.B(n_4932),
.Y(n_5301)
);

OAI21x1_ASAP7_75t_L g5302 ( 
.A1(n_4987),
.A2(n_4735),
.B(n_4729),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_5027),
.Y(n_5303)
);

AOI22xp33_ASAP7_75t_L g5304 ( 
.A1(n_5131),
.A2(n_4792),
.B1(n_4794),
.B2(n_4884),
.Y(n_5304)
);

BUFx2_ASAP7_75t_L g5305 ( 
.A(n_4997),
.Y(n_5305)
);

AO21x2_ASAP7_75t_L g5306 ( 
.A1(n_5070),
.A2(n_4640),
.B(n_4630),
.Y(n_5306)
);

INVx2_ASAP7_75t_L g5307 ( 
.A(n_4977),
.Y(n_5307)
);

AO31x2_ASAP7_75t_L g5308 ( 
.A1(n_5143),
.A2(n_4665),
.A3(n_4928),
.B(n_4846),
.Y(n_5308)
);

OAI21x1_ASAP7_75t_L g5309 ( 
.A1(n_5058),
.A2(n_4756),
.B(n_4870),
.Y(n_5309)
);

CKINVDCx11_ASAP7_75t_R g5310 ( 
.A(n_5163),
.Y(n_5310)
);

NOR2xp67_ASAP7_75t_L g5311 ( 
.A(n_5053),
.B(n_4790),
.Y(n_5311)
);

INVx2_ASAP7_75t_L g5312 ( 
.A(n_5103),
.Y(n_5312)
);

AOI21x1_ASAP7_75t_L g5313 ( 
.A1(n_5155),
.A2(n_4880),
.B(n_4642),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_5116),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_4995),
.B(n_4934),
.Y(n_5315)
);

AOI22xp33_ASAP7_75t_L g5316 ( 
.A1(n_4979),
.A2(n_4889),
.B1(n_4939),
.B2(n_4646),
.Y(n_5316)
);

OAI21x1_ASAP7_75t_L g5317 ( 
.A1(n_4999),
.A2(n_4613),
.B(n_4907),
.Y(n_5317)
);

OAI21x1_ASAP7_75t_L g5318 ( 
.A1(n_5139),
.A2(n_4731),
.B(n_4879),
.Y(n_5318)
);

OAI21xp5_ASAP7_75t_L g5319 ( 
.A1(n_5078),
.A2(n_4601),
.B(n_4797),
.Y(n_5319)
);

INVx3_ASAP7_75t_L g5320 ( 
.A(n_5132),
.Y(n_5320)
);

AND2x6_ASAP7_75t_L g5321 ( 
.A(n_4975),
.B(n_4902),
.Y(n_5321)
);

NAND2x1p5_ASAP7_75t_L g5322 ( 
.A(n_5178),
.B(n_4656),
.Y(n_5322)
);

OR2x2_ASAP7_75t_L g5323 ( 
.A(n_4973),
.B(n_4533),
.Y(n_5323)
);

AOI21x1_ASAP7_75t_L g5324 ( 
.A1(n_5011),
.A2(n_4641),
.B(n_4644),
.Y(n_5324)
);

AND2x2_ASAP7_75t_L g5325 ( 
.A(n_5220),
.B(n_4533),
.Y(n_5325)
);

O2A1O1Ixp33_ASAP7_75t_SL g5326 ( 
.A1(n_5031),
.A2(n_4887),
.B(n_4670),
.C(n_4702),
.Y(n_5326)
);

OAI21x1_ASAP7_75t_L g5327 ( 
.A1(n_5185),
.A2(n_4863),
.B(n_4622),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_5124),
.Y(n_5328)
);

NAND2x1p5_ASAP7_75t_L g5329 ( 
.A(n_5178),
.B(n_4871),
.Y(n_5329)
);

AO21x2_ASAP7_75t_L g5330 ( 
.A1(n_5077),
.A2(n_4559),
.B(n_4546),
.Y(n_5330)
);

OAI21xp5_ASAP7_75t_L g5331 ( 
.A1(n_5111),
.A2(n_4916),
.B(n_4726),
.Y(n_5331)
);

OAI21x1_ASAP7_75t_L g5332 ( 
.A1(n_5006),
.A2(n_4658),
.B(n_4844),
.Y(n_5332)
);

OR2x6_ASAP7_75t_L g5333 ( 
.A(n_5150),
.B(n_5055),
.Y(n_5333)
);

OAI21x1_ASAP7_75t_L g5334 ( 
.A1(n_5213),
.A2(n_4965),
.B(n_5127),
.Y(n_5334)
);

AO21x2_ASAP7_75t_L g5335 ( 
.A1(n_5138),
.A2(n_4572),
.B(n_4541),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_5128),
.Y(n_5336)
);

INVx2_ASAP7_75t_L g5337 ( 
.A(n_5136),
.Y(n_5337)
);

AOI22xp33_ASAP7_75t_L g5338 ( 
.A1(n_5192),
.A2(n_4889),
.B1(n_4719),
.B2(n_4816),
.Y(n_5338)
);

AO21x2_ASAP7_75t_L g5339 ( 
.A1(n_5170),
.A2(n_4759),
.B(n_4775),
.Y(n_5339)
);

OAI21xp5_ASAP7_75t_L g5340 ( 
.A1(n_5207),
.A2(n_4804),
.B(n_4795),
.Y(n_5340)
);

BUFx3_ASAP7_75t_L g5341 ( 
.A(n_4985),
.Y(n_5341)
);

INVx3_ASAP7_75t_L g5342 ( 
.A(n_5082),
.Y(n_5342)
);

AOI21xp33_ASAP7_75t_L g5343 ( 
.A1(n_4954),
.A2(n_4808),
.B(n_4848),
.Y(n_5343)
);

INVx2_ASAP7_75t_L g5344 ( 
.A(n_5140),
.Y(n_5344)
);

AOI21xp33_ASAP7_75t_L g5345 ( 
.A1(n_5091),
.A2(n_4864),
.B(n_4857),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_5000),
.Y(n_5346)
);

INVx3_ASAP7_75t_L g5347 ( 
.A(n_4968),
.Y(n_5347)
);

NAND2x1p5_ASAP7_75t_L g5348 ( 
.A(n_5037),
.B(n_4533),
.Y(n_5348)
);

AOI21xp33_ASAP7_75t_L g5349 ( 
.A1(n_5036),
.A2(n_4893),
.B(n_4872),
.Y(n_5349)
);

OAI21x1_ASAP7_75t_L g5350 ( 
.A1(n_4976),
.A2(n_4902),
.B(n_4944),
.Y(n_5350)
);

OA21x2_ASAP7_75t_L g5351 ( 
.A1(n_4991),
.A2(n_4946),
.B(n_4623),
.Y(n_5351)
);

OAI22xp5_ASAP7_75t_SL g5352 ( 
.A1(n_5119),
.A2(n_4877),
.B1(n_4836),
.B2(n_4648),
.Y(n_5352)
);

BUFx6f_ASAP7_75t_L g5353 ( 
.A(n_4963),
.Y(n_5353)
);

INVx2_ASAP7_75t_L g5354 ( 
.A(n_4989),
.Y(n_5354)
);

OAI21x1_ASAP7_75t_L g5355 ( 
.A1(n_5151),
.A2(n_4902),
.B(n_4889),
.Y(n_5355)
);

NAND2xp5_ASAP7_75t_L g5356 ( 
.A(n_5235),
.B(n_4891),
.Y(n_5356)
);

AND2x2_ASAP7_75t_L g5357 ( 
.A(n_5201),
.B(n_4648),
.Y(n_5357)
);

NOR2xp33_ASAP7_75t_L g5358 ( 
.A(n_5229),
.B(n_4877),
.Y(n_5358)
);

OAI21x1_ASAP7_75t_L g5359 ( 
.A1(n_5174),
.A2(n_4766),
.B(n_4891),
.Y(n_5359)
);

OAI21x1_ASAP7_75t_L g5360 ( 
.A1(n_5175),
.A2(n_4766),
.B(n_4718),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_5032),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_4951),
.Y(n_5362)
);

INVx3_ASAP7_75t_L g5363 ( 
.A(n_5149),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_4964),
.Y(n_5364)
);

CKINVDCx5p33_ASAP7_75t_R g5365 ( 
.A(n_5161),
.Y(n_5365)
);

NAND2xp5_ASAP7_75t_L g5366 ( 
.A(n_4998),
.B(n_4877),
.Y(n_5366)
);

INVx2_ASAP7_75t_L g5367 ( 
.A(n_5007),
.Y(n_5367)
);

OAI21x1_ASAP7_75t_L g5368 ( 
.A1(n_5176),
.A2(n_4766),
.B(n_4718),
.Y(n_5368)
);

CKINVDCx20_ASAP7_75t_R g5369 ( 
.A(n_5190),
.Y(n_5369)
);

INVx1_ASAP7_75t_L g5370 ( 
.A(n_4980),
.Y(n_5370)
);

INVx2_ASAP7_75t_L g5371 ( 
.A(n_5054),
.Y(n_5371)
);

AOI21xp5_ASAP7_75t_L g5372 ( 
.A1(n_5086),
.A2(n_4648),
.B(n_4809),
.Y(n_5372)
);

HB1xp67_ASAP7_75t_L g5373 ( 
.A(n_5051),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_5142),
.Y(n_5374)
);

AND2x4_ASAP7_75t_L g5375 ( 
.A(n_5191),
.B(n_4809),
.Y(n_5375)
);

OR2x2_ASAP7_75t_L g5376 ( 
.A(n_5204),
.B(n_4809),
.Y(n_5376)
);

BUFx6f_ASAP7_75t_L g5377 ( 
.A(n_4963),
.Y(n_5377)
);

INVx2_ASAP7_75t_L g5378 ( 
.A(n_5148),
.Y(n_5378)
);

INVx2_ASAP7_75t_SL g5379 ( 
.A(n_5191),
.Y(n_5379)
);

OAI21x1_ASAP7_75t_L g5380 ( 
.A1(n_5182),
.A2(n_4718),
.B(n_4812),
.Y(n_5380)
);

OAI21x1_ASAP7_75t_L g5381 ( 
.A1(n_5230),
.A2(n_4812),
.B(n_4869),
.Y(n_5381)
);

OAI21xp33_ASAP7_75t_L g5382 ( 
.A1(n_5232),
.A2(n_4812),
.B(n_4778),
.Y(n_5382)
);

INVx2_ASAP7_75t_L g5383 ( 
.A(n_5214),
.Y(n_5383)
);

NAND3xp33_ASAP7_75t_L g5384 ( 
.A(n_5016),
.B(n_4778),
.C(n_4869),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_4993),
.Y(n_5385)
);

INVx3_ASAP7_75t_L g5386 ( 
.A(n_5233),
.Y(n_5386)
);

CKINVDCx5p33_ASAP7_75t_R g5387 ( 
.A(n_5194),
.Y(n_5387)
);

BUFx2_ASAP7_75t_L g5388 ( 
.A(n_5100),
.Y(n_5388)
);

INVx2_ASAP7_75t_L g5389 ( 
.A(n_5084),
.Y(n_5389)
);

INVx4_ASAP7_75t_L g5390 ( 
.A(n_5215),
.Y(n_5390)
);

AND2x4_ASAP7_75t_L g5391 ( 
.A(n_5180),
.B(n_736),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_5028),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_5028),
.Y(n_5393)
);

NAND2xp5_ASAP7_75t_L g5394 ( 
.A(n_5216),
.B(n_737),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_5099),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_5125),
.Y(n_5396)
);

CKINVDCx5p33_ASAP7_75t_R g5397 ( 
.A(n_5197),
.Y(n_5397)
);

OAI21x1_ASAP7_75t_L g5398 ( 
.A1(n_5014),
.A2(n_4869),
.B(n_4778),
.Y(n_5398)
);

OA21x2_ASAP7_75t_L g5399 ( 
.A1(n_5110),
.A2(n_738),
.B(n_737),
.Y(n_5399)
);

AOI21xp5_ASAP7_75t_L g5400 ( 
.A1(n_5019),
.A2(n_739),
.B(n_737),
.Y(n_5400)
);

OAI21x1_ASAP7_75t_L g5401 ( 
.A1(n_5018),
.A2(n_740),
.B(n_739),
.Y(n_5401)
);

INVx2_ASAP7_75t_L g5402 ( 
.A(n_5222),
.Y(n_5402)
);

NOR2xp33_ASAP7_75t_L g5403 ( 
.A(n_5101),
.B(n_739),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_5135),
.Y(n_5404)
);

O2A1O1Ixp33_ASAP7_75t_SL g5405 ( 
.A1(n_5146),
.A2(n_741),
.B(n_742),
.C(n_740),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5092),
.Y(n_5406)
);

OAI21x1_ASAP7_75t_L g5407 ( 
.A1(n_5021),
.A2(n_741),
.B(n_740),
.Y(n_5407)
);

A2O1A1Ixp33_ASAP7_75t_L g5408 ( 
.A1(n_5231),
.A2(n_5098),
.B(n_5162),
.C(n_5029),
.Y(n_5408)
);

OAI21x1_ASAP7_75t_L g5409 ( 
.A1(n_5066),
.A2(n_742),
.B(n_741),
.Y(n_5409)
);

AND2x2_ASAP7_75t_L g5410 ( 
.A(n_5240),
.B(n_5105),
.Y(n_5410)
);

INVx2_ASAP7_75t_L g5411 ( 
.A(n_5258),
.Y(n_5411)
);

OAI21x1_ASAP7_75t_L g5412 ( 
.A1(n_5299),
.A2(n_5045),
.B(n_5212),
.Y(n_5412)
);

INVx2_ASAP7_75t_L g5413 ( 
.A(n_5305),
.Y(n_5413)
);

AND2x2_ASAP7_75t_L g5414 ( 
.A(n_5283),
.B(n_5105),
.Y(n_5414)
);

AOI21x1_ASAP7_75t_L g5415 ( 
.A1(n_5313),
.A2(n_5033),
.B(n_5147),
.Y(n_5415)
);

AOI22xp33_ASAP7_75t_L g5416 ( 
.A1(n_5241),
.A2(n_5243),
.B1(n_5403),
.B2(n_5390),
.Y(n_5416)
);

OAI22xp5_ASAP7_75t_L g5417 ( 
.A1(n_5255),
.A2(n_5215),
.B1(n_5147),
.B2(n_5133),
.Y(n_5417)
);

INVx2_ASAP7_75t_L g5418 ( 
.A(n_5305),
.Y(n_5418)
);

INVx2_ASAP7_75t_L g5419 ( 
.A(n_5268),
.Y(n_5419)
);

BUFx2_ASAP7_75t_R g5420 ( 
.A(n_5251),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_5252),
.Y(n_5421)
);

INVx2_ASAP7_75t_L g5422 ( 
.A(n_5242),
.Y(n_5422)
);

OR2x2_ASAP7_75t_L g5423 ( 
.A(n_5239),
.B(n_5089),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5256),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5261),
.Y(n_5425)
);

NAND2xp5_ASAP7_75t_L g5426 ( 
.A(n_5385),
.B(n_4983),
.Y(n_5426)
);

AOI22xp33_ASAP7_75t_L g5427 ( 
.A1(n_5384),
.A2(n_4983),
.B1(n_5234),
.B2(n_5114),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_5262),
.Y(n_5428)
);

CKINVDCx5p33_ASAP7_75t_R g5429 ( 
.A(n_5279),
.Y(n_5429)
);

BUFx3_ASAP7_75t_L g5430 ( 
.A(n_5298),
.Y(n_5430)
);

BUFx4f_ASAP7_75t_SL g5431 ( 
.A(n_5257),
.Y(n_5431)
);

INVx2_ASAP7_75t_L g5432 ( 
.A(n_5270),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_5297),
.Y(n_5433)
);

INVx6_ASAP7_75t_L g5434 ( 
.A(n_5298),
.Y(n_5434)
);

BUFx12f_ASAP7_75t_L g5435 ( 
.A(n_5265),
.Y(n_5435)
);

OR2x6_ASAP7_75t_L g5436 ( 
.A(n_5379),
.B(n_5333),
.Y(n_5436)
);

INVx3_ASAP7_75t_L g5437 ( 
.A(n_5333),
.Y(n_5437)
);

HB1xp67_ASAP7_75t_L g5438 ( 
.A(n_5373),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5289),
.Y(n_5439)
);

AOI21x1_ASAP7_75t_L g5440 ( 
.A1(n_5313),
.A2(n_5311),
.B(n_5324),
.Y(n_5440)
);

OAI22xp33_ASAP7_75t_L g5441 ( 
.A1(n_5293),
.A2(n_4971),
.B1(n_5085),
.B2(n_5177),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_5312),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5337),
.Y(n_5443)
);

AO21x2_ASAP7_75t_L g5444 ( 
.A1(n_5354),
.A2(n_5193),
.B(n_5039),
.Y(n_5444)
);

NAND2x1p5_ASAP7_75t_L g5445 ( 
.A(n_5253),
.B(n_5238),
.Y(n_5445)
);

INVx4_ASAP7_75t_L g5446 ( 
.A(n_5320),
.Y(n_5446)
);

AOI22xp33_ASAP7_75t_SL g5447 ( 
.A1(n_5273),
.A2(n_5236),
.B1(n_4983),
.B2(n_5134),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5344),
.Y(n_5448)
);

INVxp67_ASAP7_75t_L g5449 ( 
.A(n_5254),
.Y(n_5449)
);

AND2x2_ASAP7_75t_L g5450 ( 
.A(n_5357),
.B(n_4971),
.Y(n_5450)
);

INVx2_ASAP7_75t_L g5451 ( 
.A(n_5278),
.Y(n_5451)
);

INVx1_ASAP7_75t_L g5452 ( 
.A(n_5314),
.Y(n_5452)
);

BUFx3_ASAP7_75t_L g5453 ( 
.A(n_5341),
.Y(n_5453)
);

CKINVDCx11_ASAP7_75t_R g5454 ( 
.A(n_5237),
.Y(n_5454)
);

AOI22xp33_ASAP7_75t_SL g5455 ( 
.A1(n_5273),
.A2(n_5219),
.B1(n_5203),
.B2(n_5188),
.Y(n_5455)
);

AOI22xp5_ASAP7_75t_L g5456 ( 
.A1(n_5382),
.A2(n_5057),
.B1(n_4982),
.B2(n_5209),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_5328),
.Y(n_5457)
);

INVx11_ASAP7_75t_L g5458 ( 
.A(n_5285),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_5336),
.Y(n_5459)
);

AOI22xp33_ASAP7_75t_SL g5460 ( 
.A1(n_5386),
.A2(n_5226),
.B1(n_5202),
.B2(n_5195),
.Y(n_5460)
);

NAND2x1p5_ASAP7_75t_L g5461 ( 
.A(n_5347),
.B(n_5227),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_5272),
.Y(n_5462)
);

AOI22xp33_ASAP7_75t_L g5463 ( 
.A1(n_5247),
.A2(n_5117),
.B1(n_4988),
.B2(n_5164),
.Y(n_5463)
);

AOI22xp33_ASAP7_75t_SL g5464 ( 
.A1(n_5342),
.A2(n_5352),
.B1(n_5369),
.B2(n_5249),
.Y(n_5464)
);

BUFx4_ASAP7_75t_R g5465 ( 
.A(n_5310),
.Y(n_5465)
);

OAI22xp5_ASAP7_75t_L g5466 ( 
.A1(n_5338),
.A2(n_5062),
.B1(n_5046),
.B2(n_5206),
.Y(n_5466)
);

AOI22xp33_ASAP7_75t_L g5467 ( 
.A1(n_5276),
.A2(n_5090),
.B1(n_5115),
.B2(n_5106),
.Y(n_5467)
);

BUFx2_ASAP7_75t_L g5468 ( 
.A(n_5269),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_5346),
.Y(n_5469)
);

HB1xp67_ASAP7_75t_L g5470 ( 
.A(n_5351),
.Y(n_5470)
);

INVx2_ASAP7_75t_L g5471 ( 
.A(n_5294),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5303),
.Y(n_5472)
);

BUFx2_ASAP7_75t_L g5473 ( 
.A(n_5269),
.Y(n_5473)
);

CKINVDCx20_ASAP7_75t_R g5474 ( 
.A(n_5284),
.Y(n_5474)
);

BUFx6f_ASAP7_75t_SL g5475 ( 
.A(n_5375),
.Y(n_5475)
);

INVx2_ASAP7_75t_L g5476 ( 
.A(n_5307),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_5362),
.Y(n_5477)
);

INVx1_ASAP7_75t_SL g5478 ( 
.A(n_5274),
.Y(n_5478)
);

OAI22xp5_ASAP7_75t_L g5479 ( 
.A1(n_5365),
.A2(n_5088),
.B1(n_5095),
.B2(n_5034),
.Y(n_5479)
);

NAND2xp5_ASAP7_75t_L g5480 ( 
.A(n_5364),
.B(n_5171),
.Y(n_5480)
);

AOI22xp33_ASAP7_75t_L g5481 ( 
.A1(n_5296),
.A2(n_5167),
.B1(n_5199),
.B2(n_5059),
.Y(n_5481)
);

OR2x2_ASAP7_75t_L g5482 ( 
.A(n_5370),
.B(n_5153),
.Y(n_5482)
);

AO21x1_ASAP7_75t_L g5483 ( 
.A1(n_5391),
.A2(n_5109),
.B(n_5104),
.Y(n_5483)
);

NAND2x1p5_ASAP7_75t_L g5484 ( 
.A(n_5363),
.B(n_5100),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5290),
.Y(n_5485)
);

OAI22xp5_ASAP7_75t_L g5486 ( 
.A1(n_5387),
.A2(n_5221),
.B1(n_5158),
.B2(n_5137),
.Y(n_5486)
);

INVx2_ASAP7_75t_L g5487 ( 
.A(n_5402),
.Y(n_5487)
);

CKINVDCx5p33_ASAP7_75t_R g5488 ( 
.A(n_5397),
.Y(n_5488)
);

OAI21x1_ASAP7_75t_L g5489 ( 
.A1(n_5355),
.A2(n_5048),
.B(n_4972),
.Y(n_5489)
);

BUFx6f_ASAP7_75t_L g5490 ( 
.A(n_5353),
.Y(n_5490)
);

INVx2_ASAP7_75t_L g5491 ( 
.A(n_5323),
.Y(n_5491)
);

INVx6_ASAP7_75t_L g5492 ( 
.A(n_5375),
.Y(n_5492)
);

AOI21x1_ASAP7_75t_L g5493 ( 
.A1(n_5324),
.A2(n_5228),
.B(n_5123),
.Y(n_5493)
);

OA21x2_ASAP7_75t_L g5494 ( 
.A1(n_5360),
.A2(n_5217),
.B(n_5069),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_5361),
.Y(n_5495)
);

HB1xp67_ASAP7_75t_L g5496 ( 
.A(n_5351),
.Y(n_5496)
);

NAND2x1_ASAP7_75t_L g5497 ( 
.A(n_5321),
.B(n_5122),
.Y(n_5497)
);

OA21x2_ASAP7_75t_L g5498 ( 
.A1(n_5368),
.A2(n_5159),
.B(n_5020),
.Y(n_5498)
);

INVx2_ASAP7_75t_L g5499 ( 
.A(n_5367),
.Y(n_5499)
);

OA21x2_ASAP7_75t_L g5500 ( 
.A1(n_5380),
.A2(n_5350),
.B(n_5381),
.Y(n_5500)
);

INVx3_ASAP7_75t_L g5501 ( 
.A(n_5288),
.Y(n_5501)
);

BUFx6f_ASAP7_75t_L g5502 ( 
.A(n_5353),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_5374),
.Y(n_5503)
);

OR2x2_ASAP7_75t_L g5504 ( 
.A(n_5281),
.B(n_5056),
.Y(n_5504)
);

INVx1_ASAP7_75t_L g5505 ( 
.A(n_5356),
.Y(n_5505)
);

BUFx3_ASAP7_75t_L g5506 ( 
.A(n_5329),
.Y(n_5506)
);

NOR2x1_ASAP7_75t_SL g5507 ( 
.A(n_5389),
.B(n_4955),
.Y(n_5507)
);

OAI22xp33_ASAP7_75t_L g5508 ( 
.A1(n_5267),
.A2(n_5246),
.B1(n_5292),
.B2(n_5263),
.Y(n_5508)
);

BUFx2_ASAP7_75t_R g5509 ( 
.A(n_5315),
.Y(n_5509)
);

OAI22xp5_ASAP7_75t_L g5510 ( 
.A1(n_5316),
.A2(n_5218),
.B1(n_5144),
.B2(n_5156),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_5248),
.Y(n_5511)
);

INVx1_ASAP7_75t_L g5512 ( 
.A(n_5325),
.Y(n_5512)
);

AOI22xp33_ASAP7_75t_L g5513 ( 
.A1(n_5296),
.A2(n_5087),
.B1(n_5168),
.B2(n_5152),
.Y(n_5513)
);

INVx2_ASAP7_75t_L g5514 ( 
.A(n_5371),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_5376),
.Y(n_5515)
);

BUFx2_ASAP7_75t_L g5516 ( 
.A(n_5388),
.Y(n_5516)
);

BUFx2_ASAP7_75t_L g5517 ( 
.A(n_5321),
.Y(n_5517)
);

INVx1_ASAP7_75t_SL g5518 ( 
.A(n_5322),
.Y(n_5518)
);

AOI22xp33_ASAP7_75t_L g5519 ( 
.A1(n_5343),
.A2(n_5189),
.B1(n_5121),
.B2(n_5113),
.Y(n_5519)
);

AOI22xp33_ASAP7_75t_SL g5520 ( 
.A1(n_5391),
.A2(n_4955),
.B1(n_5196),
.B2(n_5081),
.Y(n_5520)
);

BUFx3_ASAP7_75t_L g5521 ( 
.A(n_5388),
.Y(n_5521)
);

INVx1_ASAP7_75t_SL g5522 ( 
.A(n_5295),
.Y(n_5522)
);

AND2x4_ASAP7_75t_L g5523 ( 
.A(n_5378),
.B(n_4953),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_5406),
.Y(n_5524)
);

INVx3_ASAP7_75t_L g5525 ( 
.A(n_5377),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_5366),
.Y(n_5526)
);

OAI21xp5_ASAP7_75t_L g5527 ( 
.A1(n_5300),
.A2(n_5075),
.B(n_5049),
.Y(n_5527)
);

OR2x2_ASAP7_75t_L g5528 ( 
.A(n_5383),
.B(n_5056),
.Y(n_5528)
);

OAI22xp33_ASAP7_75t_L g5529 ( 
.A1(n_5286),
.A2(n_5348),
.B1(n_5275),
.B2(n_5280),
.Y(n_5529)
);

OR2x2_ASAP7_75t_L g5530 ( 
.A(n_5395),
.B(n_5396),
.Y(n_5530)
);

AND2x2_ASAP7_75t_L g5531 ( 
.A(n_5404),
.B(n_4953),
.Y(n_5531)
);

OAI21x1_ASAP7_75t_L g5532 ( 
.A1(n_5334),
.A2(n_5072),
.B(n_5120),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_5392),
.Y(n_5533)
);

CKINVDCx20_ASAP7_75t_R g5534 ( 
.A(n_5358),
.Y(n_5534)
);

INVx2_ASAP7_75t_L g5535 ( 
.A(n_5393),
.Y(n_5535)
);

INVx1_ASAP7_75t_SL g5536 ( 
.A(n_5377),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_5472),
.Y(n_5537)
);

OR2x2_ASAP7_75t_L g5538 ( 
.A(n_5438),
.B(n_5280),
.Y(n_5538)
);

BUFx5_ASAP7_75t_L g5539 ( 
.A(n_5506),
.Y(n_5539)
);

INVx4_ASAP7_75t_R g5540 ( 
.A(n_5430),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5442),
.Y(n_5541)
);

INVx6_ASAP7_75t_L g5542 ( 
.A(n_5434),
.Y(n_5542)
);

AOI22xp33_ASAP7_75t_L g5543 ( 
.A1(n_5450),
.A2(n_5275),
.B1(n_5271),
.B2(n_5291),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_5443),
.Y(n_5544)
);

AOI22xp33_ASAP7_75t_SL g5545 ( 
.A1(n_5446),
.A2(n_5321),
.B1(n_5399),
.B2(n_5335),
.Y(n_5545)
);

OAI21xp5_ASAP7_75t_SL g5546 ( 
.A1(n_5464),
.A2(n_5304),
.B(n_5400),
.Y(n_5546)
);

INVx2_ASAP7_75t_L g5547 ( 
.A(n_5419),
.Y(n_5547)
);

AOI22xp33_ASAP7_75t_L g5548 ( 
.A1(n_5441),
.A2(n_5345),
.B1(n_5399),
.B2(n_5339),
.Y(n_5548)
);

AND2x2_ASAP7_75t_L g5549 ( 
.A(n_5522),
.B(n_5266),
.Y(n_5549)
);

NAND2xp5_ASAP7_75t_L g5550 ( 
.A(n_5531),
.B(n_5330),
.Y(n_5550)
);

AND2x2_ASAP7_75t_L g5551 ( 
.A(n_5468),
.B(n_5359),
.Y(n_5551)
);

OAI22xp5_ASAP7_75t_L g5552 ( 
.A1(n_5436),
.A2(n_5408),
.B1(n_5372),
.B2(n_5394),
.Y(n_5552)
);

AOI22xp33_ASAP7_75t_L g5553 ( 
.A1(n_5416),
.A2(n_5508),
.B1(n_5417),
.B2(n_5527),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_5448),
.Y(n_5554)
);

AOI22xp33_ASAP7_75t_L g5555 ( 
.A1(n_5520),
.A2(n_5340),
.B1(n_5349),
.B2(n_5287),
.Y(n_5555)
);

OAI21xp5_ASAP7_75t_L g5556 ( 
.A1(n_5415),
.A2(n_5332),
.B(n_5282),
.Y(n_5556)
);

AOI22xp33_ASAP7_75t_SL g5557 ( 
.A1(n_5437),
.A2(n_5306),
.B1(n_5398),
.B2(n_5245),
.Y(n_5557)
);

INVx2_ASAP7_75t_L g5558 ( 
.A(n_5411),
.Y(n_5558)
);

AOI22xp33_ASAP7_75t_L g5559 ( 
.A1(n_5427),
.A2(n_5331),
.B1(n_5319),
.B2(n_5302),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5524),
.Y(n_5560)
);

AOI222xp33_ASAP7_75t_L g5561 ( 
.A1(n_5486),
.A2(n_5327),
.B1(n_5318),
.B2(n_5317),
.C1(n_5301),
.C2(n_5401),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_5462),
.Y(n_5562)
);

AOI22xp33_ASAP7_75t_L g5563 ( 
.A1(n_5460),
.A2(n_5244),
.B1(n_5309),
.B2(n_5260),
.Y(n_5563)
);

AOI22xp33_ASAP7_75t_SL g5564 ( 
.A1(n_5436),
.A2(n_5264),
.B1(n_5277),
.B2(n_5407),
.Y(n_5564)
);

OAI22xp5_ASAP7_75t_L g5565 ( 
.A1(n_5509),
.A2(n_4990),
.B1(n_5250),
.B2(n_5208),
.Y(n_5565)
);

OAI22xp5_ASAP7_75t_L g5566 ( 
.A1(n_5447),
.A2(n_5208),
.B1(n_5405),
.B2(n_5096),
.Y(n_5566)
);

HB1xp67_ASAP7_75t_L g5567 ( 
.A(n_5468),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_5530),
.Y(n_5568)
);

INVx2_ASAP7_75t_L g5569 ( 
.A(n_5473),
.Y(n_5569)
);

HB1xp67_ASAP7_75t_L g5570 ( 
.A(n_5473),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_5469),
.Y(n_5571)
);

INVx2_ASAP7_75t_L g5572 ( 
.A(n_5422),
.Y(n_5572)
);

INVx8_ASAP7_75t_L g5573 ( 
.A(n_5435),
.Y(n_5573)
);

BUFx4f_ASAP7_75t_SL g5574 ( 
.A(n_5474),
.Y(n_5574)
);

AOI22xp33_ASAP7_75t_L g5575 ( 
.A1(n_5483),
.A2(n_5259),
.B1(n_5409),
.B2(n_5108),
.Y(n_5575)
);

OAI222xp33_ASAP7_75t_L g5576 ( 
.A1(n_5529),
.A2(n_5225),
.B1(n_5326),
.B2(n_4984),
.C1(n_5187),
.C2(n_5145),
.Y(n_5576)
);

OAI21xp5_ASAP7_75t_SL g5577 ( 
.A1(n_5445),
.A2(n_4984),
.B(n_5173),
.Y(n_5577)
);

AOI22xp33_ASAP7_75t_L g5578 ( 
.A1(n_5510),
.A2(n_5107),
.B1(n_5157),
.B2(n_5130),
.Y(n_5578)
);

AOI22xp33_ASAP7_75t_L g5579 ( 
.A1(n_5481),
.A2(n_5463),
.B1(n_5466),
.B2(n_5467),
.Y(n_5579)
);

AOI22xp33_ASAP7_75t_L g5580 ( 
.A1(n_5513),
.A2(n_5444),
.B1(n_5511),
.B2(n_5426),
.Y(n_5580)
);

BUFx2_ASAP7_75t_L g5581 ( 
.A(n_5453),
.Y(n_5581)
);

OAI22xp5_ASAP7_75t_L g5582 ( 
.A1(n_5518),
.A2(n_5225),
.B1(n_5145),
.B2(n_5198),
.Y(n_5582)
);

AOI22xp5_ASAP7_75t_L g5583 ( 
.A1(n_5456),
.A2(n_5479),
.B1(n_5410),
.B2(n_5449),
.Y(n_5583)
);

AOI22xp33_ASAP7_75t_SL g5584 ( 
.A1(n_5507),
.A2(n_5205),
.B1(n_5211),
.B2(n_5200),
.Y(n_5584)
);

AOI22xp33_ASAP7_75t_SL g5585 ( 
.A1(n_5475),
.A2(n_5169),
.B1(n_5179),
.B2(n_5126),
.Y(n_5585)
);

INVx2_ASAP7_75t_L g5586 ( 
.A(n_5432),
.Y(n_5586)
);

AOI22xp33_ASAP7_75t_L g5587 ( 
.A1(n_5455),
.A2(n_5166),
.B1(n_5308),
.B2(n_5008),
.Y(n_5587)
);

AND2x2_ASAP7_75t_L g5588 ( 
.A(n_5491),
.B(n_5187),
.Y(n_5588)
);

AOI222xp33_ASAP7_75t_L g5589 ( 
.A1(n_5485),
.A2(n_5308),
.B1(n_746),
.B2(n_744),
.C1(n_747),
.C2(n_745),
.Y(n_5589)
);

BUFx3_ASAP7_75t_L g5590 ( 
.A(n_5431),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5477),
.Y(n_5591)
);

AOI22xp33_ASAP7_75t_L g5592 ( 
.A1(n_5512),
.A2(n_5308),
.B1(n_5017),
.B2(n_4974),
.Y(n_5592)
);

AOI22xp33_ASAP7_75t_L g5593 ( 
.A1(n_5515),
.A2(n_5017),
.B1(n_4974),
.B2(n_5004),
.Y(n_5593)
);

OR2x2_ASAP7_75t_L g5594 ( 
.A(n_5413),
.B(n_5004),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_5421),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_5451),
.Y(n_5596)
);

INVx2_ASAP7_75t_L g5597 ( 
.A(n_5471),
.Y(n_5597)
);

OR2x2_ASAP7_75t_L g5598 ( 
.A(n_5418),
.B(n_743),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5476),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_5535),
.Y(n_5600)
);

AOI22xp33_ASAP7_75t_L g5601 ( 
.A1(n_5519),
.A2(n_744),
.B1(n_746),
.B2(n_743),
.Y(n_5601)
);

INVx2_ASAP7_75t_SL g5602 ( 
.A(n_5434),
.Y(n_5602)
);

AOI22xp33_ASAP7_75t_SL g5603 ( 
.A1(n_5470),
.A2(n_747),
.B1(n_748),
.B2(n_746),
.Y(n_5603)
);

AOI222xp33_ASAP7_75t_L g5604 ( 
.A1(n_5480),
.A2(n_750),
.B1(n_748),
.B2(n_751),
.C1(n_749),
.C2(n_747),
.Y(n_5604)
);

AOI22xp33_ASAP7_75t_L g5605 ( 
.A1(n_5505),
.A2(n_5494),
.B1(n_5526),
.B2(n_5478),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5424),
.Y(n_5606)
);

BUFx6f_ASAP7_75t_L g5607 ( 
.A(n_5490),
.Y(n_5607)
);

HB1xp67_ASAP7_75t_L g5608 ( 
.A(n_5496),
.Y(n_5608)
);

AOI22xp33_ASAP7_75t_L g5609 ( 
.A1(n_5494),
.A2(n_749),
.B1(n_750),
.B2(n_748),
.Y(n_5609)
);

NAND2xp5_ASAP7_75t_L g5610 ( 
.A(n_5495),
.B(n_749),
.Y(n_5610)
);

INVx4_ASAP7_75t_L g5611 ( 
.A(n_5465),
.Y(n_5611)
);

INVx2_ASAP7_75t_L g5612 ( 
.A(n_5528),
.Y(n_5612)
);

AOI22xp33_ASAP7_75t_L g5613 ( 
.A1(n_5461),
.A2(n_751),
.B1(n_752),
.B2(n_750),
.Y(n_5613)
);

NAND2xp5_ASAP7_75t_L g5614 ( 
.A(n_5503),
.B(n_751),
.Y(n_5614)
);

BUFx12f_ASAP7_75t_L g5615 ( 
.A(n_5429),
.Y(n_5615)
);

OAI22xp5_ASAP7_75t_SL g5616 ( 
.A1(n_5488),
.A2(n_754),
.B1(n_755),
.B2(n_753),
.Y(n_5616)
);

AOI22xp33_ASAP7_75t_SL g5617 ( 
.A1(n_5517),
.A2(n_754),
.B1(n_755),
.B2(n_753),
.Y(n_5617)
);

INVxp67_ASAP7_75t_SL g5618 ( 
.A(n_5516),
.Y(n_5618)
);

AOI22xp33_ASAP7_75t_L g5619 ( 
.A1(n_5504),
.A2(n_755),
.B1(n_756),
.B2(n_754),
.Y(n_5619)
);

AOI22xp33_ASAP7_75t_SL g5620 ( 
.A1(n_5517),
.A2(n_758),
.B1(n_759),
.B2(n_757),
.Y(n_5620)
);

BUFx4f_ASAP7_75t_SL g5621 ( 
.A(n_5534),
.Y(n_5621)
);

INVx6_ASAP7_75t_L g5622 ( 
.A(n_5490),
.Y(n_5622)
);

AOI22xp33_ASAP7_75t_SL g5623 ( 
.A1(n_5492),
.A2(n_758),
.B1(n_759),
.B2(n_757),
.Y(n_5623)
);

AOI22xp33_ASAP7_75t_L g5624 ( 
.A1(n_5414),
.A2(n_759),
.B1(n_760),
.B2(n_757),
.Y(n_5624)
);

NAND2xp5_ASAP7_75t_SL g5625 ( 
.A(n_5440),
.B(n_17),
.Y(n_5625)
);

AND2x2_ASAP7_75t_L g5626 ( 
.A(n_5521),
.B(n_760),
.Y(n_5626)
);

INVx1_ASAP7_75t_L g5627 ( 
.A(n_5425),
.Y(n_5627)
);

BUFx4f_ASAP7_75t_SL g5628 ( 
.A(n_5420),
.Y(n_5628)
);

AOI22xp33_ASAP7_75t_L g5629 ( 
.A1(n_5497),
.A2(n_762),
.B1(n_763),
.B2(n_760),
.Y(n_5629)
);

AOI22xp33_ASAP7_75t_L g5630 ( 
.A1(n_5533),
.A2(n_764),
.B1(n_765),
.B2(n_762),
.Y(n_5630)
);

AOI22xp33_ASAP7_75t_L g5631 ( 
.A1(n_5423),
.A2(n_765),
.B1(n_766),
.B2(n_764),
.Y(n_5631)
);

BUFx4f_ASAP7_75t_SL g5632 ( 
.A(n_5454),
.Y(n_5632)
);

INVx2_ASAP7_75t_L g5633 ( 
.A(n_5487),
.Y(n_5633)
);

HB1xp67_ASAP7_75t_L g5634 ( 
.A(n_5499),
.Y(n_5634)
);

AND2x2_ASAP7_75t_L g5635 ( 
.A(n_5514),
.B(n_764),
.Y(n_5635)
);

AOI22xp33_ASAP7_75t_SL g5636 ( 
.A1(n_5492),
.A2(n_766),
.B1(n_767),
.B2(n_765),
.Y(n_5636)
);

INVx2_ASAP7_75t_L g5637 ( 
.A(n_5523),
.Y(n_5637)
);

CKINVDCx11_ASAP7_75t_R g5638 ( 
.A(n_5458),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_5428),
.Y(n_5639)
);

OAI21xp5_ASAP7_75t_SL g5640 ( 
.A1(n_5501),
.A2(n_768),
.B(n_767),
.Y(n_5640)
);

NAND2xp5_ASAP7_75t_L g5641 ( 
.A(n_5543),
.B(n_5433),
.Y(n_5641)
);

INVx1_ASAP7_75t_L g5642 ( 
.A(n_5537),
.Y(n_5642)
);

INVxp67_ASAP7_75t_L g5643 ( 
.A(n_5581),
.Y(n_5643)
);

AND2x4_ASAP7_75t_L g5644 ( 
.A(n_5611),
.B(n_5536),
.Y(n_5644)
);

NAND2xp33_ASAP7_75t_R g5645 ( 
.A(n_5628),
.B(n_5412),
.Y(n_5645)
);

OR2x6_ASAP7_75t_L g5646 ( 
.A(n_5573),
.B(n_5484),
.Y(n_5646)
);

INVx1_ASAP7_75t_L g5647 ( 
.A(n_5541),
.Y(n_5647)
);

AND2x4_ASAP7_75t_L g5648 ( 
.A(n_5611),
.B(n_5525),
.Y(n_5648)
);

BUFx3_ASAP7_75t_L g5649 ( 
.A(n_5573),
.Y(n_5649)
);

OR2x6_ASAP7_75t_L g5650 ( 
.A(n_5542),
.B(n_5493),
.Y(n_5650)
);

AND2x4_ASAP7_75t_L g5651 ( 
.A(n_5602),
.B(n_5502),
.Y(n_5651)
);

XNOR2x2_ASAP7_75t_L g5652 ( 
.A(n_5556),
.B(n_5482),
.Y(n_5652)
);

AND2x2_ASAP7_75t_L g5653 ( 
.A(n_5549),
.B(n_5523),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_5544),
.Y(n_5654)
);

BUFx3_ASAP7_75t_L g5655 ( 
.A(n_5574),
.Y(n_5655)
);

OR2x6_ASAP7_75t_L g5656 ( 
.A(n_5542),
.B(n_5502),
.Y(n_5656)
);

NAND2xp33_ASAP7_75t_R g5657 ( 
.A(n_5540),
.B(n_5626),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_5554),
.Y(n_5658)
);

BUFx3_ASAP7_75t_L g5659 ( 
.A(n_5632),
.Y(n_5659)
);

BUFx10_ASAP7_75t_L g5660 ( 
.A(n_5622),
.Y(n_5660)
);

NAND2xp5_ASAP7_75t_L g5661 ( 
.A(n_5583),
.B(n_5439),
.Y(n_5661)
);

NOR2xp33_ASAP7_75t_R g5662 ( 
.A(n_5638),
.B(n_18),
.Y(n_5662)
);

NAND2xp33_ASAP7_75t_R g5663 ( 
.A(n_5539),
.B(n_5500),
.Y(n_5663)
);

NOR2xp33_ASAP7_75t_R g5664 ( 
.A(n_5621),
.B(n_18),
.Y(n_5664)
);

BUFx2_ASAP7_75t_L g5665 ( 
.A(n_5539),
.Y(n_5665)
);

NAND2xp33_ASAP7_75t_SL g5666 ( 
.A(n_5567),
.B(n_5452),
.Y(n_5666)
);

AND2x4_ASAP7_75t_L g5667 ( 
.A(n_5568),
.B(n_5457),
.Y(n_5667)
);

NAND2xp33_ASAP7_75t_R g5668 ( 
.A(n_5539),
.B(n_5500),
.Y(n_5668)
);

NAND2xp5_ASAP7_75t_L g5669 ( 
.A(n_5588),
.B(n_5459),
.Y(n_5669)
);

INVx2_ASAP7_75t_L g5670 ( 
.A(n_5634),
.Y(n_5670)
);

AND2x4_ASAP7_75t_L g5671 ( 
.A(n_5590),
.B(n_5532),
.Y(n_5671)
);

NAND2xp33_ASAP7_75t_R g5672 ( 
.A(n_5539),
.B(n_5498),
.Y(n_5672)
);

NAND2xp5_ASAP7_75t_L g5673 ( 
.A(n_5550),
.B(n_5498),
.Y(n_5673)
);

AND2x4_ASAP7_75t_L g5674 ( 
.A(n_5618),
.B(n_5607),
.Y(n_5674)
);

BUFx3_ASAP7_75t_L g5675 ( 
.A(n_5615),
.Y(n_5675)
);

NAND2xp5_ASAP7_75t_L g5676 ( 
.A(n_5555),
.B(n_5489),
.Y(n_5676)
);

AND2x4_ASAP7_75t_L g5677 ( 
.A(n_5607),
.B(n_5635),
.Y(n_5677)
);

NAND2xp5_ASAP7_75t_L g5678 ( 
.A(n_5580),
.B(n_5548),
.Y(n_5678)
);

NAND2xp33_ASAP7_75t_R g5679 ( 
.A(n_5539),
.B(n_18),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5595),
.Y(n_5680)
);

HB1xp67_ASAP7_75t_L g5681 ( 
.A(n_5570),
.Y(n_5681)
);

NAND2xp5_ASAP7_75t_L g5682 ( 
.A(n_5612),
.B(n_769),
.Y(n_5682)
);

NAND2xp5_ASAP7_75t_SL g5683 ( 
.A(n_5545),
.B(n_18),
.Y(n_5683)
);

NOR2xp33_ASAP7_75t_R g5684 ( 
.A(n_5622),
.B(n_19),
.Y(n_5684)
);

AND2x4_ASAP7_75t_L g5685 ( 
.A(n_5607),
.B(n_769),
.Y(n_5685)
);

NOR2xp33_ASAP7_75t_R g5686 ( 
.A(n_5553),
.B(n_19),
.Y(n_5686)
);

NAND2xp5_ASAP7_75t_L g5687 ( 
.A(n_5605),
.B(n_770),
.Y(n_5687)
);

NAND2xp5_ASAP7_75t_SL g5688 ( 
.A(n_5557),
.B(n_19),
.Y(n_5688)
);

NAND2xp33_ASAP7_75t_R g5689 ( 
.A(n_5538),
.B(n_19),
.Y(n_5689)
);

NAND2xp5_ASAP7_75t_L g5690 ( 
.A(n_5579),
.B(n_770),
.Y(n_5690)
);

BUFx10_ASAP7_75t_L g5691 ( 
.A(n_5640),
.Y(n_5691)
);

BUFx6f_ASAP7_75t_L g5692 ( 
.A(n_5625),
.Y(n_5692)
);

NOR2xp33_ASAP7_75t_R g5693 ( 
.A(n_5559),
.B(n_20),
.Y(n_5693)
);

NOR2xp33_ASAP7_75t_R g5694 ( 
.A(n_5629),
.B(n_20),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_5606),
.Y(n_5695)
);

AND2x2_ASAP7_75t_L g5696 ( 
.A(n_5551),
.B(n_20),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_5627),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5639),
.Y(n_5698)
);

BUFx10_ASAP7_75t_L g5699 ( 
.A(n_5616),
.Y(n_5699)
);

XOR2xp5_ASAP7_75t_L g5700 ( 
.A(n_5565),
.B(n_20),
.Y(n_5700)
);

INVxp67_ASAP7_75t_L g5701 ( 
.A(n_5552),
.Y(n_5701)
);

NOR2xp33_ASAP7_75t_R g5702 ( 
.A(n_5613),
.B(n_21),
.Y(n_5702)
);

NOR2xp33_ASAP7_75t_R g5703 ( 
.A(n_5598),
.B(n_21),
.Y(n_5703)
);

INVxp67_ASAP7_75t_L g5704 ( 
.A(n_5610),
.Y(n_5704)
);

INVx2_ASAP7_75t_L g5705 ( 
.A(n_5594),
.Y(n_5705)
);

AND2x4_ASAP7_75t_L g5706 ( 
.A(n_5569),
.B(n_771),
.Y(n_5706)
);

NAND2xp5_ASAP7_75t_SL g5707 ( 
.A(n_5564),
.B(n_21),
.Y(n_5707)
);

INVx2_ASAP7_75t_L g5708 ( 
.A(n_5600),
.Y(n_5708)
);

INVx3_ASAP7_75t_L g5709 ( 
.A(n_5547),
.Y(n_5709)
);

AND2x2_ASAP7_75t_L g5710 ( 
.A(n_5637),
.B(n_22),
.Y(n_5710)
);

XNOR2xp5_ASAP7_75t_L g5711 ( 
.A(n_5617),
.B(n_22),
.Y(n_5711)
);

INVx3_ASAP7_75t_L g5712 ( 
.A(n_5572),
.Y(n_5712)
);

NOR2xp33_ASAP7_75t_R g5713 ( 
.A(n_5614),
.B(n_22),
.Y(n_5713)
);

BUFx8_ASAP7_75t_SL g5714 ( 
.A(n_5558),
.Y(n_5714)
);

NOR2xp33_ASAP7_75t_R g5715 ( 
.A(n_5619),
.B(n_22),
.Y(n_5715)
);

NAND2xp33_ASAP7_75t_R g5716 ( 
.A(n_5546),
.B(n_23),
.Y(n_5716)
);

AND2x2_ASAP7_75t_L g5717 ( 
.A(n_5644),
.B(n_5608),
.Y(n_5717)
);

AND2x2_ASAP7_75t_L g5718 ( 
.A(n_5648),
.B(n_5563),
.Y(n_5718)
);

BUFx3_ASAP7_75t_L g5719 ( 
.A(n_5659),
.Y(n_5719)
);

BUFx2_ASAP7_75t_L g5720 ( 
.A(n_5656),
.Y(n_5720)
);

INVxp67_ASAP7_75t_SL g5721 ( 
.A(n_5679),
.Y(n_5721)
);

AND2x2_ASAP7_75t_L g5722 ( 
.A(n_5643),
.B(n_5561),
.Y(n_5722)
);

AND2x2_ASAP7_75t_L g5723 ( 
.A(n_5674),
.B(n_5633),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5647),
.Y(n_5724)
);

INVx3_ASAP7_75t_L g5725 ( 
.A(n_5646),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_5654),
.Y(n_5726)
);

AND2x2_ASAP7_75t_L g5727 ( 
.A(n_5653),
.B(n_5560),
.Y(n_5727)
);

BUFx3_ASAP7_75t_L g5728 ( 
.A(n_5649),
.Y(n_5728)
);

NAND2xp5_ASAP7_75t_L g5729 ( 
.A(n_5701),
.B(n_5575),
.Y(n_5729)
);

NOR4xp25_ASAP7_75t_SL g5730 ( 
.A(n_5645),
.B(n_5577),
.C(n_5571),
.D(n_5562),
.Y(n_5730)
);

OAI21xp33_ASAP7_75t_L g5731 ( 
.A1(n_5678),
.A2(n_5587),
.B(n_5584),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5681),
.Y(n_5732)
);

NAND2x1p5_ASAP7_75t_L g5733 ( 
.A(n_5685),
.B(n_5591),
.Y(n_5733)
);

BUFx2_ASAP7_75t_L g5734 ( 
.A(n_5656),
.Y(n_5734)
);

INVx4_ASAP7_75t_SL g5735 ( 
.A(n_5646),
.Y(n_5735)
);

INVx2_ASAP7_75t_L g5736 ( 
.A(n_5712),
.Y(n_5736)
);

INVx2_ASAP7_75t_L g5737 ( 
.A(n_5709),
.Y(n_5737)
);

AO21x2_ASAP7_75t_L g5738 ( 
.A1(n_5676),
.A2(n_5576),
.B(n_5582),
.Y(n_5738)
);

BUFx6f_ASAP7_75t_L g5739 ( 
.A(n_5675),
.Y(n_5739)
);

INVx2_ASAP7_75t_L g5740 ( 
.A(n_5670),
.Y(n_5740)
);

NOR2x1p5_ASAP7_75t_L g5741 ( 
.A(n_5655),
.B(n_5586),
.Y(n_5741)
);

INVx2_ASAP7_75t_L g5742 ( 
.A(n_5705),
.Y(n_5742)
);

HB1xp67_ASAP7_75t_L g5743 ( 
.A(n_5689),
.Y(n_5743)
);

INVx2_ASAP7_75t_L g5744 ( 
.A(n_5708),
.Y(n_5744)
);

INVx2_ASAP7_75t_L g5745 ( 
.A(n_5667),
.Y(n_5745)
);

INVxp67_ASAP7_75t_L g5746 ( 
.A(n_5696),
.Y(n_5746)
);

BUFx3_ASAP7_75t_L g5747 ( 
.A(n_5714),
.Y(n_5747)
);

AND2x2_ASAP7_75t_L g5748 ( 
.A(n_5671),
.B(n_5596),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5658),
.Y(n_5749)
);

HB1xp67_ASAP7_75t_L g5750 ( 
.A(n_5642),
.Y(n_5750)
);

INVx1_ASAP7_75t_L g5751 ( 
.A(n_5680),
.Y(n_5751)
);

NAND2xp5_ASAP7_75t_L g5752 ( 
.A(n_5641),
.B(n_5592),
.Y(n_5752)
);

INVx1_ASAP7_75t_L g5753 ( 
.A(n_5695),
.Y(n_5753)
);

BUFx3_ASAP7_75t_L g5754 ( 
.A(n_5651),
.Y(n_5754)
);

INVx2_ASAP7_75t_L g5755 ( 
.A(n_5665),
.Y(n_5755)
);

AND2x2_ASAP7_75t_L g5756 ( 
.A(n_5660),
.B(n_5597),
.Y(n_5756)
);

CKINVDCx5p33_ASAP7_75t_R g5757 ( 
.A(n_5662),
.Y(n_5757)
);

INVx2_ASAP7_75t_L g5758 ( 
.A(n_5697),
.Y(n_5758)
);

AOI22xp5_ASAP7_75t_L g5759 ( 
.A1(n_5716),
.A2(n_5566),
.B1(n_5589),
.B2(n_5585),
.Y(n_5759)
);

AND2x2_ASAP7_75t_L g5760 ( 
.A(n_5677),
.B(n_5599),
.Y(n_5760)
);

INVx2_ASAP7_75t_L g5761 ( 
.A(n_5698),
.Y(n_5761)
);

INVx1_ASAP7_75t_L g5762 ( 
.A(n_5669),
.Y(n_5762)
);

AND2x4_ASAP7_75t_L g5763 ( 
.A(n_5650),
.B(n_5578),
.Y(n_5763)
);

OR2x6_ASAP7_75t_L g5764 ( 
.A(n_5707),
.B(n_5623),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_5682),
.Y(n_5765)
);

AND2x2_ASAP7_75t_L g5766 ( 
.A(n_5704),
.B(n_5593),
.Y(n_5766)
);

HB1xp67_ASAP7_75t_L g5767 ( 
.A(n_5692),
.Y(n_5767)
);

AND2x2_ASAP7_75t_L g5768 ( 
.A(n_5710),
.B(n_5624),
.Y(n_5768)
);

OR2x2_ASAP7_75t_L g5769 ( 
.A(n_5661),
.B(n_5609),
.Y(n_5769)
);

INVxp67_ASAP7_75t_SL g5770 ( 
.A(n_5692),
.Y(n_5770)
);

AND2x2_ASAP7_75t_L g5771 ( 
.A(n_5650),
.B(n_5601),
.Y(n_5771)
);

OR2x2_ASAP7_75t_L g5772 ( 
.A(n_5673),
.B(n_5631),
.Y(n_5772)
);

NOR2x1_ASAP7_75t_SL g5773 ( 
.A(n_5683),
.B(n_5620),
.Y(n_5773)
);

NOR2x1_ASAP7_75t_SL g5774 ( 
.A(n_5688),
.B(n_5636),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5687),
.Y(n_5775)
);

INVx2_ASAP7_75t_SL g5776 ( 
.A(n_5684),
.Y(n_5776)
);

AO21x2_ASAP7_75t_L g5777 ( 
.A1(n_5700),
.A2(n_5664),
.B(n_5686),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_5706),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_5690),
.Y(n_5779)
);

AND2x2_ASAP7_75t_L g5780 ( 
.A(n_5691),
.B(n_5604),
.Y(n_5780)
);

HB1xp67_ASAP7_75t_L g5781 ( 
.A(n_5657),
.Y(n_5781)
);

AND2x2_ASAP7_75t_L g5782 ( 
.A(n_5699),
.B(n_5703),
.Y(n_5782)
);

BUFx6f_ASAP7_75t_L g5783 ( 
.A(n_5711),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_5666),
.Y(n_5784)
);

NOR2x1_ASAP7_75t_SL g5785 ( 
.A(n_5652),
.B(n_5603),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5693),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_5713),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_5694),
.Y(n_5788)
);

INVx2_ASAP7_75t_L g5789 ( 
.A(n_5672),
.Y(n_5789)
);

NAND2xp5_ASAP7_75t_L g5790 ( 
.A(n_5715),
.B(n_5630),
.Y(n_5790)
);

INVx1_ASAP7_75t_L g5791 ( 
.A(n_5702),
.Y(n_5791)
);

AND2x4_ASAP7_75t_L g5792 ( 
.A(n_5663),
.B(n_771),
.Y(n_5792)
);

INVx2_ASAP7_75t_L g5793 ( 
.A(n_5668),
.Y(n_5793)
);

CKINVDCx5p33_ASAP7_75t_R g5794 ( 
.A(n_5659),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_5647),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5647),
.Y(n_5796)
);

INVx3_ASAP7_75t_L g5797 ( 
.A(n_5646),
.Y(n_5797)
);

INVx3_ASAP7_75t_L g5798 ( 
.A(n_5646),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5647),
.Y(n_5799)
);

AND2x2_ASAP7_75t_L g5800 ( 
.A(n_5644),
.B(n_23),
.Y(n_5800)
);

HB1xp67_ASAP7_75t_L g5801 ( 
.A(n_5681),
.Y(n_5801)
);

NAND2xp5_ASAP7_75t_L g5802 ( 
.A(n_5701),
.B(n_23),
.Y(n_5802)
);

HB1xp67_ASAP7_75t_L g5803 ( 
.A(n_5681),
.Y(n_5803)
);

AND2x2_ASAP7_75t_SL g5804 ( 
.A(n_5792),
.B(n_771),
.Y(n_5804)
);

NAND2xp5_ASAP7_75t_L g5805 ( 
.A(n_5779),
.B(n_23),
.Y(n_5805)
);

INVx2_ASAP7_75t_L g5806 ( 
.A(n_5741),
.Y(n_5806)
);

BUFx2_ASAP7_75t_L g5807 ( 
.A(n_5735),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5801),
.Y(n_5808)
);

INVx2_ASAP7_75t_L g5809 ( 
.A(n_5740),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5744),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5803),
.Y(n_5811)
);

BUFx2_ASAP7_75t_L g5812 ( 
.A(n_5735),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_5732),
.Y(n_5813)
);

INVx2_ASAP7_75t_SL g5814 ( 
.A(n_5747),
.Y(n_5814)
);

AND2x2_ASAP7_75t_L g5815 ( 
.A(n_5725),
.B(n_24),
.Y(n_5815)
);

BUFx2_ASAP7_75t_L g5816 ( 
.A(n_5725),
.Y(n_5816)
);

INVx2_ASAP7_75t_SL g5817 ( 
.A(n_5719),
.Y(n_5817)
);

INVx2_ASAP7_75t_L g5818 ( 
.A(n_5717),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5742),
.Y(n_5819)
);

NAND2xp5_ASAP7_75t_L g5820 ( 
.A(n_5779),
.B(n_5775),
.Y(n_5820)
);

AND2x2_ASAP7_75t_L g5821 ( 
.A(n_5797),
.B(n_24),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5750),
.Y(n_5822)
);

AND2x2_ASAP7_75t_L g5823 ( 
.A(n_5797),
.B(n_24),
.Y(n_5823)
);

INVx2_ASAP7_75t_L g5824 ( 
.A(n_5733),
.Y(n_5824)
);

NOR2xp33_ASAP7_75t_L g5825 ( 
.A(n_5739),
.B(n_25),
.Y(n_5825)
);

INVx2_ASAP7_75t_L g5826 ( 
.A(n_5755),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_5802),
.Y(n_5827)
);

INVx1_ASAP7_75t_L g5828 ( 
.A(n_5767),
.Y(n_5828)
);

INVx1_ASAP7_75t_L g5829 ( 
.A(n_5724),
.Y(n_5829)
);

OR2x2_ASAP7_75t_L g5830 ( 
.A(n_5772),
.B(n_25),
.Y(n_5830)
);

INVx1_ASAP7_75t_L g5831 ( 
.A(n_5724),
.Y(n_5831)
);

OAI22xp5_ASAP7_75t_L g5832 ( 
.A1(n_5781),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_5832)
);

INVx1_ASAP7_75t_L g5833 ( 
.A(n_5726),
.Y(n_5833)
);

HB1xp67_ASAP7_75t_L g5834 ( 
.A(n_5743),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5726),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5795),
.Y(n_5836)
);

INVx2_ASAP7_75t_L g5837 ( 
.A(n_5723),
.Y(n_5837)
);

AND2x2_ASAP7_75t_L g5838 ( 
.A(n_5798),
.B(n_26),
.Y(n_5838)
);

AND2x4_ASAP7_75t_L g5839 ( 
.A(n_5798),
.B(n_772),
.Y(n_5839)
);

BUFx2_ASAP7_75t_SL g5840 ( 
.A(n_5728),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5795),
.Y(n_5841)
);

OR2x2_ASAP7_75t_L g5842 ( 
.A(n_5769),
.B(n_26),
.Y(n_5842)
);

INVx1_ASAP7_75t_L g5843 ( 
.A(n_5796),
.Y(n_5843)
);

INVxp67_ASAP7_75t_SL g5844 ( 
.A(n_5774),
.Y(n_5844)
);

NAND2xp5_ASAP7_75t_L g5845 ( 
.A(n_5775),
.B(n_26),
.Y(n_5845)
);

NAND2xp5_ASAP7_75t_L g5846 ( 
.A(n_5731),
.B(n_27),
.Y(n_5846)
);

NAND3xp33_ASAP7_75t_SL g5847 ( 
.A(n_5730),
.B(n_28),
.C(n_29),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5796),
.Y(n_5848)
);

AND2x2_ASAP7_75t_L g5849 ( 
.A(n_5720),
.B(n_28),
.Y(n_5849)
);

AND2x2_ASAP7_75t_L g5850 ( 
.A(n_5734),
.B(n_28),
.Y(n_5850)
);

BUFx2_ASAP7_75t_L g5851 ( 
.A(n_5754),
.Y(n_5851)
);

NAND2xp5_ASAP7_75t_L g5852 ( 
.A(n_5780),
.B(n_29),
.Y(n_5852)
);

BUFx2_ASAP7_75t_L g5853 ( 
.A(n_5770),
.Y(n_5853)
);

OR2x2_ASAP7_75t_L g5854 ( 
.A(n_5762),
.B(n_29),
.Y(n_5854)
);

OR2x2_ASAP7_75t_L g5855 ( 
.A(n_5729),
.B(n_30),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5799),
.Y(n_5856)
);

NAND2xp5_ASAP7_75t_L g5857 ( 
.A(n_5766),
.B(n_5722),
.Y(n_5857)
);

INVx2_ASAP7_75t_L g5858 ( 
.A(n_5758),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5799),
.Y(n_5859)
);

HB1xp67_ASAP7_75t_L g5860 ( 
.A(n_5761),
.Y(n_5860)
);

HB1xp67_ASAP7_75t_L g5861 ( 
.A(n_5749),
.Y(n_5861)
);

NAND2xp5_ASAP7_75t_L g5862 ( 
.A(n_5721),
.B(n_30),
.Y(n_5862)
);

INVx1_ASAP7_75t_L g5863 ( 
.A(n_5751),
.Y(n_5863)
);

INVx2_ASAP7_75t_L g5864 ( 
.A(n_5778),
.Y(n_5864)
);

NOR2xp33_ASAP7_75t_R g5865 ( 
.A(n_5794),
.B(n_30),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_5753),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5800),
.Y(n_5867)
);

HB1xp67_ASAP7_75t_L g5868 ( 
.A(n_5765),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5746),
.Y(n_5869)
);

AND2x4_ASAP7_75t_SL g5870 ( 
.A(n_5739),
.B(n_30),
.Y(n_5870)
);

NAND2xp5_ASAP7_75t_L g5871 ( 
.A(n_5759),
.B(n_31),
.Y(n_5871)
);

NAND2xp5_ASAP7_75t_SL g5872 ( 
.A(n_5792),
.B(n_31),
.Y(n_5872)
);

AND2x2_ASAP7_75t_L g5873 ( 
.A(n_5718),
.B(n_31),
.Y(n_5873)
);

HB1xp67_ASAP7_75t_L g5874 ( 
.A(n_5788),
.Y(n_5874)
);

INVx3_ASAP7_75t_L g5875 ( 
.A(n_5739),
.Y(n_5875)
);

AND2x2_ASAP7_75t_L g5876 ( 
.A(n_5771),
.B(n_31),
.Y(n_5876)
);

NAND2xp5_ASAP7_75t_L g5877 ( 
.A(n_5785),
.B(n_32),
.Y(n_5877)
);

INVx1_ASAP7_75t_L g5878 ( 
.A(n_5756),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_5776),
.Y(n_5879)
);

BUFx3_ASAP7_75t_L g5880 ( 
.A(n_5757),
.Y(n_5880)
);

BUFx3_ASAP7_75t_L g5881 ( 
.A(n_5787),
.Y(n_5881)
);

CKINVDCx5p33_ASAP7_75t_R g5882 ( 
.A(n_5783),
.Y(n_5882)
);

AND2x4_ASAP7_75t_L g5883 ( 
.A(n_5745),
.B(n_772),
.Y(n_5883)
);

HB1xp67_ASAP7_75t_L g5884 ( 
.A(n_5791),
.Y(n_5884)
);

HB1xp67_ASAP7_75t_L g5885 ( 
.A(n_5793),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5768),
.Y(n_5886)
);

OR2x2_ASAP7_75t_L g5887 ( 
.A(n_5738),
.B(n_32),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5727),
.Y(n_5888)
);

NAND2xp5_ASAP7_75t_L g5889 ( 
.A(n_5785),
.B(n_32),
.Y(n_5889)
);

AND2x4_ASAP7_75t_L g5890 ( 
.A(n_5782),
.B(n_772),
.Y(n_5890)
);

AND2x2_ASAP7_75t_L g5891 ( 
.A(n_5763),
.B(n_32),
.Y(n_5891)
);

INVxp67_ASAP7_75t_SL g5892 ( 
.A(n_5774),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5736),
.Y(n_5893)
);

NAND2xp5_ASAP7_75t_L g5894 ( 
.A(n_5752),
.B(n_33),
.Y(n_5894)
);

NOR3xp33_ASAP7_75t_L g5895 ( 
.A(n_5786),
.B(n_33),
.C(n_34),
.Y(n_5895)
);

INVx2_ASAP7_75t_L g5896 ( 
.A(n_5737),
.Y(n_5896)
);

INVx1_ASAP7_75t_L g5897 ( 
.A(n_5760),
.Y(n_5897)
);

NAND2xp5_ASAP7_75t_L g5898 ( 
.A(n_5763),
.B(n_33),
.Y(n_5898)
);

INVx1_ASAP7_75t_L g5899 ( 
.A(n_5790),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5786),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_5784),
.Y(n_5901)
);

INVxp67_ASAP7_75t_SL g5902 ( 
.A(n_5773),
.Y(n_5902)
);

INVx1_ASAP7_75t_L g5903 ( 
.A(n_5748),
.Y(n_5903)
);

INVx1_ASAP7_75t_L g5904 ( 
.A(n_5773),
.Y(n_5904)
);

AND2x2_ASAP7_75t_L g5905 ( 
.A(n_5789),
.B(n_5777),
.Y(n_5905)
);

NOR2xp33_ASAP7_75t_L g5906 ( 
.A(n_5783),
.B(n_34),
.Y(n_5906)
);

AND2x2_ASAP7_75t_L g5907 ( 
.A(n_5764),
.B(n_34),
.Y(n_5907)
);

AND2x2_ASAP7_75t_L g5908 ( 
.A(n_5764),
.B(n_35),
.Y(n_5908)
);

INVx1_ASAP7_75t_L g5909 ( 
.A(n_5783),
.Y(n_5909)
);

INVx2_ASAP7_75t_L g5910 ( 
.A(n_5741),
.Y(n_5910)
);

OR2x2_ASAP7_75t_L g5911 ( 
.A(n_5772),
.B(n_35),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5803),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5803),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5801),
.Y(n_5914)
);

INVx2_ASAP7_75t_L g5915 ( 
.A(n_5881),
.Y(n_5915)
);

AND2x2_ASAP7_75t_L g5916 ( 
.A(n_5840),
.B(n_5807),
.Y(n_5916)
);

INVx1_ASAP7_75t_SL g5917 ( 
.A(n_5812),
.Y(n_5917)
);

INVx3_ASAP7_75t_L g5918 ( 
.A(n_5880),
.Y(n_5918)
);

AND2x2_ASAP7_75t_L g5919 ( 
.A(n_5817),
.B(n_35),
.Y(n_5919)
);

INVx2_ASAP7_75t_L g5920 ( 
.A(n_5853),
.Y(n_5920)
);

AND2x2_ASAP7_75t_L g5921 ( 
.A(n_5851),
.B(n_35),
.Y(n_5921)
);

INVx2_ASAP7_75t_L g5922 ( 
.A(n_5816),
.Y(n_5922)
);

AND2x4_ASAP7_75t_L g5923 ( 
.A(n_5814),
.B(n_773),
.Y(n_5923)
);

NOR2x1_ASAP7_75t_L g5924 ( 
.A(n_5875),
.B(n_36),
.Y(n_5924)
);

NAND2xp5_ASAP7_75t_L g5925 ( 
.A(n_5834),
.B(n_36),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5815),
.Y(n_5926)
);

AND2x2_ASAP7_75t_L g5927 ( 
.A(n_5909),
.B(n_36),
.Y(n_5927)
);

AND2x2_ASAP7_75t_L g5928 ( 
.A(n_5909),
.B(n_36),
.Y(n_5928)
);

NAND2xp5_ASAP7_75t_L g5929 ( 
.A(n_5891),
.B(n_37),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5839),
.Y(n_5930)
);

AND2x2_ASAP7_75t_L g5931 ( 
.A(n_5875),
.B(n_37),
.Y(n_5931)
);

AND2x2_ASAP7_75t_L g5932 ( 
.A(n_5879),
.B(n_37),
.Y(n_5932)
);

OR2x2_ASAP7_75t_L g5933 ( 
.A(n_5898),
.B(n_37),
.Y(n_5933)
);

NAND2xp5_ASAP7_75t_L g5934 ( 
.A(n_5876),
.B(n_38),
.Y(n_5934)
);

AND2x2_ASAP7_75t_L g5935 ( 
.A(n_5806),
.B(n_5910),
.Y(n_5935)
);

INVx2_ASAP7_75t_SL g5936 ( 
.A(n_5882),
.Y(n_5936)
);

AND2x2_ASAP7_75t_L g5937 ( 
.A(n_5902),
.B(n_38),
.Y(n_5937)
);

NAND2xp5_ASAP7_75t_L g5938 ( 
.A(n_5874),
.B(n_38),
.Y(n_5938)
);

HB1xp67_ASAP7_75t_L g5939 ( 
.A(n_5884),
.Y(n_5939)
);

NAND2xp5_ASAP7_75t_L g5940 ( 
.A(n_5873),
.B(n_5900),
.Y(n_5940)
);

AND2x2_ASAP7_75t_L g5941 ( 
.A(n_5844),
.B(n_38),
.Y(n_5941)
);

NAND2xp5_ASAP7_75t_L g5942 ( 
.A(n_5886),
.B(n_39),
.Y(n_5942)
);

INVx2_ASAP7_75t_L g5943 ( 
.A(n_5839),
.Y(n_5943)
);

NAND2xp5_ASAP7_75t_L g5944 ( 
.A(n_5899),
.B(n_39),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5821),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_5892),
.B(n_39),
.Y(n_5946)
);

HB1xp67_ASAP7_75t_L g5947 ( 
.A(n_5849),
.Y(n_5947)
);

AND2x2_ASAP7_75t_L g5948 ( 
.A(n_5905),
.B(n_39),
.Y(n_5948)
);

OAI221xp5_ASAP7_75t_SL g5949 ( 
.A1(n_5904),
.A2(n_775),
.B1(n_776),
.B2(n_774),
.C(n_773),
.Y(n_5949)
);

NAND2x1p5_ASAP7_75t_L g5950 ( 
.A(n_5872),
.B(n_5804),
.Y(n_5950)
);

AND2x2_ASAP7_75t_L g5951 ( 
.A(n_5878),
.B(n_40),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5823),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5838),
.Y(n_5953)
);

NAND2xp5_ASAP7_75t_L g5954 ( 
.A(n_5877),
.B(n_40),
.Y(n_5954)
);

AND2x2_ASAP7_75t_L g5955 ( 
.A(n_5890),
.B(n_40),
.Y(n_5955)
);

INVx2_ASAP7_75t_L g5956 ( 
.A(n_5828),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5850),
.Y(n_5957)
);

AND2x4_ASAP7_75t_SL g5958 ( 
.A(n_5890),
.B(n_40),
.Y(n_5958)
);

NOR2xp33_ASAP7_75t_L g5959 ( 
.A(n_5889),
.B(n_5857),
.Y(n_5959)
);

OR2x2_ASAP7_75t_L g5960 ( 
.A(n_5842),
.B(n_41),
.Y(n_5960)
);

AND2x2_ASAP7_75t_L g5961 ( 
.A(n_5824),
.B(n_41),
.Y(n_5961)
);

INVx2_ASAP7_75t_L g5962 ( 
.A(n_5896),
.Y(n_5962)
);

HB1xp67_ASAP7_75t_L g5963 ( 
.A(n_5808),
.Y(n_5963)
);

AND2x2_ASAP7_75t_L g5964 ( 
.A(n_5837),
.B(n_41),
.Y(n_5964)
);

INVx2_ASAP7_75t_L g5965 ( 
.A(n_5826),
.Y(n_5965)
);

INVx1_ASAP7_75t_L g5966 ( 
.A(n_5808),
.Y(n_5966)
);

OR2x2_ASAP7_75t_L g5967 ( 
.A(n_5830),
.B(n_5911),
.Y(n_5967)
);

NAND2xp5_ASAP7_75t_L g5968 ( 
.A(n_5827),
.B(n_42),
.Y(n_5968)
);

OR2x2_ASAP7_75t_L g5969 ( 
.A(n_5852),
.B(n_42),
.Y(n_5969)
);

OR2x2_ASAP7_75t_L g5970 ( 
.A(n_5871),
.B(n_42),
.Y(n_5970)
);

AND2x2_ASAP7_75t_L g5971 ( 
.A(n_5818),
.B(n_43),
.Y(n_5971)
);

OR2x2_ASAP7_75t_L g5972 ( 
.A(n_5894),
.B(n_43),
.Y(n_5972)
);

AND2x2_ASAP7_75t_L g5973 ( 
.A(n_5907),
.B(n_43),
.Y(n_5973)
);

AND2x2_ASAP7_75t_L g5974 ( 
.A(n_5908),
.B(n_43),
.Y(n_5974)
);

HB1xp67_ASAP7_75t_L g5975 ( 
.A(n_5912),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_5912),
.Y(n_5976)
);

NAND2xp5_ASAP7_75t_L g5977 ( 
.A(n_5887),
.B(n_44),
.Y(n_5977)
);

AND2x4_ASAP7_75t_L g5978 ( 
.A(n_5864),
.B(n_773),
.Y(n_5978)
);

AND2x4_ASAP7_75t_SL g5979 ( 
.A(n_5867),
.B(n_44),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5913),
.Y(n_5980)
);

INVx1_ASAP7_75t_L g5981 ( 
.A(n_5913),
.Y(n_5981)
);

AND2x2_ASAP7_75t_L g5982 ( 
.A(n_5885),
.B(n_44),
.Y(n_5982)
);

INVx1_ASAP7_75t_L g5983 ( 
.A(n_5862),
.Y(n_5983)
);

HB1xp67_ASAP7_75t_L g5984 ( 
.A(n_5811),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_5914),
.Y(n_5985)
);

AND2x2_ASAP7_75t_L g5986 ( 
.A(n_5897),
.B(n_44),
.Y(n_5986)
);

NAND2xp5_ASAP7_75t_L g5987 ( 
.A(n_5846),
.B(n_45),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5868),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5819),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5861),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5869),
.Y(n_5991)
);

NAND2xp5_ASAP7_75t_L g5992 ( 
.A(n_5855),
.B(n_45),
.Y(n_5992)
);

INVx2_ASAP7_75t_L g5993 ( 
.A(n_5809),
.Y(n_5993)
);

NAND2xp5_ASAP7_75t_L g5994 ( 
.A(n_5888),
.B(n_45),
.Y(n_5994)
);

NAND2xp5_ASAP7_75t_L g5995 ( 
.A(n_5901),
.B(n_45),
.Y(n_5995)
);

NAND2xp5_ASAP7_75t_L g5996 ( 
.A(n_5820),
.B(n_46),
.Y(n_5996)
);

AND2x2_ASAP7_75t_L g5997 ( 
.A(n_5903),
.B(n_46),
.Y(n_5997)
);

AND2x2_ASAP7_75t_L g5998 ( 
.A(n_5893),
.B(n_46),
.Y(n_5998)
);

AND2x2_ASAP7_75t_L g5999 ( 
.A(n_5883),
.B(n_46),
.Y(n_5999)
);

NAND2xp5_ASAP7_75t_L g6000 ( 
.A(n_5822),
.B(n_47),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5859),
.Y(n_6001)
);

NAND2xp5_ASAP7_75t_L g6002 ( 
.A(n_5813),
.B(n_47),
.Y(n_6002)
);

AND2x2_ASAP7_75t_L g6003 ( 
.A(n_5883),
.B(n_47),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5859),
.Y(n_6004)
);

INVx2_ASAP7_75t_L g6005 ( 
.A(n_5810),
.Y(n_6005)
);

AND2x4_ASAP7_75t_L g6006 ( 
.A(n_5870),
.B(n_774),
.Y(n_6006)
);

AND2x4_ASAP7_75t_L g6007 ( 
.A(n_5916),
.B(n_5825),
.Y(n_6007)
);

AND2x2_ASAP7_75t_L g6008 ( 
.A(n_5918),
.B(n_5906),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5921),
.Y(n_6009)
);

BUFx3_ASAP7_75t_L g6010 ( 
.A(n_5918),
.Y(n_6010)
);

OR2x2_ASAP7_75t_L g6011 ( 
.A(n_5925),
.B(n_5832),
.Y(n_6011)
);

AND2x2_ASAP7_75t_L g6012 ( 
.A(n_5936),
.B(n_5915),
.Y(n_6012)
);

AND2x2_ASAP7_75t_L g6013 ( 
.A(n_5917),
.B(n_5865),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5963),
.Y(n_6014)
);

AND2x2_ASAP7_75t_L g6015 ( 
.A(n_5937),
.B(n_5860),
.Y(n_6015)
);

AND2x2_ASAP7_75t_L g6016 ( 
.A(n_5941),
.B(n_5805),
.Y(n_6016)
);

AND2x2_ASAP7_75t_L g6017 ( 
.A(n_5946),
.B(n_5845),
.Y(n_6017)
);

AND2x2_ASAP7_75t_L g6018 ( 
.A(n_5948),
.B(n_5854),
.Y(n_6018)
);

INVx2_ASAP7_75t_L g6019 ( 
.A(n_5920),
.Y(n_6019)
);

OR2x2_ASAP7_75t_L g6020 ( 
.A(n_5967),
.B(n_5858),
.Y(n_6020)
);

BUFx3_ASAP7_75t_L g6021 ( 
.A(n_5919),
.Y(n_6021)
);

INVx2_ASAP7_75t_SL g6022 ( 
.A(n_5931),
.Y(n_6022)
);

INVxp67_ASAP7_75t_SL g6023 ( 
.A(n_5938),
.Y(n_6023)
);

AND2x4_ASAP7_75t_L g6024 ( 
.A(n_5935),
.B(n_5930),
.Y(n_6024)
);

AND2x2_ASAP7_75t_L g6025 ( 
.A(n_5950),
.B(n_5895),
.Y(n_6025)
);

AND2x2_ASAP7_75t_L g6026 ( 
.A(n_5927),
.B(n_5863),
.Y(n_6026)
);

AND2x4_ASAP7_75t_SL g6027 ( 
.A(n_5961),
.B(n_5866),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_5928),
.B(n_5829),
.Y(n_6028)
);

AND2x4_ASAP7_75t_L g6029 ( 
.A(n_5943),
.B(n_5856),
.Y(n_6029)
);

NAND2xp5_ASAP7_75t_L g6030 ( 
.A(n_5922),
.B(n_5831),
.Y(n_6030)
);

OR2x2_ASAP7_75t_L g6031 ( 
.A(n_5957),
.B(n_5847),
.Y(n_6031)
);

INVx1_ASAP7_75t_L g6032 ( 
.A(n_5939),
.Y(n_6032)
);

INVx3_ASAP7_75t_L g6033 ( 
.A(n_5923),
.Y(n_6033)
);

INVx1_ASAP7_75t_L g6034 ( 
.A(n_5982),
.Y(n_6034)
);

HB1xp67_ASAP7_75t_L g6035 ( 
.A(n_5975),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_5923),
.Y(n_6036)
);

INVx2_ASAP7_75t_L g6037 ( 
.A(n_5965),
.Y(n_6037)
);

INVx2_ASAP7_75t_SL g6038 ( 
.A(n_5958),
.Y(n_6038)
);

INVx2_ASAP7_75t_L g6039 ( 
.A(n_5962),
.Y(n_6039)
);

AND2x2_ASAP7_75t_L g6040 ( 
.A(n_5947),
.B(n_5833),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5998),
.B(n_5835),
.Y(n_6041)
);

AND2x2_ASAP7_75t_L g6042 ( 
.A(n_5932),
.B(n_5836),
.Y(n_6042)
);

AND2x2_ASAP7_75t_L g6043 ( 
.A(n_5945),
.B(n_5841),
.Y(n_6043)
);

INVxp67_ASAP7_75t_L g6044 ( 
.A(n_5924),
.Y(n_6044)
);

AND2x2_ASAP7_75t_L g6045 ( 
.A(n_5945),
.B(n_5843),
.Y(n_6045)
);

AND2x2_ASAP7_75t_L g6046 ( 
.A(n_5952),
.B(n_5848),
.Y(n_6046)
);

INVx2_ASAP7_75t_L g6047 ( 
.A(n_5989),
.Y(n_6047)
);

NAND2x1p5_ASAP7_75t_L g6048 ( 
.A(n_6006),
.B(n_774),
.Y(n_6048)
);

AND2x2_ASAP7_75t_L g6049 ( 
.A(n_5952),
.B(n_47),
.Y(n_6049)
);

NOR2xp67_ASAP7_75t_L g6050 ( 
.A(n_5988),
.B(n_48),
.Y(n_6050)
);

AOI22xp33_ASAP7_75t_L g6051 ( 
.A1(n_5959),
.A2(n_776),
.B1(n_777),
.B2(n_775),
.Y(n_6051)
);

INVx2_ASAP7_75t_L g6052 ( 
.A(n_5993),
.Y(n_6052)
);

INVx1_ASAP7_75t_L g6053 ( 
.A(n_5984),
.Y(n_6053)
);

NAND2xp5_ASAP7_75t_L g6054 ( 
.A(n_5953),
.B(n_5978),
.Y(n_6054)
);

AND2x2_ASAP7_75t_L g6055 ( 
.A(n_5953),
.B(n_48),
.Y(n_6055)
);

AND4x1_ASAP7_75t_L g6056 ( 
.A(n_5983),
.B(n_51),
.C(n_49),
.D(n_50),
.Y(n_6056)
);

NOR2xp33_ASAP7_75t_R g6057 ( 
.A(n_5955),
.B(n_49),
.Y(n_6057)
);

OR2x2_ASAP7_75t_L g6058 ( 
.A(n_5942),
.B(n_49),
.Y(n_6058)
);

NAND2xp5_ASAP7_75t_L g6059 ( 
.A(n_5978),
.B(n_49),
.Y(n_6059)
);

INVx4_ASAP7_75t_L g6060 ( 
.A(n_6006),
.Y(n_6060)
);

AND2x2_ASAP7_75t_L g6061 ( 
.A(n_5951),
.B(n_50),
.Y(n_6061)
);

INVx2_ASAP7_75t_L g6062 ( 
.A(n_6005),
.Y(n_6062)
);

NAND2xp5_ASAP7_75t_L g6063 ( 
.A(n_5926),
.B(n_5988),
.Y(n_6063)
);

AOI22xp5_ASAP7_75t_L g6064 ( 
.A1(n_5940),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_5964),
.Y(n_6065)
);

NAND2xp5_ASAP7_75t_L g6066 ( 
.A(n_5956),
.B(n_5986),
.Y(n_6066)
);

INVx1_ASAP7_75t_L g6067 ( 
.A(n_5971),
.Y(n_6067)
);

AND2x2_ASAP7_75t_L g6068 ( 
.A(n_5997),
.B(n_50),
.Y(n_6068)
);

NAND2xp5_ASAP7_75t_SL g6069 ( 
.A(n_5990),
.B(n_5985),
.Y(n_6069)
);

INVx5_ASAP7_75t_L g6070 ( 
.A(n_5973),
.Y(n_6070)
);

NAND2xp5_ASAP7_75t_L g6071 ( 
.A(n_5990),
.B(n_5991),
.Y(n_6071)
);

INVx2_ASAP7_75t_L g6072 ( 
.A(n_5979),
.Y(n_6072)
);

INVx2_ASAP7_75t_L g6073 ( 
.A(n_5960),
.Y(n_6073)
);

AND2x4_ASAP7_75t_L g6074 ( 
.A(n_5966),
.B(n_51),
.Y(n_6074)
);

AND2x2_ASAP7_75t_L g6075 ( 
.A(n_5974),
.B(n_52),
.Y(n_6075)
);

INVx1_ASAP7_75t_L g6076 ( 
.A(n_5999),
.Y(n_6076)
);

AND2x2_ASAP7_75t_L g6077 ( 
.A(n_5944),
.B(n_52),
.Y(n_6077)
);

NAND2xp5_ASAP7_75t_L g6078 ( 
.A(n_5968),
.B(n_52),
.Y(n_6078)
);

INVx2_ASAP7_75t_L g6079 ( 
.A(n_5976),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_6003),
.Y(n_6080)
);

NAND2xp5_ASAP7_75t_L g6081 ( 
.A(n_5995),
.B(n_53),
.Y(n_6081)
);

NAND2xp33_ASAP7_75t_R g6082 ( 
.A(n_5970),
.B(n_53),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_5977),
.Y(n_6083)
);

OR2x2_ASAP7_75t_L g6084 ( 
.A(n_6000),
.B(n_53),
.Y(n_6084)
);

AND2x2_ASAP7_75t_L g6085 ( 
.A(n_5994),
.B(n_54),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_5969),
.B(n_5972),
.Y(n_6086)
);

NOR2xp33_ASAP7_75t_L g6087 ( 
.A(n_6002),
.B(n_54),
.Y(n_6087)
);

OR2x2_ASAP7_75t_L g6088 ( 
.A(n_5996),
.B(n_54),
.Y(n_6088)
);

AND2x2_ASAP7_75t_L g6089 ( 
.A(n_5992),
.B(n_54),
.Y(n_6089)
);

AND2x2_ASAP7_75t_L g6090 ( 
.A(n_5933),
.B(n_55),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_5976),
.Y(n_6091)
);

AND2x2_ASAP7_75t_L g6092 ( 
.A(n_5987),
.B(n_55),
.Y(n_6092)
);

NAND2xp5_ASAP7_75t_SL g6093 ( 
.A(n_5980),
.B(n_55),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_5981),
.B(n_55),
.Y(n_6094)
);

OR2x2_ASAP7_75t_L g6095 ( 
.A(n_5954),
.B(n_56),
.Y(n_6095)
);

OR2x2_ASAP7_75t_L g6096 ( 
.A(n_5934),
.B(n_56),
.Y(n_6096)
);

INVx2_ASAP7_75t_L g6097 ( 
.A(n_5981),
.Y(n_6097)
);

OR2x2_ASAP7_75t_L g6098 ( 
.A(n_5929),
.B(n_56),
.Y(n_6098)
);

OR2x2_ASAP7_75t_L g6099 ( 
.A(n_5949),
.B(n_57),
.Y(n_6099)
);

AND2x2_ASAP7_75t_L g6100 ( 
.A(n_6001),
.B(n_58),
.Y(n_6100)
);

NAND2xp5_ASAP7_75t_L g6101 ( 
.A(n_6001),
.B(n_58),
.Y(n_6101)
);

OR2x2_ASAP7_75t_L g6102 ( 
.A(n_6004),
.B(n_58),
.Y(n_6102)
);

AND2x2_ASAP7_75t_L g6103 ( 
.A(n_6004),
.B(n_59),
.Y(n_6103)
);

NOR2x1_ASAP7_75t_L g6104 ( 
.A(n_5918),
.B(n_59),
.Y(n_6104)
);

INVx2_ASAP7_75t_L g6105 ( 
.A(n_5915),
.Y(n_6105)
);

INVx1_ASAP7_75t_L g6106 ( 
.A(n_5921),
.Y(n_6106)
);

INVxp67_ASAP7_75t_L g6107 ( 
.A(n_5916),
.Y(n_6107)
);

AND2x2_ASAP7_75t_L g6108 ( 
.A(n_5916),
.B(n_59),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_5921),
.Y(n_6109)
);

NAND2xp5_ASAP7_75t_L g6110 ( 
.A(n_5937),
.B(n_60),
.Y(n_6110)
);

AND2x2_ASAP7_75t_L g6111 ( 
.A(n_5916),
.B(n_60),
.Y(n_6111)
);

BUFx2_ASAP7_75t_L g6112 ( 
.A(n_5916),
.Y(n_6112)
);

INVx2_ASAP7_75t_L g6113 ( 
.A(n_5915),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_6108),
.Y(n_6114)
);

NAND2xp5_ASAP7_75t_L g6115 ( 
.A(n_6111),
.B(n_61),
.Y(n_6115)
);

AND2x2_ASAP7_75t_L g6116 ( 
.A(n_6112),
.B(n_61),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_6112),
.Y(n_6117)
);

OR2x2_ASAP7_75t_L g6118 ( 
.A(n_6019),
.B(n_61),
.Y(n_6118)
);

OR2x2_ASAP7_75t_L g6119 ( 
.A(n_6105),
.B(n_61),
.Y(n_6119)
);

INVx1_ASAP7_75t_L g6120 ( 
.A(n_6020),
.Y(n_6120)
);

AND2x2_ASAP7_75t_L g6121 ( 
.A(n_6013),
.B(n_62),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_6059),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_6113),
.Y(n_6123)
);

NAND2xp5_ASAP7_75t_L g6124 ( 
.A(n_6107),
.B(n_6015),
.Y(n_6124)
);

AND2x4_ASAP7_75t_SL g6125 ( 
.A(n_6012),
.B(n_6060),
.Y(n_6125)
);

NAND2xp5_ASAP7_75t_L g6126 ( 
.A(n_6033),
.B(n_62),
.Y(n_6126)
);

AND2x2_ASAP7_75t_L g6127 ( 
.A(n_6010),
.B(n_6008),
.Y(n_6127)
);

AND2x2_ASAP7_75t_L g6128 ( 
.A(n_6007),
.B(n_62),
.Y(n_6128)
);

A2O1A1Ixp33_ASAP7_75t_SL g6129 ( 
.A1(n_6032),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_6129)
);

OR2x2_ASAP7_75t_L g6130 ( 
.A(n_6099),
.B(n_63),
.Y(n_6130)
);

OR2x2_ASAP7_75t_L g6131 ( 
.A(n_6031),
.B(n_63),
.Y(n_6131)
);

INVx2_ASAP7_75t_L g6132 ( 
.A(n_6038),
.Y(n_6132)
);

AND2x4_ASAP7_75t_L g6133 ( 
.A(n_6007),
.B(n_63),
.Y(n_6133)
);

OR2x2_ASAP7_75t_L g6134 ( 
.A(n_6036),
.B(n_64),
.Y(n_6134)
);

NAND2xp5_ASAP7_75t_L g6135 ( 
.A(n_6033),
.B(n_65),
.Y(n_6135)
);

INVx1_ASAP7_75t_L g6136 ( 
.A(n_6035),
.Y(n_6136)
);

INVx3_ASAP7_75t_L g6137 ( 
.A(n_6024),
.Y(n_6137)
);

OR2x2_ASAP7_75t_L g6138 ( 
.A(n_6009),
.B(n_65),
.Y(n_6138)
);

OR2x2_ASAP7_75t_L g6139 ( 
.A(n_6106),
.B(n_65),
.Y(n_6139)
);

INVx2_ASAP7_75t_L g6140 ( 
.A(n_6024),
.Y(n_6140)
);

OR2x2_ASAP7_75t_L g6141 ( 
.A(n_6109),
.B(n_65),
.Y(n_6141)
);

AND2x2_ASAP7_75t_L g6142 ( 
.A(n_6060),
.B(n_66),
.Y(n_6142)
);

AOI22xp5_ASAP7_75t_L g6143 ( 
.A1(n_6025),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_6143)
);

AND2x2_ASAP7_75t_L g6144 ( 
.A(n_6070),
.B(n_66),
.Y(n_6144)
);

O2A1O1Ixp33_ASAP7_75t_L g6145 ( 
.A1(n_6044),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_6145)
);

OR2x2_ASAP7_75t_L g6146 ( 
.A(n_6034),
.B(n_67),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_6090),
.Y(n_6147)
);

AND2x2_ASAP7_75t_L g6148 ( 
.A(n_6070),
.B(n_67),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_6037),
.Y(n_6149)
);

NAND3xp33_ASAP7_75t_SL g6150 ( 
.A(n_6064),
.B(n_68),
.C(n_69),
.Y(n_6150)
);

INVxp67_ASAP7_75t_L g6151 ( 
.A(n_6082),
.Y(n_6151)
);

NAND2xp5_ASAP7_75t_L g6152 ( 
.A(n_6016),
.B(n_68),
.Y(n_6152)
);

AND2x4_ASAP7_75t_L g6153 ( 
.A(n_6072),
.B(n_69),
.Y(n_6153)
);

OR2x2_ASAP7_75t_L g6154 ( 
.A(n_6102),
.B(n_69),
.Y(n_6154)
);

AND2x4_ASAP7_75t_L g6155 ( 
.A(n_6022),
.B(n_70),
.Y(n_6155)
);

OR2x2_ASAP7_75t_L g6156 ( 
.A(n_6039),
.B(n_6047),
.Y(n_6156)
);

INVx2_ASAP7_75t_L g6157 ( 
.A(n_6048),
.Y(n_6157)
);

NAND3xp33_ASAP7_75t_L g6158 ( 
.A(n_6014),
.B(n_70),
.C(n_71),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_6052),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_6062),
.Y(n_6160)
);

NAND2xp5_ASAP7_75t_L g6161 ( 
.A(n_6017),
.B(n_70),
.Y(n_6161)
);

AND2x2_ASAP7_75t_L g6162 ( 
.A(n_6070),
.B(n_70),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_6074),
.Y(n_6163)
);

AND2x2_ASAP7_75t_L g6164 ( 
.A(n_6049),
.B(n_71),
.Y(n_6164)
);

AND2x2_ASAP7_75t_L g6165 ( 
.A(n_6055),
.B(n_71),
.Y(n_6165)
);

NAND2xp5_ASAP7_75t_L g6166 ( 
.A(n_6018),
.B(n_72),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_6074),
.Y(n_6167)
);

AND2x2_ASAP7_75t_L g6168 ( 
.A(n_6021),
.B(n_72),
.Y(n_6168)
);

NAND2xp5_ASAP7_75t_L g6169 ( 
.A(n_6050),
.B(n_72),
.Y(n_6169)
);

INVx1_ASAP7_75t_L g6170 ( 
.A(n_6110),
.Y(n_6170)
);

AND2x4_ASAP7_75t_L g6171 ( 
.A(n_6027),
.B(n_73),
.Y(n_6171)
);

AND2x2_ASAP7_75t_L g6172 ( 
.A(n_6026),
.B(n_73),
.Y(n_6172)
);

AND2x2_ASAP7_75t_L g6173 ( 
.A(n_6086),
.B(n_73),
.Y(n_6173)
);

INVx1_ASAP7_75t_L g6174 ( 
.A(n_6054),
.Y(n_6174)
);

HB1xp67_ASAP7_75t_L g6175 ( 
.A(n_6053),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_6053),
.Y(n_6176)
);

AND2x2_ASAP7_75t_L g6177 ( 
.A(n_6028),
.B(n_73),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_6014),
.Y(n_6178)
);

AOI22xp5_ASAP7_75t_L g6179 ( 
.A1(n_6065),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_6061),
.Y(n_6180)
);

INVx1_ASAP7_75t_L g6181 ( 
.A(n_6068),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_6089),
.Y(n_6182)
);

INVx2_ASAP7_75t_L g6183 ( 
.A(n_6029),
.Y(n_6183)
);

NAND2xp33_ASAP7_75t_L g6184 ( 
.A(n_6104),
.B(n_74),
.Y(n_6184)
);

AND2x2_ASAP7_75t_L g6185 ( 
.A(n_6042),
.B(n_74),
.Y(n_6185)
);

AND2x2_ASAP7_75t_L g6186 ( 
.A(n_6041),
.B(n_74),
.Y(n_6186)
);

NAND2xp5_ASAP7_75t_L g6187 ( 
.A(n_6100),
.B(n_75),
.Y(n_6187)
);

AND2x2_ASAP7_75t_L g6188 ( 
.A(n_6073),
.B(n_75),
.Y(n_6188)
);

INVx1_ASAP7_75t_L g6189 ( 
.A(n_6096),
.Y(n_6189)
);

NAND2xp5_ASAP7_75t_L g6190 ( 
.A(n_6103),
.B(n_75),
.Y(n_6190)
);

INVx2_ASAP7_75t_L g6191 ( 
.A(n_6029),
.Y(n_6191)
);

AND2x2_ASAP7_75t_L g6192 ( 
.A(n_6067),
.B(n_76),
.Y(n_6192)
);

AND2x4_ASAP7_75t_L g6193 ( 
.A(n_6076),
.B(n_76),
.Y(n_6193)
);

INVx1_ASAP7_75t_L g6194 ( 
.A(n_6098),
.Y(n_6194)
);

INVxp67_ASAP7_75t_SL g6195 ( 
.A(n_6095),
.Y(n_6195)
);

NAND2xp5_ASAP7_75t_L g6196 ( 
.A(n_6080),
.B(n_76),
.Y(n_6196)
);

OAI21xp33_ASAP7_75t_L g6197 ( 
.A1(n_6063),
.A2(n_6066),
.B(n_6023),
.Y(n_6197)
);

NAND2xp5_ASAP7_75t_L g6198 ( 
.A(n_6051),
.B(n_77),
.Y(n_6198)
);

AND2x2_ASAP7_75t_L g6199 ( 
.A(n_6083),
.B(n_77),
.Y(n_6199)
);

INVx1_ASAP7_75t_L g6200 ( 
.A(n_6075),
.Y(n_6200)
);

AND2x2_ASAP7_75t_L g6201 ( 
.A(n_6077),
.B(n_77),
.Y(n_6201)
);

INVx1_ASAP7_75t_SL g6202 ( 
.A(n_6057),
.Y(n_6202)
);

AND2x2_ASAP7_75t_L g6203 ( 
.A(n_6085),
.B(n_78),
.Y(n_6203)
);

NAND2xp5_ASAP7_75t_L g6204 ( 
.A(n_6040),
.B(n_78),
.Y(n_6204)
);

AND2x4_ASAP7_75t_SL g6205 ( 
.A(n_6092),
.B(n_79),
.Y(n_6205)
);

AND2x4_ASAP7_75t_L g6206 ( 
.A(n_6043),
.B(n_79),
.Y(n_6206)
);

INVx2_ASAP7_75t_SL g6207 ( 
.A(n_6058),
.Y(n_6207)
);

NAND2xp5_ASAP7_75t_L g6208 ( 
.A(n_6045),
.B(n_80),
.Y(n_6208)
);

AND2x2_ASAP7_75t_L g6209 ( 
.A(n_6046),
.B(n_80),
.Y(n_6209)
);

NAND2xp5_ASAP7_75t_L g6210 ( 
.A(n_6087),
.B(n_80),
.Y(n_6210)
);

AND2x2_ASAP7_75t_L g6211 ( 
.A(n_6011),
.B(n_81),
.Y(n_6211)
);

INVx2_ASAP7_75t_L g6212 ( 
.A(n_6084),
.Y(n_6212)
);

NAND2x1_ASAP7_75t_L g6213 ( 
.A(n_6030),
.B(n_81),
.Y(n_6213)
);

INVx1_ASAP7_75t_L g6214 ( 
.A(n_6071),
.Y(n_6214)
);

INVx1_ASAP7_75t_L g6215 ( 
.A(n_6088),
.Y(n_6215)
);

INVxp67_ASAP7_75t_L g6216 ( 
.A(n_6116),
.Y(n_6216)
);

INVx1_ASAP7_75t_L g6217 ( 
.A(n_6142),
.Y(n_6217)
);

HB1xp67_ASAP7_75t_L g6218 ( 
.A(n_6120),
.Y(n_6218)
);

INVx1_ASAP7_75t_L g6219 ( 
.A(n_6144),
.Y(n_6219)
);

AND2x2_ASAP7_75t_L g6220 ( 
.A(n_6125),
.B(n_6127),
.Y(n_6220)
);

INVxp67_ASAP7_75t_L g6221 ( 
.A(n_6148),
.Y(n_6221)
);

INVx1_ASAP7_75t_L g6222 ( 
.A(n_6162),
.Y(n_6222)
);

OR2x2_ASAP7_75t_L g6223 ( 
.A(n_6132),
.B(n_6094),
.Y(n_6223)
);

INVx2_ASAP7_75t_L g6224 ( 
.A(n_6137),
.Y(n_6224)
);

AND2x2_ASAP7_75t_L g6225 ( 
.A(n_6121),
.B(n_6093),
.Y(n_6225)
);

NAND2xp5_ASAP7_75t_L g6226 ( 
.A(n_6153),
.B(n_6056),
.Y(n_6226)
);

INVx1_ASAP7_75t_L g6227 ( 
.A(n_6168),
.Y(n_6227)
);

INVx2_ASAP7_75t_L g6228 ( 
.A(n_6156),
.Y(n_6228)
);

INVx1_ASAP7_75t_L g6229 ( 
.A(n_6128),
.Y(n_6229)
);

INVx1_ASAP7_75t_SL g6230 ( 
.A(n_6119),
.Y(n_6230)
);

AND2x2_ASAP7_75t_L g6231 ( 
.A(n_6173),
.B(n_6078),
.Y(n_6231)
);

AND2x2_ASAP7_75t_L g6232 ( 
.A(n_6172),
.B(n_6209),
.Y(n_6232)
);

OR2x2_ASAP7_75t_L g6233 ( 
.A(n_6124),
.B(n_6117),
.Y(n_6233)
);

NAND2xp5_ASAP7_75t_L g6234 ( 
.A(n_6202),
.B(n_6101),
.Y(n_6234)
);

INVx1_ASAP7_75t_SL g6235 ( 
.A(n_6133),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_6126),
.Y(n_6236)
);

NAND4xp25_ASAP7_75t_L g6237 ( 
.A(n_6151),
.B(n_6069),
.C(n_6091),
.D(n_6079),
.Y(n_6237)
);

AND2x4_ASAP7_75t_L g6238 ( 
.A(n_6140),
.B(n_6097),
.Y(n_6238)
);

INVx1_ASAP7_75t_L g6239 ( 
.A(n_6135),
.Y(n_6239)
);

OR2x2_ASAP7_75t_L g6240 ( 
.A(n_6130),
.B(n_6081),
.Y(n_6240)
);

BUFx2_ASAP7_75t_L g6241 ( 
.A(n_6155),
.Y(n_6241)
);

OR2x2_ASAP7_75t_L g6242 ( 
.A(n_6204),
.B(n_81),
.Y(n_6242)
);

AND2x2_ASAP7_75t_L g6243 ( 
.A(n_6177),
.B(n_81),
.Y(n_6243)
);

INVx2_ASAP7_75t_L g6244 ( 
.A(n_6171),
.Y(n_6244)
);

AND2x2_ASAP7_75t_L g6245 ( 
.A(n_6185),
.B(n_82),
.Y(n_6245)
);

NAND2xp33_ASAP7_75t_L g6246 ( 
.A(n_6157),
.B(n_82),
.Y(n_6246)
);

NAND2xp5_ASAP7_75t_L g6247 ( 
.A(n_6155),
.B(n_82),
.Y(n_6247)
);

OAI22xp33_ASAP7_75t_L g6248 ( 
.A1(n_6131),
.A2(n_82),
.B1(n_777),
.B2(n_776),
.Y(n_6248)
);

NAND2xp5_ASAP7_75t_L g6249 ( 
.A(n_6205),
.B(n_777),
.Y(n_6249)
);

INVx1_ASAP7_75t_L g6250 ( 
.A(n_6188),
.Y(n_6250)
);

NAND2xp5_ASAP7_75t_L g6251 ( 
.A(n_6211),
.B(n_778),
.Y(n_6251)
);

INVxp67_ASAP7_75t_SL g6252 ( 
.A(n_6175),
.Y(n_6252)
);

NAND2xp5_ASAP7_75t_L g6253 ( 
.A(n_6171),
.B(n_778),
.Y(n_6253)
);

INVx2_ASAP7_75t_L g6254 ( 
.A(n_6183),
.Y(n_6254)
);

NAND2xp5_ASAP7_75t_L g6255 ( 
.A(n_6206),
.B(n_6186),
.Y(n_6255)
);

OR2x2_ASAP7_75t_L g6256 ( 
.A(n_6166),
.B(n_779),
.Y(n_6256)
);

AND2x2_ASAP7_75t_L g6257 ( 
.A(n_6192),
.B(n_779),
.Y(n_6257)
);

AND2x2_ASAP7_75t_L g6258 ( 
.A(n_6199),
.B(n_779),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_6123),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_6206),
.Y(n_6260)
);

AOI22xp5_ASAP7_75t_L g6261 ( 
.A1(n_6184),
.A2(n_782),
.B1(n_780),
.B2(n_781),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_6134),
.Y(n_6262)
);

INVx2_ASAP7_75t_SL g6263 ( 
.A(n_6191),
.Y(n_6263)
);

NAND2x1p5_ASAP7_75t_L g6264 ( 
.A(n_6193),
.B(n_780),
.Y(n_6264)
);

INVx2_ASAP7_75t_L g6265 ( 
.A(n_6149),
.Y(n_6265)
);

NOR2xp33_ASAP7_75t_SL g6266 ( 
.A(n_6163),
.B(n_780),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_6118),
.Y(n_6267)
);

INVx2_ASAP7_75t_SL g6268 ( 
.A(n_6159),
.Y(n_6268)
);

INVxp67_ASAP7_75t_L g6269 ( 
.A(n_6164),
.Y(n_6269)
);

NAND2x1p5_ASAP7_75t_L g6270 ( 
.A(n_6193),
.B(n_781),
.Y(n_6270)
);

OAI22xp33_ASAP7_75t_L g6271 ( 
.A1(n_6213),
.A2(n_784),
.B1(n_782),
.B2(n_783),
.Y(n_6271)
);

NAND2xp5_ASAP7_75t_L g6272 ( 
.A(n_6165),
.B(n_784),
.Y(n_6272)
);

NOR2xp33_ASAP7_75t_SL g6273 ( 
.A(n_6167),
.B(n_6160),
.Y(n_6273)
);

HB1xp67_ASAP7_75t_L g6274 ( 
.A(n_6136),
.Y(n_6274)
);

NAND2xp5_ASAP7_75t_L g6275 ( 
.A(n_6129),
.B(n_785),
.Y(n_6275)
);

INVx1_ASAP7_75t_L g6276 ( 
.A(n_6201),
.Y(n_6276)
);

AND2x4_ASAP7_75t_L g6277 ( 
.A(n_6207),
.B(n_785),
.Y(n_6277)
);

AND2x4_ASAP7_75t_L g6278 ( 
.A(n_6212),
.B(n_785),
.Y(n_6278)
);

AND2x2_ASAP7_75t_L g6279 ( 
.A(n_6114),
.B(n_786),
.Y(n_6279)
);

INVx2_ASAP7_75t_L g6280 ( 
.A(n_6203),
.Y(n_6280)
);

NAND2xp33_ASAP7_75t_L g6281 ( 
.A(n_6154),
.B(n_786),
.Y(n_6281)
);

AND2x2_ASAP7_75t_L g6282 ( 
.A(n_6180),
.B(n_787),
.Y(n_6282)
);

INVx2_ASAP7_75t_SL g6283 ( 
.A(n_6146),
.Y(n_6283)
);

NAND2xp5_ASAP7_75t_L g6284 ( 
.A(n_6195),
.B(n_787),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_6115),
.Y(n_6285)
);

A2O1A1Ixp33_ASAP7_75t_L g6286 ( 
.A1(n_6197),
.A2(n_789),
.B(n_787),
.C(n_788),
.Y(n_6286)
);

OR2x2_ASAP7_75t_L g6287 ( 
.A(n_6208),
.B(n_788),
.Y(n_6287)
);

CKINVDCx14_ASAP7_75t_R g6288 ( 
.A(n_6150),
.Y(n_6288)
);

INVx2_ASAP7_75t_L g6289 ( 
.A(n_6138),
.Y(n_6289)
);

INVx1_ASAP7_75t_L g6290 ( 
.A(n_6187),
.Y(n_6290)
);

INVx1_ASAP7_75t_SL g6291 ( 
.A(n_6139),
.Y(n_6291)
);

AND2x2_ASAP7_75t_L g6292 ( 
.A(n_6181),
.B(n_788),
.Y(n_6292)
);

AND2x2_ASAP7_75t_L g6293 ( 
.A(n_6200),
.B(n_790),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_6190),
.Y(n_6294)
);

AOI211xp5_ASAP7_75t_SL g6295 ( 
.A1(n_6174),
.A2(n_792),
.B(n_790),
.C(n_791),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_6141),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_6152),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_6161),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_6169),
.Y(n_6299)
);

INVx1_ASAP7_75t_SL g6300 ( 
.A(n_6210),
.Y(n_6300)
);

INVx1_ASAP7_75t_SL g6301 ( 
.A(n_6189),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_6147),
.Y(n_6302)
);

INVx1_ASAP7_75t_L g6303 ( 
.A(n_6158),
.Y(n_6303)
);

AND2x2_ASAP7_75t_L g6304 ( 
.A(n_6182),
.B(n_790),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_6178),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_6176),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_6198),
.Y(n_6307)
);

OR2x6_ASAP7_75t_L g6308 ( 
.A(n_6145),
.B(n_791),
.Y(n_6308)
);

OR2x2_ASAP7_75t_L g6309 ( 
.A(n_6196),
.B(n_791),
.Y(n_6309)
);

INVx2_ASAP7_75t_L g6310 ( 
.A(n_6194),
.Y(n_6310)
);

INVx2_ASAP7_75t_L g6311 ( 
.A(n_6215),
.Y(n_6311)
);

INVx2_ASAP7_75t_SL g6312 ( 
.A(n_6170),
.Y(n_6312)
);

OAI22xp5_ASAP7_75t_L g6313 ( 
.A1(n_6288),
.A2(n_6214),
.B1(n_6143),
.B2(n_6122),
.Y(n_6313)
);

AOI21xp33_ASAP7_75t_L g6314 ( 
.A1(n_6220),
.A2(n_6179),
.B(n_793),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_6241),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_6247),
.Y(n_6316)
);

INVx1_ASAP7_75t_L g6317 ( 
.A(n_6228),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6253),
.Y(n_6318)
);

XOR2x2_ASAP7_75t_L g6319 ( 
.A(n_6226),
.B(n_793),
.Y(n_6319)
);

OAI21xp33_ASAP7_75t_L g6320 ( 
.A1(n_6273),
.A2(n_793),
.B(n_794),
.Y(n_6320)
);

AOI22xp5_ASAP7_75t_L g6321 ( 
.A1(n_6263),
.A2(n_6224),
.B1(n_6235),
.B2(n_6243),
.Y(n_6321)
);

AOI22xp5_ASAP7_75t_L g6322 ( 
.A1(n_6245),
.A2(n_796),
.B1(n_794),
.B2(n_795),
.Y(n_6322)
);

AOI22xp5_ASAP7_75t_L g6323 ( 
.A1(n_6266),
.A2(n_6246),
.B1(n_6254),
.B2(n_6244),
.Y(n_6323)
);

INVx2_ASAP7_75t_L g6324 ( 
.A(n_6238),
.Y(n_6324)
);

OAI22xp33_ASAP7_75t_L g6325 ( 
.A1(n_6308),
.A2(n_797),
.B1(n_795),
.B2(n_796),
.Y(n_6325)
);

AOI22xp5_ASAP7_75t_L g6326 ( 
.A1(n_6232),
.A2(n_797),
.B1(n_795),
.B2(n_796),
.Y(n_6326)
);

XNOR2xp5_ASAP7_75t_L g6327 ( 
.A(n_6261),
.B(n_798),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_6218),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_6264),
.Y(n_6329)
);

INVx2_ASAP7_75t_L g6330 ( 
.A(n_6238),
.Y(n_6330)
);

NAND3xp33_ASAP7_75t_L g6331 ( 
.A(n_6286),
.B(n_798),
.C(n_799),
.Y(n_6331)
);

INVx1_ASAP7_75t_SL g6332 ( 
.A(n_6278),
.Y(n_6332)
);

OAI21xp33_ASAP7_75t_L g6333 ( 
.A1(n_6233),
.A2(n_798),
.B(n_799),
.Y(n_6333)
);

AOI22xp5_ASAP7_75t_L g6334 ( 
.A1(n_6279),
.A2(n_6282),
.B1(n_6293),
.B2(n_6292),
.Y(n_6334)
);

INVx1_ASAP7_75t_L g6335 ( 
.A(n_6270),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_L g6336 ( 
.A(n_6257),
.B(n_800),
.Y(n_6336)
);

INVx2_ASAP7_75t_L g6337 ( 
.A(n_6268),
.Y(n_6337)
);

NAND2xp5_ASAP7_75t_L g6338 ( 
.A(n_6295),
.B(n_800),
.Y(n_6338)
);

INVx1_ASAP7_75t_L g6339 ( 
.A(n_6277),
.Y(n_6339)
);

XOR2x2_ASAP7_75t_L g6340 ( 
.A(n_6255),
.B(n_801),
.Y(n_6340)
);

AOI22xp5_ASAP7_75t_L g6341 ( 
.A1(n_6304),
.A2(n_803),
.B1(n_801),
.B2(n_802),
.Y(n_6341)
);

NOR2xp33_ASAP7_75t_L g6342 ( 
.A(n_6216),
.B(n_801),
.Y(n_6342)
);

NOR2xp33_ASAP7_75t_L g6343 ( 
.A(n_6221),
.B(n_802),
.Y(n_6343)
);

AOI22xp5_ASAP7_75t_L g6344 ( 
.A1(n_6225),
.A2(n_804),
.B1(n_802),
.B2(n_803),
.Y(n_6344)
);

INVx1_ASAP7_75t_L g6345 ( 
.A(n_6277),
.Y(n_6345)
);

NOR2x1_ASAP7_75t_SL g6346 ( 
.A(n_6265),
.B(n_804),
.Y(n_6346)
);

OAI21xp5_ASAP7_75t_L g6347 ( 
.A1(n_6269),
.A2(n_804),
.B(n_805),
.Y(n_6347)
);

NAND2xp5_ASAP7_75t_L g6348 ( 
.A(n_6258),
.B(n_805),
.Y(n_6348)
);

OAI22xp33_ASAP7_75t_L g6349 ( 
.A1(n_6308),
.A2(n_807),
.B1(n_805),
.B2(n_806),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_6249),
.Y(n_6350)
);

AOI22xp5_ASAP7_75t_L g6351 ( 
.A1(n_6301),
.A2(n_809),
.B1(n_807),
.B2(n_808),
.Y(n_6351)
);

AOI21xp33_ASAP7_75t_SL g6352 ( 
.A1(n_6271),
.A2(n_1067),
.B(n_807),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_6278),
.Y(n_6353)
);

HB1xp67_ASAP7_75t_L g6354 ( 
.A(n_6274),
.Y(n_6354)
);

AOI22x1_ASAP7_75t_SL g6355 ( 
.A1(n_6303),
.A2(n_810),
.B1(n_808),
.B2(n_809),
.Y(n_6355)
);

O2A1O1Ixp33_ASAP7_75t_SL g6356 ( 
.A1(n_6284),
.A2(n_6234),
.B(n_6219),
.C(n_6222),
.Y(n_6356)
);

XNOR2x1_ASAP7_75t_SL g6357 ( 
.A(n_6312),
.B(n_808),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_6252),
.Y(n_6358)
);

NAND3xp33_ASAP7_75t_SL g6359 ( 
.A(n_6300),
.B(n_809),
.C(n_810),
.Y(n_6359)
);

NOR2xp33_ASAP7_75t_R g6360 ( 
.A(n_6260),
.B(n_810),
.Y(n_6360)
);

INVx1_ASAP7_75t_SL g6361 ( 
.A(n_6223),
.Y(n_6361)
);

AOI21xp33_ASAP7_75t_L g6362 ( 
.A1(n_6259),
.A2(n_811),
.B(n_813),
.Y(n_6362)
);

OAI22xp5_ASAP7_75t_L g6363 ( 
.A1(n_6217),
.A2(n_814),
.B1(n_811),
.B2(n_813),
.Y(n_6363)
);

OAI21xp33_ASAP7_75t_L g6364 ( 
.A1(n_6227),
.A2(n_811),
.B(n_813),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_6272),
.Y(n_6365)
);

OAI22xp5_ASAP7_75t_L g6366 ( 
.A1(n_6276),
.A2(n_6291),
.B1(n_6242),
.B2(n_6230),
.Y(n_6366)
);

AOI211x1_ASAP7_75t_L g6367 ( 
.A1(n_6237),
.A2(n_816),
.B(n_814),
.C(n_815),
.Y(n_6367)
);

AOI21xp5_ASAP7_75t_L g6368 ( 
.A1(n_6281),
.A2(n_6275),
.B(n_6251),
.Y(n_6368)
);

OR2x2_ASAP7_75t_L g6369 ( 
.A(n_6256),
.B(n_815),
.Y(n_6369)
);

OAI21xp5_ASAP7_75t_L g6370 ( 
.A1(n_6250),
.A2(n_816),
.B(n_817),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_6287),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_6280),
.Y(n_6372)
);

INVx2_ASAP7_75t_L g6373 ( 
.A(n_6310),
.Y(n_6373)
);

OAI21xp33_ASAP7_75t_L g6374 ( 
.A1(n_6262),
.A2(n_6283),
.B(n_6296),
.Y(n_6374)
);

OAI21xp5_ASAP7_75t_L g6375 ( 
.A1(n_6229),
.A2(n_6267),
.B(n_6302),
.Y(n_6375)
);

AOI22xp5_ASAP7_75t_L g6376 ( 
.A1(n_6231),
.A2(n_818),
.B1(n_816),
.B2(n_817),
.Y(n_6376)
);

AOI21xp33_ASAP7_75t_L g6377 ( 
.A1(n_6311),
.A2(n_817),
.B(n_818),
.Y(n_6377)
);

OAI21xp33_ASAP7_75t_L g6378 ( 
.A1(n_6289),
.A2(n_818),
.B(n_819),
.Y(n_6378)
);

INVx1_ASAP7_75t_L g6379 ( 
.A(n_6324),
.Y(n_6379)
);

AOI21xp5_ASAP7_75t_L g6380 ( 
.A1(n_6338),
.A2(n_6348),
.B(n_6336),
.Y(n_6380)
);

AOI211xp5_ASAP7_75t_L g6381 ( 
.A1(n_6314),
.A2(n_6248),
.B(n_6307),
.C(n_6298),
.Y(n_6381)
);

OAI31xp33_ASAP7_75t_L g6382 ( 
.A1(n_6357),
.A2(n_6297),
.A3(n_6239),
.B(n_6236),
.Y(n_6382)
);

OAI22xp5_ASAP7_75t_L g6383 ( 
.A1(n_6321),
.A2(n_6240),
.B1(n_6309),
.B2(n_6285),
.Y(n_6383)
);

NAND3xp33_ASAP7_75t_L g6384 ( 
.A(n_6317),
.B(n_6306),
.C(n_6305),
.Y(n_6384)
);

OAI22xp5_ASAP7_75t_L g6385 ( 
.A1(n_6323),
.A2(n_6294),
.B1(n_6290),
.B2(n_6299),
.Y(n_6385)
);

AOI221xp5_ASAP7_75t_L g6386 ( 
.A1(n_6367),
.A2(n_821),
.B1(n_819),
.B2(n_820),
.C(n_822),
.Y(n_6386)
);

OAI21xp33_ASAP7_75t_L g6387 ( 
.A1(n_6315),
.A2(n_819),
.B(n_820),
.Y(n_6387)
);

OAI22xp5_ASAP7_75t_L g6388 ( 
.A1(n_6330),
.A2(n_823),
.B1(n_821),
.B2(n_822),
.Y(n_6388)
);

NAND2xp5_ASAP7_75t_L g6389 ( 
.A(n_6332),
.B(n_821),
.Y(n_6389)
);

AND2x2_ASAP7_75t_L g6390 ( 
.A(n_6337),
.B(n_822),
.Y(n_6390)
);

NAND2xp5_ASAP7_75t_L g6391 ( 
.A(n_6358),
.B(n_823),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6346),
.Y(n_6392)
);

NAND2xp5_ASAP7_75t_L g6393 ( 
.A(n_6339),
.B(n_823),
.Y(n_6393)
);

AND2x2_ASAP7_75t_L g6394 ( 
.A(n_6361),
.B(n_824),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_6354),
.Y(n_6395)
);

INVxp67_ASAP7_75t_L g6396 ( 
.A(n_6343),
.Y(n_6396)
);

OAI211xp5_ASAP7_75t_SL g6397 ( 
.A1(n_6374),
.A2(n_826),
.B(n_824),
.C(n_825),
.Y(n_6397)
);

OAI332xp33_ASAP7_75t_L g6398 ( 
.A1(n_6313),
.A2(n_824),
.A3(n_825),
.B1(n_826),
.B2(n_827),
.B3(n_828),
.C1(n_829),
.C2(n_830),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_6345),
.Y(n_6399)
);

NAND2xp5_ASAP7_75t_L g6400 ( 
.A(n_6325),
.B(n_825),
.Y(n_6400)
);

OAI21xp33_ASAP7_75t_L g6401 ( 
.A1(n_6319),
.A2(n_827),
.B(n_828),
.Y(n_6401)
);

NOR4xp25_ASAP7_75t_L g6402 ( 
.A(n_6328),
.B(n_829),
.C(n_827),
.D(n_828),
.Y(n_6402)
);

OR2x2_ASAP7_75t_L g6403 ( 
.A(n_6353),
.B(n_829),
.Y(n_6403)
);

INVx2_ASAP7_75t_SL g6404 ( 
.A(n_6373),
.Y(n_6404)
);

NAND2xp5_ASAP7_75t_L g6405 ( 
.A(n_6349),
.B(n_830),
.Y(n_6405)
);

OAI22xp33_ASAP7_75t_SL g6406 ( 
.A1(n_6369),
.A2(n_832),
.B1(n_830),
.B2(n_831),
.Y(n_6406)
);

INVxp67_ASAP7_75t_L g6407 ( 
.A(n_6342),
.Y(n_6407)
);

AOI22xp5_ASAP7_75t_L g6408 ( 
.A1(n_6372),
.A2(n_833),
.B1(n_831),
.B2(n_832),
.Y(n_6408)
);

INVx2_ASAP7_75t_L g6409 ( 
.A(n_6329),
.Y(n_6409)
);

INVx2_ASAP7_75t_L g6410 ( 
.A(n_6335),
.Y(n_6410)
);

AOI22xp5_ASAP7_75t_L g6411 ( 
.A1(n_6359),
.A2(n_834),
.B1(n_831),
.B2(n_833),
.Y(n_6411)
);

AOI22xp5_ASAP7_75t_L g6412 ( 
.A1(n_6320),
.A2(n_835),
.B1(n_833),
.B2(n_834),
.Y(n_6412)
);

INVxp67_ASAP7_75t_L g6413 ( 
.A(n_6355),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_6351),
.Y(n_6414)
);

NAND2xp5_ASAP7_75t_L g6415 ( 
.A(n_6352),
.B(n_835),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_6327),
.Y(n_6416)
);

AOI22xp33_ASAP7_75t_L g6417 ( 
.A1(n_6331),
.A2(n_1062),
.B1(n_837),
.B2(n_835),
.Y(n_6417)
);

OAI31xp33_ASAP7_75t_L g6418 ( 
.A1(n_6333),
.A2(n_838),
.A3(n_836),
.B(n_837),
.Y(n_6418)
);

AOI22xp5_ASAP7_75t_L g6419 ( 
.A1(n_6366),
.A2(n_838),
.B1(n_836),
.B2(n_837),
.Y(n_6419)
);

NAND2xp5_ASAP7_75t_SL g6420 ( 
.A(n_6352),
.B(n_836),
.Y(n_6420)
);

NAND2xp5_ASAP7_75t_L g6421 ( 
.A(n_6334),
.B(n_838),
.Y(n_6421)
);

AOI321xp33_ASAP7_75t_L g6422 ( 
.A1(n_6318),
.A2(n_841),
.A3(n_843),
.B1(n_839),
.B2(n_840),
.C(n_842),
.Y(n_6422)
);

INVx1_ASAP7_75t_SL g6423 ( 
.A(n_6360),
.Y(n_6423)
);

BUFx2_ASAP7_75t_L g6424 ( 
.A(n_6370),
.Y(n_6424)
);

XNOR2xp5_ASAP7_75t_L g6425 ( 
.A(n_6340),
.B(n_839),
.Y(n_6425)
);

OAI22xp5_ASAP7_75t_L g6426 ( 
.A1(n_6344),
.A2(n_841),
.B1(n_839),
.B2(n_840),
.Y(n_6426)
);

NAND2xp5_ASAP7_75t_L g6427 ( 
.A(n_6341),
.B(n_840),
.Y(n_6427)
);

OAI322xp33_ASAP7_75t_L g6428 ( 
.A1(n_6371),
.A2(n_841),
.A3(n_842),
.B1(n_843),
.B2(n_844),
.C1(n_845),
.C2(n_846),
.Y(n_6428)
);

INVx1_ASAP7_75t_L g6429 ( 
.A(n_6363),
.Y(n_6429)
);

AOI21xp33_ASAP7_75t_L g6430 ( 
.A1(n_6378),
.A2(n_842),
.B(n_843),
.Y(n_6430)
);

INVxp67_ASAP7_75t_SL g6431 ( 
.A(n_6326),
.Y(n_6431)
);

OAI22xp5_ASAP7_75t_L g6432 ( 
.A1(n_6376),
.A2(n_846),
.B1(n_844),
.B2(n_845),
.Y(n_6432)
);

INVx1_ASAP7_75t_L g6433 ( 
.A(n_6364),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_6322),
.Y(n_6434)
);

NOR2xp33_ASAP7_75t_L g6435 ( 
.A(n_6377),
.B(n_845),
.Y(n_6435)
);

AOI22xp5_ASAP7_75t_L g6436 ( 
.A1(n_6316),
.A2(n_848),
.B1(n_846),
.B2(n_847),
.Y(n_6436)
);

HB1xp67_ASAP7_75t_L g6437 ( 
.A(n_6375),
.Y(n_6437)
);

NAND2xp5_ASAP7_75t_L g6438 ( 
.A(n_6368),
.B(n_847),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6347),
.Y(n_6439)
);

AND2x2_ASAP7_75t_L g6440 ( 
.A(n_6350),
.B(n_847),
.Y(n_6440)
);

AOI21xp5_ASAP7_75t_L g6441 ( 
.A1(n_6356),
.A2(n_848),
.B(n_849),
.Y(n_6441)
);

OR2x2_ASAP7_75t_L g6442 ( 
.A(n_6365),
.B(n_848),
.Y(n_6442)
);

AOI21xp5_ASAP7_75t_L g6443 ( 
.A1(n_6362),
.A2(n_849),
.B(n_850),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_6392),
.Y(n_6444)
);

INVx1_ASAP7_75t_SL g6445 ( 
.A(n_6379),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6390),
.Y(n_6446)
);

AOI22xp5_ASAP7_75t_L g6447 ( 
.A1(n_6413),
.A2(n_852),
.B1(n_850),
.B2(n_851),
.Y(n_6447)
);

OR2x2_ASAP7_75t_L g6448 ( 
.A(n_6404),
.B(n_850),
.Y(n_6448)
);

OAI322xp33_ASAP7_75t_L g6449 ( 
.A1(n_6395),
.A2(n_851),
.A3(n_852),
.B1(n_853),
.B2(n_855),
.C1(n_856),
.C2(n_857),
.Y(n_6449)
);

OR2x2_ASAP7_75t_L g6450 ( 
.A(n_6403),
.B(n_6389),
.Y(n_6450)
);

AOI22xp5_ASAP7_75t_L g6451 ( 
.A1(n_6409),
.A2(n_853),
.B1(n_851),
.B2(n_852),
.Y(n_6451)
);

AOI211xp5_ASAP7_75t_L g6452 ( 
.A1(n_6430),
.A2(n_857),
.B(n_855),
.C(n_856),
.Y(n_6452)
);

OAI322xp33_ASAP7_75t_L g6453 ( 
.A1(n_6410),
.A2(n_856),
.A3(n_857),
.B1(n_858),
.B2(n_859),
.C1(n_860),
.C2(n_861),
.Y(n_6453)
);

OAI22xp5_ASAP7_75t_L g6454 ( 
.A1(n_6419),
.A2(n_860),
.B1(n_858),
.B2(n_859),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_6394),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6393),
.Y(n_6456)
);

INVxp67_ASAP7_75t_L g6457 ( 
.A(n_6420),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_6400),
.Y(n_6458)
);

AOI22xp5_ASAP7_75t_L g6459 ( 
.A1(n_6401),
.A2(n_860),
.B1(n_858),
.B2(n_859),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_6405),
.Y(n_6460)
);

OAI332xp33_ASAP7_75t_L g6461 ( 
.A1(n_6423),
.A2(n_861),
.A3(n_862),
.B1(n_863),
.B2(n_864),
.B3(n_865),
.C1(n_866),
.C2(n_867),
.Y(n_6461)
);

AND2x2_ASAP7_75t_L g6462 ( 
.A(n_6440),
.B(n_861),
.Y(n_6462)
);

NAND2xp5_ASAP7_75t_L g6463 ( 
.A(n_6441),
.B(n_862),
.Y(n_6463)
);

AOI22xp5_ASAP7_75t_L g6464 ( 
.A1(n_6414),
.A2(n_864),
.B1(n_862),
.B2(n_863),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_6438),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_6391),
.Y(n_6466)
);

OAI22xp5_ASAP7_75t_L g6467 ( 
.A1(n_6425),
.A2(n_867),
.B1(n_865),
.B2(n_866),
.Y(n_6467)
);

OAI33xp33_ASAP7_75t_L g6468 ( 
.A1(n_6383),
.A2(n_867),
.A3(n_868),
.B1(n_869),
.B2(n_870),
.B3(n_871),
.Y(n_6468)
);

AOI31xp33_ASAP7_75t_L g6469 ( 
.A1(n_6386),
.A2(n_870),
.A3(n_868),
.B(n_869),
.Y(n_6469)
);

AOI22xp5_ASAP7_75t_L g6470 ( 
.A1(n_6435),
.A2(n_871),
.B1(n_868),
.B2(n_870),
.Y(n_6470)
);

OAI32xp33_ASAP7_75t_L g6471 ( 
.A1(n_6442),
.A2(n_874),
.A3(n_872),
.B1(n_873),
.B2(n_875),
.Y(n_6471)
);

NAND2xp5_ASAP7_75t_L g6472 ( 
.A(n_6402),
.B(n_872),
.Y(n_6472)
);

NAND2xp5_ASAP7_75t_L g6473 ( 
.A(n_6411),
.B(n_6382),
.Y(n_6473)
);

OAI322xp33_ASAP7_75t_L g6474 ( 
.A1(n_6433),
.A2(n_873),
.A3(n_874),
.B1(n_875),
.B2(n_876),
.C1(n_877),
.C2(n_878),
.Y(n_6474)
);

INVx1_ASAP7_75t_L g6475 ( 
.A(n_6415),
.Y(n_6475)
);

OAI32xp33_ASAP7_75t_L g6476 ( 
.A1(n_6429),
.A2(n_876),
.A3(n_873),
.B1(n_874),
.B2(n_877),
.Y(n_6476)
);

AOI21xp33_ASAP7_75t_L g6477 ( 
.A1(n_6406),
.A2(n_1062),
.B(n_878),
.Y(n_6477)
);

INVx2_ASAP7_75t_SL g6478 ( 
.A(n_6399),
.Y(n_6478)
);

OAI21xp5_ASAP7_75t_L g6479 ( 
.A1(n_6443),
.A2(n_879),
.B(n_880),
.Y(n_6479)
);

NOR3xp33_ASAP7_75t_SL g6480 ( 
.A(n_6397),
.B(n_1061),
.C(n_879),
.Y(n_6480)
);

NAND2xp5_ASAP7_75t_L g6481 ( 
.A(n_6411),
.B(n_879),
.Y(n_6481)
);

INVx1_ASAP7_75t_L g6482 ( 
.A(n_6388),
.Y(n_6482)
);

NAND2xp5_ASAP7_75t_L g6483 ( 
.A(n_6417),
.B(n_880),
.Y(n_6483)
);

INVx2_ASAP7_75t_SL g6484 ( 
.A(n_6421),
.Y(n_6484)
);

AOI22xp5_ASAP7_75t_L g6485 ( 
.A1(n_6431),
.A2(n_883),
.B1(n_881),
.B2(n_882),
.Y(n_6485)
);

OAI321xp33_ASAP7_75t_L g6486 ( 
.A1(n_6385),
.A2(n_882),
.A3(n_883),
.B1(n_884),
.B2(n_885),
.C(n_886),
.Y(n_6486)
);

CKINVDCx16_ASAP7_75t_R g6487 ( 
.A(n_6412),
.Y(n_6487)
);

AOI322xp5_ASAP7_75t_L g6488 ( 
.A1(n_6434),
.A2(n_6416),
.A3(n_6439),
.B1(n_6437),
.B2(n_6396),
.C1(n_6407),
.C2(n_6424),
.Y(n_6488)
);

NOR2xp33_ASAP7_75t_L g6489 ( 
.A(n_6468),
.B(n_6398),
.Y(n_6489)
);

OAI21xp33_ASAP7_75t_L g6490 ( 
.A1(n_6473),
.A2(n_6387),
.B(n_6427),
.Y(n_6490)
);

NOR2xp33_ASAP7_75t_L g6491 ( 
.A(n_6444),
.B(n_6384),
.Y(n_6491)
);

AOI22xp5_ASAP7_75t_SL g6492 ( 
.A1(n_6463),
.A2(n_6426),
.B1(n_6432),
.B2(n_6380),
.Y(n_6492)
);

AOI21xp33_ASAP7_75t_SL g6493 ( 
.A1(n_6469),
.A2(n_6418),
.B(n_6408),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_6448),
.Y(n_6494)
);

AND2x2_ASAP7_75t_L g6495 ( 
.A(n_6445),
.B(n_6381),
.Y(n_6495)
);

OA22x2_ASAP7_75t_L g6496 ( 
.A1(n_6464),
.A2(n_6436),
.B1(n_6422),
.B2(n_6428),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_6481),
.Y(n_6497)
);

NAND2xp5_ASAP7_75t_SL g6498 ( 
.A(n_6487),
.B(n_882),
.Y(n_6498)
);

NOR2x1_ASAP7_75t_L g6499 ( 
.A(n_6465),
.B(n_883),
.Y(n_6499)
);

NAND2xp5_ASAP7_75t_L g6500 ( 
.A(n_6462),
.B(n_884),
.Y(n_6500)
);

NAND2x1_ASAP7_75t_L g6501 ( 
.A(n_6478),
.B(n_884),
.Y(n_6501)
);

INVx1_ASAP7_75t_L g6502 ( 
.A(n_6483),
.Y(n_6502)
);

NOR3xp33_ASAP7_75t_L g6503 ( 
.A(n_6461),
.B(n_885),
.C(n_886),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_6447),
.Y(n_6504)
);

OAI21xp5_ASAP7_75t_SL g6505 ( 
.A1(n_6459),
.A2(n_885),
.B(n_886),
.Y(n_6505)
);

AOI21xp33_ASAP7_75t_L g6506 ( 
.A1(n_6476),
.A2(n_887),
.B(n_888),
.Y(n_6506)
);

INVx1_ASAP7_75t_SL g6507 ( 
.A(n_6450),
.Y(n_6507)
);

AOI221xp5_ASAP7_75t_L g6508 ( 
.A1(n_6471),
.A2(n_889),
.B1(n_887),
.B2(n_888),
.C(n_890),
.Y(n_6508)
);

XNOR2xp5_ASAP7_75t_L g6509 ( 
.A(n_6480),
.B(n_887),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_6453),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_6474),
.Y(n_6511)
);

NAND3xp33_ASAP7_75t_L g6512 ( 
.A(n_6488),
.B(n_888),
.C(n_889),
.Y(n_6512)
);

AOI211xp5_ASAP7_75t_L g6513 ( 
.A1(n_6477),
.A2(n_891),
.B(n_889),
.C(n_890),
.Y(n_6513)
);

NAND3xp33_ASAP7_75t_L g6514 ( 
.A(n_6485),
.B(n_890),
.C(n_891),
.Y(n_6514)
);

AOI221xp5_ASAP7_75t_L g6515 ( 
.A1(n_6486),
.A2(n_893),
.B1(n_891),
.B2(n_892),
.C(n_894),
.Y(n_6515)
);

NOR2xp33_ASAP7_75t_L g6516 ( 
.A(n_6472),
.B(n_892),
.Y(n_6516)
);

AND2x2_ASAP7_75t_L g6517 ( 
.A(n_6455),
.B(n_892),
.Y(n_6517)
);

AOI211xp5_ASAP7_75t_L g6518 ( 
.A1(n_6449),
.A2(n_895),
.B(n_893),
.C(n_894),
.Y(n_6518)
);

AND2x2_ASAP7_75t_L g6519 ( 
.A(n_6446),
.B(n_893),
.Y(n_6519)
);

INVx2_ASAP7_75t_L g6520 ( 
.A(n_6482),
.Y(n_6520)
);

AOI211x1_ASAP7_75t_L g6521 ( 
.A1(n_6479),
.A2(n_897),
.B(n_895),
.C(n_896),
.Y(n_6521)
);

NAND2x1p5_ASAP7_75t_L g6522 ( 
.A(n_6470),
.B(n_896),
.Y(n_6522)
);

NAND2xp5_ASAP7_75t_L g6523 ( 
.A(n_6451),
.B(n_896),
.Y(n_6523)
);

AND2x2_ASAP7_75t_L g6524 ( 
.A(n_6457),
.B(n_897),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_6454),
.Y(n_6525)
);

INVx1_ASAP7_75t_SL g6526 ( 
.A(n_6458),
.Y(n_6526)
);

NOR3x1_ASAP7_75t_L g6527 ( 
.A(n_6467),
.B(n_897),
.C(n_898),
.Y(n_6527)
);

OAI211xp5_ASAP7_75t_SL g6528 ( 
.A1(n_6452),
.A2(n_900),
.B(n_898),
.C(n_899),
.Y(n_6528)
);

NOR4xp25_ASAP7_75t_L g6529 ( 
.A(n_6460),
.B(n_6475),
.C(n_6466),
.D(n_6484),
.Y(n_6529)
);

OAI21xp5_ASAP7_75t_L g6530 ( 
.A1(n_6456),
.A2(n_898),
.B(n_899),
.Y(n_6530)
);

AOI21xp5_ASAP7_75t_L g6531 ( 
.A1(n_6476),
.A2(n_900),
.B(n_901),
.Y(n_6531)
);

NAND2xp5_ASAP7_75t_SL g6532 ( 
.A(n_6444),
.B(n_900),
.Y(n_6532)
);

AOI21xp5_ASAP7_75t_L g6533 ( 
.A1(n_6476),
.A2(n_901),
.B(n_902),
.Y(n_6533)
);

NAND2xp5_ASAP7_75t_L g6534 ( 
.A(n_6444),
.B(n_902),
.Y(n_6534)
);

OAI211xp5_ASAP7_75t_L g6535 ( 
.A1(n_6464),
.A2(n_904),
.B(n_902),
.C(n_903),
.Y(n_6535)
);

INVx2_ASAP7_75t_L g6536 ( 
.A(n_6444),
.Y(n_6536)
);

AND2x4_ASAP7_75t_L g6537 ( 
.A(n_6536),
.B(n_903),
.Y(n_6537)
);

AOI211xp5_ASAP7_75t_L g6538 ( 
.A1(n_6506),
.A2(n_905),
.B(n_903),
.C(n_904),
.Y(n_6538)
);

AOI22xp5_ASAP7_75t_L g6539 ( 
.A1(n_6503),
.A2(n_1059),
.B1(n_906),
.B2(n_904),
.Y(n_6539)
);

NOR3x1_ASAP7_75t_L g6540 ( 
.A(n_6512),
.B(n_905),
.C(n_906),
.Y(n_6540)
);

NAND2xp5_ASAP7_75t_SL g6541 ( 
.A(n_6511),
.B(n_906),
.Y(n_6541)
);

AOI22xp33_ASAP7_75t_L g6542 ( 
.A1(n_6510),
.A2(n_909),
.B1(n_907),
.B2(n_908),
.Y(n_6542)
);

NOR2xp33_ASAP7_75t_L g6543 ( 
.A(n_6520),
.B(n_907),
.Y(n_6543)
);

AOI211xp5_ASAP7_75t_L g6544 ( 
.A1(n_6493),
.A2(n_909),
.B(n_907),
.C(n_908),
.Y(n_6544)
);

NAND4xp25_ASAP7_75t_L g6545 ( 
.A(n_6489),
.B(n_912),
.C(n_910),
.D(n_911),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_6524),
.B(n_6517),
.Y(n_6546)
);

OAI221xp5_ASAP7_75t_L g6547 ( 
.A1(n_6505),
.A2(n_910),
.B1(n_911),
.B2(n_912),
.C(n_913),
.Y(n_6547)
);

O2A1O1Ixp5_ASAP7_75t_SL g6548 ( 
.A1(n_6498),
.A2(n_913),
.B(n_910),
.C(n_912),
.Y(n_6548)
);

AOI21xp5_ASAP7_75t_L g6549 ( 
.A1(n_6531),
.A2(n_913),
.B(n_914),
.Y(n_6549)
);

INVx1_ASAP7_75t_L g6550 ( 
.A(n_6501),
.Y(n_6550)
);

AOI211xp5_ASAP7_75t_L g6551 ( 
.A1(n_6528),
.A2(n_916),
.B(n_914),
.C(n_915),
.Y(n_6551)
);

NAND2xp5_ASAP7_75t_L g6552 ( 
.A(n_6519),
.B(n_914),
.Y(n_6552)
);

OAI22xp5_ASAP7_75t_L g6553 ( 
.A1(n_6509),
.A2(n_917),
.B1(n_915),
.B2(n_916),
.Y(n_6553)
);

AOI221xp5_ASAP7_75t_L g6554 ( 
.A1(n_6491),
.A2(n_915),
.B1(n_916),
.B2(n_917),
.C(n_918),
.Y(n_6554)
);

AOI221xp5_ASAP7_75t_SL g6555 ( 
.A1(n_6490),
.A2(n_6515),
.B1(n_6533),
.B2(n_6507),
.C(n_6518),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_6495),
.Y(n_6556)
);

O2A1O1Ixp33_ASAP7_75t_L g6557 ( 
.A1(n_6532),
.A2(n_920),
.B(n_918),
.C(n_919),
.Y(n_6557)
);

INVx2_ASAP7_75t_SL g6558 ( 
.A(n_6494),
.Y(n_6558)
);

AOI21xp5_ASAP7_75t_L g6559 ( 
.A1(n_6500),
.A2(n_918),
.B(n_920),
.Y(n_6559)
);

AOI22xp5_ASAP7_75t_L g6560 ( 
.A1(n_6516),
.A2(n_1059),
.B1(n_922),
.B2(n_920),
.Y(n_6560)
);

HB1xp67_ASAP7_75t_L g6561 ( 
.A(n_6499),
.Y(n_6561)
);

NAND3xp33_ASAP7_75t_SL g6562 ( 
.A(n_6513),
.B(n_921),
.C(n_922),
.Y(n_6562)
);

NAND2xp5_ASAP7_75t_L g6563 ( 
.A(n_6537),
.B(n_6542),
.Y(n_6563)
);

OAI221xp5_ASAP7_75t_L g6564 ( 
.A1(n_6539),
.A2(n_6508),
.B1(n_6530),
.B2(n_6534),
.C(n_6535),
.Y(n_6564)
);

AOI221xp5_ASAP7_75t_L g6565 ( 
.A1(n_6553),
.A2(n_6529),
.B1(n_6521),
.B2(n_6514),
.C(n_6504),
.Y(n_6565)
);

NOR2xp33_ASAP7_75t_L g6566 ( 
.A(n_6545),
.B(n_6526),
.Y(n_6566)
);

NOR3x1_ASAP7_75t_L g6567 ( 
.A(n_6547),
.B(n_6523),
.C(n_6525),
.Y(n_6567)
);

OAI221xp5_ASAP7_75t_L g6568 ( 
.A1(n_6554),
.A2(n_6522),
.B1(n_6497),
.B2(n_6502),
.C(n_6492),
.Y(n_6568)
);

NAND2xp5_ASAP7_75t_SL g6569 ( 
.A(n_6544),
.B(n_6496),
.Y(n_6569)
);

AOI21xp5_ASAP7_75t_L g6570 ( 
.A1(n_6541),
.A2(n_6499),
.B(n_6527),
.Y(n_6570)
);

AND2x2_ASAP7_75t_L g6571 ( 
.A(n_6556),
.B(n_921),
.Y(n_6571)
);

AOI211xp5_ASAP7_75t_L g6572 ( 
.A1(n_6562),
.A2(n_6543),
.B(n_6549),
.C(n_6557),
.Y(n_6572)
);

NAND4xp25_ASAP7_75t_SL g6573 ( 
.A(n_6555),
.B(n_924),
.C(n_922),
.D(n_923),
.Y(n_6573)
);

AOI22xp5_ASAP7_75t_L g6574 ( 
.A1(n_6558),
.A2(n_926),
.B1(n_923),
.B2(n_925),
.Y(n_6574)
);

AOI21xp33_ASAP7_75t_SL g6575 ( 
.A1(n_6552),
.A2(n_923),
.B(n_925),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6537),
.Y(n_6576)
);

OAI211xp5_ASAP7_75t_L g6577 ( 
.A1(n_6538),
.A2(n_6551),
.B(n_6560),
.C(n_6559),
.Y(n_6577)
);

OAI222xp33_ASAP7_75t_L g6578 ( 
.A1(n_6550),
.A2(n_6546),
.B1(n_6561),
.B2(n_6540),
.C1(n_6548),
.C2(n_929),
.Y(n_6578)
);

AOI221xp5_ASAP7_75t_L g6579 ( 
.A1(n_6553),
.A2(n_925),
.B1(n_926),
.B2(n_927),
.C(n_928),
.Y(n_6579)
);

AOI322xp5_ASAP7_75t_L g6580 ( 
.A1(n_6542),
.A2(n_926),
.A3(n_927),
.B1(n_928),
.B2(n_929),
.C1(n_930),
.C2(n_931),
.Y(n_6580)
);

AOI21xp33_ASAP7_75t_L g6581 ( 
.A1(n_6557),
.A2(n_927),
.B(n_929),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_6537),
.Y(n_6582)
);

AND3x1_ASAP7_75t_L g6583 ( 
.A(n_6544),
.B(n_930),
.C(n_931),
.Y(n_6583)
);

OAI21xp5_ASAP7_75t_L g6584 ( 
.A1(n_6549),
.A2(n_930),
.B(n_931),
.Y(n_6584)
);

O2A1O1Ixp33_ASAP7_75t_L g6585 ( 
.A1(n_6541),
.A2(n_934),
.B(n_932),
.C(n_933),
.Y(n_6585)
);

NAND4xp75_ASAP7_75t_L g6586 ( 
.A(n_6540),
.B(n_934),
.C(n_932),
.D(n_933),
.Y(n_6586)
);

NOR2xp33_ASAP7_75t_L g6587 ( 
.A(n_6573),
.B(n_932),
.Y(n_6587)
);

NOR2xp33_ASAP7_75t_L g6588 ( 
.A(n_6578),
.B(n_933),
.Y(n_6588)
);

AOI21xp33_ASAP7_75t_SL g6589 ( 
.A1(n_6569),
.A2(n_6568),
.B(n_6566),
.Y(n_6589)
);

INVx1_ASAP7_75t_L g6590 ( 
.A(n_6571),
.Y(n_6590)
);

OAI211xp5_ASAP7_75t_L g6591 ( 
.A1(n_6565),
.A2(n_936),
.B(n_934),
.C(n_935),
.Y(n_6591)
);

OAI211xp5_ASAP7_75t_L g6592 ( 
.A1(n_6581),
.A2(n_937),
.B(n_935),
.C(n_936),
.Y(n_6592)
);

AOI211xp5_ASAP7_75t_L g6593 ( 
.A1(n_6575),
.A2(n_938),
.B(n_935),
.C(n_937),
.Y(n_6593)
);

NAND4xp25_ASAP7_75t_L g6594 ( 
.A(n_6567),
.B(n_6572),
.C(n_6579),
.D(n_6580),
.Y(n_6594)
);

AOI222xp33_ASAP7_75t_L g6595 ( 
.A1(n_6584),
.A2(n_6576),
.B1(n_6582),
.B2(n_6564),
.C1(n_6563),
.C2(n_6577),
.Y(n_6595)
);

NOR3xp33_ASAP7_75t_L g6596 ( 
.A(n_6585),
.B(n_1056),
.C(n_937),
.Y(n_6596)
);

O2A1O1Ixp33_ASAP7_75t_L g6597 ( 
.A1(n_6570),
.A2(n_942),
.B(n_938),
.C(n_941),
.Y(n_6597)
);

INVxp33_ASAP7_75t_L g6598 ( 
.A(n_6586),
.Y(n_6598)
);

NOR2x1_ASAP7_75t_L g6599 ( 
.A(n_6583),
.B(n_938),
.Y(n_6599)
);

NAND3xp33_ASAP7_75t_SL g6600 ( 
.A(n_6574),
.B(n_941),
.C(n_943),
.Y(n_6600)
);

OAI221xp5_ASAP7_75t_SL g6601 ( 
.A1(n_6580),
.A2(n_941),
.B1(n_943),
.B2(n_944),
.C(n_945),
.Y(n_6601)
);

OAI211xp5_ASAP7_75t_L g6602 ( 
.A1(n_6565),
.A2(n_946),
.B(n_944),
.C(n_945),
.Y(n_6602)
);

OAI22xp5_ASAP7_75t_L g6603 ( 
.A1(n_6568),
.A2(n_946),
.B1(n_944),
.B2(n_945),
.Y(n_6603)
);

INVx1_ASAP7_75t_L g6604 ( 
.A(n_6571),
.Y(n_6604)
);

NOR2xp33_ASAP7_75t_R g6605 ( 
.A(n_6573),
.B(n_946),
.Y(n_6605)
);

INVxp67_ASAP7_75t_L g6606 ( 
.A(n_6571),
.Y(n_6606)
);

NOR2x1p5_ASAP7_75t_L g6607 ( 
.A(n_6594),
.B(n_947),
.Y(n_6607)
);

INVxp33_ASAP7_75t_L g6608 ( 
.A(n_6605),
.Y(n_6608)
);

XNOR2x1_ASAP7_75t_L g6609 ( 
.A(n_6599),
.B(n_947),
.Y(n_6609)
);

NOR3xp33_ASAP7_75t_L g6610 ( 
.A(n_6591),
.B(n_948),
.C(n_949),
.Y(n_6610)
);

NAND2xp5_ASAP7_75t_L g6611 ( 
.A(n_6588),
.B(n_948),
.Y(n_6611)
);

NAND4xp75_ASAP7_75t_L g6612 ( 
.A(n_6587),
.B(n_6590),
.C(n_6604),
.D(n_6589),
.Y(n_6612)
);

NOR2x1_ASAP7_75t_L g6613 ( 
.A(n_6602),
.B(n_949),
.Y(n_6613)
);

INVx2_ASAP7_75t_SL g6614 ( 
.A(n_6603),
.Y(n_6614)
);

NOR2x1_ASAP7_75t_L g6615 ( 
.A(n_6600),
.B(n_6592),
.Y(n_6615)
);

NAND3xp33_ASAP7_75t_SL g6616 ( 
.A(n_6595),
.B(n_950),
.C(n_951),
.Y(n_6616)
);

NOR2xp67_ASAP7_75t_L g6617 ( 
.A(n_6606),
.B(n_950),
.Y(n_6617)
);

INVx1_ASAP7_75t_L g6618 ( 
.A(n_6597),
.Y(n_6618)
);

AOI22xp5_ASAP7_75t_L g6619 ( 
.A1(n_6596),
.A2(n_952),
.B1(n_950),
.B2(n_951),
.Y(n_6619)
);

NOR2x1_ASAP7_75t_L g6620 ( 
.A(n_6598),
.B(n_6601),
.Y(n_6620)
);

NOR2x1_ASAP7_75t_SL g6621 ( 
.A(n_6593),
.B(n_951),
.Y(n_6621)
);

NOR3xp33_ASAP7_75t_L g6622 ( 
.A(n_6591),
.B(n_952),
.C(n_953),
.Y(n_6622)
);

NAND2xp5_ASAP7_75t_L g6623 ( 
.A(n_6588),
.B(n_1056),
.Y(n_6623)
);

NOR3xp33_ASAP7_75t_L g6624 ( 
.A(n_6591),
.B(n_952),
.C(n_954),
.Y(n_6624)
);

INVx2_ASAP7_75t_L g6625 ( 
.A(n_6590),
.Y(n_6625)
);

NAND4xp75_ASAP7_75t_L g6626 ( 
.A(n_6599),
.B(n_956),
.C(n_954),
.D(n_955),
.Y(n_6626)
);

NAND2xp5_ASAP7_75t_L g6627 ( 
.A(n_6617),
.B(n_6610),
.Y(n_6627)
);

NOR3x2_ASAP7_75t_L g6628 ( 
.A(n_6612),
.B(n_1056),
.C(n_955),
.Y(n_6628)
);

NOR3xp33_ASAP7_75t_L g6629 ( 
.A(n_6616),
.B(n_955),
.C(n_956),
.Y(n_6629)
);

NOR2x1_ASAP7_75t_L g6630 ( 
.A(n_6607),
.B(n_957),
.Y(n_6630)
);

NOR2xp33_ASAP7_75t_L g6631 ( 
.A(n_6608),
.B(n_957),
.Y(n_6631)
);

NOR2xp67_ASAP7_75t_L g6632 ( 
.A(n_6618),
.B(n_957),
.Y(n_6632)
);

NOR2x1_ASAP7_75t_L g6633 ( 
.A(n_6626),
.B(n_958),
.Y(n_6633)
);

AND2x2_ASAP7_75t_L g6634 ( 
.A(n_6625),
.B(n_958),
.Y(n_6634)
);

NOR2x1p5_ASAP7_75t_L g6635 ( 
.A(n_6611),
.B(n_959),
.Y(n_6635)
);

OAI22xp5_ASAP7_75t_L g6636 ( 
.A1(n_6623),
.A2(n_961),
.B1(n_959),
.B2(n_960),
.Y(n_6636)
);

NOR2x1_ASAP7_75t_L g6637 ( 
.A(n_6613),
.B(n_959),
.Y(n_6637)
);

NOR2x1_ASAP7_75t_L g6638 ( 
.A(n_6620),
.B(n_960),
.Y(n_6638)
);

NOR2x1_ASAP7_75t_L g6639 ( 
.A(n_6609),
.B(n_960),
.Y(n_6639)
);

NAND4xp75_ASAP7_75t_L g6640 ( 
.A(n_6615),
.B(n_963),
.C(n_961),
.D(n_962),
.Y(n_6640)
);

INVx1_ASAP7_75t_L g6641 ( 
.A(n_6619),
.Y(n_6641)
);

NOR3x2_ASAP7_75t_L g6642 ( 
.A(n_6621),
.B(n_961),
.C(n_962),
.Y(n_6642)
);

CKINVDCx5p33_ASAP7_75t_R g6643 ( 
.A(n_6614),
.Y(n_6643)
);

NOR3xp33_ASAP7_75t_L g6644 ( 
.A(n_6622),
.B(n_963),
.C(n_964),
.Y(n_6644)
);

NOR2x1_ASAP7_75t_L g6645 ( 
.A(n_6624),
.B(n_964),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6611),
.Y(n_6646)
);

NOR3x2_ASAP7_75t_L g6647 ( 
.A(n_6612),
.B(n_1055),
.C(n_964),
.Y(n_6647)
);

AND2x4_ASAP7_75t_L g6648 ( 
.A(n_6625),
.B(n_965),
.Y(n_6648)
);

NAND2xp5_ASAP7_75t_L g6649 ( 
.A(n_6617),
.B(n_965),
.Y(n_6649)
);

XNOR2x1_ASAP7_75t_L g6650 ( 
.A(n_6643),
.B(n_6639),
.Y(n_6650)
);

AND2x4_ASAP7_75t_L g6651 ( 
.A(n_6634),
.B(n_966),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_6628),
.Y(n_6652)
);

AND2x4_ASAP7_75t_L g6653 ( 
.A(n_6646),
.B(n_966),
.Y(n_6653)
);

OAI22xp5_ASAP7_75t_L g6654 ( 
.A1(n_6649),
.A2(n_969),
.B1(n_967),
.B2(n_968),
.Y(n_6654)
);

AND2x2_ASAP7_75t_L g6655 ( 
.A(n_6648),
.B(n_6630),
.Y(n_6655)
);

NAND2x1p5_ASAP7_75t_L g6656 ( 
.A(n_6641),
.B(n_967),
.Y(n_6656)
);

AOI221xp5_ASAP7_75t_L g6657 ( 
.A1(n_6636),
.A2(n_1055),
.B1(n_969),
.B2(n_970),
.C(n_971),
.Y(n_6657)
);

NAND2x1p5_ASAP7_75t_L g6658 ( 
.A(n_6648),
.B(n_968),
.Y(n_6658)
);

AND3x2_ASAP7_75t_L g6659 ( 
.A(n_6644),
.B(n_968),
.C(n_970),
.Y(n_6659)
);

INVx1_ASAP7_75t_L g6660 ( 
.A(n_6647),
.Y(n_6660)
);

HB1xp67_ASAP7_75t_L g6661 ( 
.A(n_6632),
.Y(n_6661)
);

INVx1_ASAP7_75t_L g6662 ( 
.A(n_6640),
.Y(n_6662)
);

NOR4xp25_ASAP7_75t_L g6663 ( 
.A(n_6627),
.B(n_970),
.C(n_971),
.D(n_972),
.Y(n_6663)
);

NOR2xp33_ASAP7_75t_L g6664 ( 
.A(n_6650),
.B(n_6631),
.Y(n_6664)
);

XNOR2xp5_ASAP7_75t_L g6665 ( 
.A(n_6651),
.B(n_6642),
.Y(n_6665)
);

NAND3xp33_ASAP7_75t_SL g6666 ( 
.A(n_6657),
.B(n_6629),
.C(n_6635),
.Y(n_6666)
);

NOR2xp33_ASAP7_75t_R g6667 ( 
.A(n_6659),
.B(n_6645),
.Y(n_6667)
);

NAND2xp33_ASAP7_75t_SL g6668 ( 
.A(n_6655),
.B(n_6637),
.Y(n_6668)
);

XOR2xp5_ASAP7_75t_L g6669 ( 
.A(n_6654),
.B(n_6638),
.Y(n_6669)
);

NAND2xp33_ASAP7_75t_SL g6670 ( 
.A(n_6652),
.B(n_6633),
.Y(n_6670)
);

NAND2xp33_ASAP7_75t_SL g6671 ( 
.A(n_6660),
.B(n_971),
.Y(n_6671)
);

NOR2xp33_ASAP7_75t_R g6672 ( 
.A(n_6662),
.B(n_1055),
.Y(n_6672)
);

OAI21xp5_ASAP7_75t_SL g6673 ( 
.A1(n_6653),
.A2(n_972),
.B(n_974),
.Y(n_6673)
);

NAND2xp33_ASAP7_75t_SL g6674 ( 
.A(n_6661),
.B(n_972),
.Y(n_6674)
);

INVx1_ASAP7_75t_L g6675 ( 
.A(n_6672),
.Y(n_6675)
);

NOR2x1_ASAP7_75t_L g6676 ( 
.A(n_6666),
.B(n_6658),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_6671),
.Y(n_6677)
);

INVx1_ASAP7_75t_L g6678 ( 
.A(n_6673),
.Y(n_6678)
);

INVx1_ASAP7_75t_L g6679 ( 
.A(n_6674),
.Y(n_6679)
);

OAI22x1_ASAP7_75t_L g6680 ( 
.A1(n_6676),
.A2(n_6664),
.B1(n_6665),
.B2(n_6669),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_6675),
.Y(n_6681)
);

INVx2_ASAP7_75t_L g6682 ( 
.A(n_6678),
.Y(n_6682)
);

INVx1_ASAP7_75t_L g6683 ( 
.A(n_6677),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6680),
.Y(n_6684)
);

HB1xp67_ASAP7_75t_L g6685 ( 
.A(n_6682),
.Y(n_6685)
);

INVx2_ASAP7_75t_L g6686 ( 
.A(n_6684),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_6686),
.Y(n_6687)
);

INVxp67_ASAP7_75t_L g6688 ( 
.A(n_6687),
.Y(n_6688)
);

NAND2xp5_ASAP7_75t_L g6689 ( 
.A(n_6688),
.B(n_6683),
.Y(n_6689)
);

AOI21x1_ASAP7_75t_L g6690 ( 
.A1(n_6689),
.A2(n_6685),
.B(n_6681),
.Y(n_6690)
);

AND4x1_ASAP7_75t_L g6691 ( 
.A(n_6690),
.B(n_6670),
.C(n_6668),
.D(n_6679),
.Y(n_6691)
);

AOI22xp33_ASAP7_75t_L g6692 ( 
.A1(n_6691),
.A2(n_6667),
.B1(n_6656),
.B2(n_6663),
.Y(n_6692)
);

XNOR2xp5_ASAP7_75t_L g6693 ( 
.A(n_6692),
.B(n_975),
.Y(n_6693)
);

O2A1O1Ixp33_ASAP7_75t_L g6694 ( 
.A1(n_6693),
.A2(n_975),
.B(n_976),
.C(n_977),
.Y(n_6694)
);

AOI211xp5_ASAP7_75t_L g6695 ( 
.A1(n_6694),
.A2(n_976),
.B(n_977),
.C(n_978),
.Y(n_6695)
);


endmodule