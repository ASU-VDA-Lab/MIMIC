module fake_jpeg_2209_n_200 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_200);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_27),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_60),
.Y(n_89)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_0),
.B(n_1),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_84),
.A2(n_64),
.B1(n_67),
.B2(n_56),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_70),
.B1(n_3),
.B2(n_5),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_67),
.B(n_69),
.C(n_65),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_68),
.B(n_66),
.C(n_59),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_99),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_52),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_52),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_58),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_65),
.C(n_63),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_114),
.Y(n_121)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_7),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_53),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_107),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2x1p5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_83),
.B1(n_76),
.B2(n_74),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_118),
.B1(n_119),
.B2(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_74),
.B1(n_66),
.B2(n_68),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_116),
.B1(n_88),
.B2(n_91),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_62),
.B(n_69),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_5),
.C(n_6),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_57),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_2),
.B(n_3),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_18),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_107),
.B1(n_109),
.B2(n_115),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_28),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_140),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_91),
.B1(n_93),
.B2(n_8),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_131),
.B1(n_11),
.B2(n_12),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_6),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_8),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_10),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_157),
.B1(n_50),
.B2(n_45),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_118),
.B(n_31),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_165),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_29),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_163),
.Y(n_166)
);

AOI21x1_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_32),
.B(n_49),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_162),
.B(n_39),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_164),
.B1(n_126),
.B2(n_127),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_14),
.B(n_16),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_14),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_161),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_R g161 ( 
.A(n_142),
.B(n_19),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_20),
.A3(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_26),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_36),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_40),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_123),
.B1(n_126),
.B2(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_168),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_160),
.B1(n_145),
.B2(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_175),
.B(n_177),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_148),
.B(n_41),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_179),
.B(n_151),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_46),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_186),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_170),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_189),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_163),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_190),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_167),
.B1(n_168),
.B2(n_174),
.Y(n_191)
);

AOI31xp67_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_183),
.A3(n_180),
.B(n_172),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_188),
.B(n_155),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_196),
.B(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_169),
.B(n_159),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_164),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_153),
.Y(n_200)
);


endmodule