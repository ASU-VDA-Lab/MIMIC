module real_aes_1608_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_810, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_810;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g208 ( .A(n_0), .B(n_130), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_1), .B(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_2), .B(n_136), .Y(n_149) );
INVx1_ASAP7_75t_L g123 ( .A(n_3), .Y(n_123) );
NAND2xp33_ASAP7_75t_SL g200 ( .A(n_4), .B(n_134), .Y(n_200) );
INVx1_ASAP7_75t_L g181 ( .A(n_5), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_6), .B(n_154), .Y(n_527) );
INVx1_ASAP7_75t_L g507 ( .A(n_7), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g779 ( .A(n_8), .Y(n_779) );
AND2x2_ASAP7_75t_L g147 ( .A(n_9), .B(n_140), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_10), .Y(n_474) );
INVx2_ASAP7_75t_L g141 ( .A(n_11), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_12), .Y(n_760) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_13), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_13), .B(n_27), .Y(n_703) );
INVx1_ASAP7_75t_L g535 ( .A(n_14), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g790 ( .A1(n_15), .A2(n_27), .B1(n_757), .B2(n_791), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_15), .Y(n_791) );
AOI221x1_ASAP7_75t_L g194 ( .A1(n_16), .A2(n_118), .B1(n_195), .B2(n_197), .C(n_199), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_17), .B(n_136), .Y(n_169) );
INVx1_ASAP7_75t_L g766 ( .A(n_18), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_19), .B(n_786), .Y(n_797) );
INVx1_ASAP7_75t_L g533 ( .A(n_20), .Y(n_533) );
INVx1_ASAP7_75t_SL g456 ( .A(n_21), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_22), .B(n_137), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_23), .A2(n_118), .B(n_151), .Y(n_150) );
AOI221xp5_ASAP7_75t_SL g161 ( .A1(n_24), .A2(n_40), .B1(n_118), .B2(n_136), .C(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_25), .B(n_130), .Y(n_152) );
AOI33xp33_ASAP7_75t_L g493 ( .A1(n_26), .A2(n_52), .A3(n_184), .B1(n_190), .B2(n_494), .B3(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g757 ( .A(n_27), .Y(n_757) );
INVx1_ASAP7_75t_L g467 ( .A(n_28), .Y(n_467) );
OR2x2_ASAP7_75t_L g142 ( .A(n_29), .B(n_89), .Y(n_142) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_29), .A2(n_89), .B(n_141), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_30), .B(n_126), .Y(n_173) );
INVxp67_ASAP7_75t_L g193 ( .A(n_31), .Y(n_193) );
AND2x2_ASAP7_75t_L g224 ( .A(n_32), .B(n_139), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_33), .B(n_182), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_34), .A2(n_118), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_35), .B(n_126), .Y(n_163) );
AND2x2_ASAP7_75t_L g119 ( .A(n_36), .B(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g134 ( .A(n_36), .B(n_123), .Y(n_134) );
INVx1_ASAP7_75t_L g189 ( .A(n_36), .Y(n_189) );
OR2x6_ASAP7_75t_L g764 ( .A(n_37), .B(n_765), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_38), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_39), .B(n_182), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_41), .A2(n_154), .B1(n_198), .B2(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_42), .B(n_525), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_43), .A2(n_81), .B1(n_118), .B2(n_187), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_44), .B(n_137), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_45), .B(n_130), .Y(n_222) );
AOI222xp33_ASAP7_75t_L g101 ( .A1(n_46), .A2(n_102), .B1(n_772), .B2(n_783), .C1(n_798), .C2(n_800), .Y(n_101) );
XNOR2xp5_ASAP7_75t_L g787 ( .A(n_46), .B(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_47), .B(n_174), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_48), .B(n_137), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_49), .Y(n_520) );
AND2x2_ASAP7_75t_L g211 ( .A(n_50), .B(n_139), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_51), .B(n_139), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_53), .B(n_137), .Y(n_485) );
INVx1_ASAP7_75t_L g122 ( .A(n_54), .Y(n_122) );
INVx1_ASAP7_75t_L g132 ( .A(n_54), .Y(n_132) );
AND2x2_ASAP7_75t_L g486 ( .A(n_55), .B(n_139), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g505 ( .A1(n_56), .A2(n_74), .B1(n_182), .B2(n_187), .C(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_57), .B(n_182), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_58), .B(n_136), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_59), .B(n_198), .Y(n_476) );
AOI21xp5_ASAP7_75t_SL g445 ( .A1(n_60), .A2(n_187), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g143 ( .A(n_61), .B(n_139), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_62), .B(n_126), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_63), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_64), .B(n_140), .Y(n_176) );
INVx1_ASAP7_75t_L g530 ( .A(n_65), .Y(n_530) );
XNOR2xp5_ASAP7_75t_L g759 ( .A(n_66), .B(n_760), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_67), .A2(n_118), .B(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g484 ( .A(n_68), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_69), .B(n_126), .Y(n_153) );
AND2x2_ASAP7_75t_SL g261 ( .A(n_70), .B(n_174), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_71), .A2(n_187), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g120 ( .A(n_72), .Y(n_120) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_73), .B(n_182), .Y(n_496) );
AND2x2_ASAP7_75t_L g458 ( .A(n_75), .B(n_197), .Y(n_458) );
INVx1_ASAP7_75t_L g531 ( .A(n_76), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_77), .A2(n_187), .B(n_455), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_78), .A2(n_187), .B(n_257), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_79), .B(n_136), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_80), .A2(n_84), .B1(n_136), .B2(n_182), .Y(n_259) );
INVx1_ASAP7_75t_L g767 ( .A(n_82), .Y(n_767) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_83), .B(n_197), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_85), .A2(n_187), .B1(n_491), .B2(n_492), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_86), .B(n_130), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_87), .B(n_130), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g117 ( .A1(n_88), .A2(n_118), .B(n_124), .Y(n_117) );
INVx1_ASAP7_75t_L g447 ( .A(n_90), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_91), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g497 ( .A(n_92), .B(n_197), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_93), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_94), .A2(n_465), .B(n_466), .C(n_468), .Y(n_464) );
INVxp67_ASAP7_75t_L g196 ( .A(n_95), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_96), .B(n_136), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_97), .B(n_126), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_98), .A2(n_118), .B(n_171), .Y(n_170) );
BUFx2_ASAP7_75t_L g780 ( .A(n_99), .Y(n_780) );
BUFx2_ASAP7_75t_SL g806 ( .A(n_99), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_100), .B(n_137), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_763), .B1(n_768), .B2(n_769), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_759), .B1(n_761), .B2(n_762), .Y(n_103) );
INVx1_ASAP7_75t_L g761 ( .A(n_104), .Y(n_761) );
OAI21x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_107), .B(n_433), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g758 ( .A(n_106), .Y(n_758) );
OR2x2_ASAP7_75t_L g771 ( .A(n_106), .B(n_764), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_106), .B(n_763), .Y(n_782) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_372), .Y(n_107) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_109), .B(n_265), .C(n_316), .Y(n_108) );
OAI211xp5_ASAP7_75t_SL g109 ( .A1(n_110), .A2(n_155), .B(n_212), .C(n_243), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_144), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_114), .B(n_217), .Y(n_380) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g225 ( .A(n_115), .B(n_146), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_115), .B(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g242 ( .A(n_115), .B(n_232), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_115), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g279 ( .A(n_115), .B(n_255), .Y(n_279) );
INVx2_ASAP7_75t_L g305 ( .A(n_115), .Y(n_305) );
AND2x4_ASAP7_75t_L g314 ( .A(n_115), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g419 ( .A(n_115), .B(n_286), .Y(n_419) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_138), .B(n_143), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_135), .Y(n_116) );
AND2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
BUFx3_ASAP7_75t_L g186 ( .A(n_119), .Y(n_186) );
AND2x6_ASAP7_75t_L g130 ( .A(n_120), .B(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g191 ( .A(n_120), .Y(n_191) );
AND2x4_ASAP7_75t_L g187 ( .A(n_121), .B(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AND2x4_ASAP7_75t_L g126 ( .A(n_122), .B(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g184 ( .A(n_122), .Y(n_184) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_123), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_129), .B(n_133), .Y(n_124) );
INVxp67_ASAP7_75t_L g536 ( .A(n_126), .Y(n_536) );
AND2x4_ASAP7_75t_L g137 ( .A(n_127), .B(n_131), .Y(n_137) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVxp67_ASAP7_75t_L g534 ( .A(n_130), .Y(n_534) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_133), .A2(n_152), .B(n_153), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_133), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_133), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_133), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_133), .A2(n_221), .B(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_133), .A2(n_447), .B(n_448), .C(n_449), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_SL g455 ( .A1(n_133), .A2(n_448), .B(n_456), .C(n_457), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_133), .A2(n_448), .B(n_484), .C(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g491 ( .A(n_133), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g506 ( .A1(n_133), .A2(n_448), .B(n_507), .C(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_133), .A2(n_523), .B(n_524), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_133), .B(n_154), .Y(n_537) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g136 ( .A(n_134), .B(n_137), .Y(n_136) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_134), .Y(n_468) );
INVx1_ASAP7_75t_L g201 ( .A(n_137), .Y(n_201) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_138), .A2(n_218), .B(n_224), .Y(n_217) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_138), .A2(n_218), .B(n_224), .Y(n_232) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_138), .A2(n_452), .B(n_458), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_139), .Y(n_138) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_139), .A2(n_161), .B(n_165), .Y(n_160) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x4_ASAP7_75t_L g154 ( .A(n_141), .B(n_142), .Y(n_154) );
AND2x2_ASAP7_75t_L g303 ( .A(n_144), .B(n_304), .Y(n_303) );
OAI32xp33_ASAP7_75t_L g386 ( .A1(n_144), .A2(n_308), .A3(n_312), .B1(n_319), .B2(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_144), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g240 ( .A(n_145), .B(n_241), .Y(n_240) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_145), .B(n_235), .C(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g339 ( .A(n_145), .B(n_242), .Y(n_339) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_146), .Y(n_229) );
INVx5_ASAP7_75t_L g264 ( .A(n_146), .Y(n_264) );
AND2x4_ASAP7_75t_L g320 ( .A(n_146), .B(n_232), .Y(n_320) );
OR2x2_ASAP7_75t_L g335 ( .A(n_146), .B(n_255), .Y(n_335) );
OR2x2_ASAP7_75t_L g361 ( .A(n_146), .B(n_217), .Y(n_361) );
AND2x2_ASAP7_75t_L g369 ( .A(n_146), .B(n_315), .Y(n_369) );
AND2x4_ASAP7_75t_SL g394 ( .A(n_146), .B(n_314), .Y(n_394) );
OR2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_154), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_154), .B(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_154), .B(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_154), .B(n_196), .Y(n_195) );
NOR3xp33_ASAP7_75t_L g199 ( .A(n_154), .B(n_200), .C(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_154), .A2(n_445), .B(n_450), .Y(n_444) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_156), .B(n_314), .Y(n_390) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_166), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_157), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OR2x6_ASAP7_75t_SL g214 ( .A(n_158), .B(n_215), .Y(n_214) );
INVxp67_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g239 ( .A(n_159), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_159), .B(n_274), .Y(n_292) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_159), .Y(n_430) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g247 ( .A(n_160), .Y(n_247) );
AND2x2_ASAP7_75t_L g272 ( .A(n_160), .B(n_203), .Y(n_272) );
INVx2_ASAP7_75t_L g300 ( .A(n_160), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_160), .B(n_167), .Y(n_341) );
BUFx3_ASAP7_75t_L g365 ( .A(n_160), .Y(n_365) );
OR2x2_ASAP7_75t_L g377 ( .A(n_160), .B(n_167), .Y(n_377) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_160), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_166), .A2(n_408), .B1(n_411), .B2(n_412), .Y(n_407) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_177), .Y(n_166) );
INVx1_ASAP7_75t_L g235 ( .A(n_167), .Y(n_235) );
OR2x2_ASAP7_75t_L g246 ( .A(n_167), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g253 ( .A(n_167), .Y(n_253) );
AND2x4_ASAP7_75t_SL g270 ( .A(n_167), .B(n_178), .Y(n_270) );
AND2x4_ASAP7_75t_L g275 ( .A(n_167), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g284 ( .A(n_167), .Y(n_284) );
OR2x2_ASAP7_75t_L g290 ( .A(n_167), .B(n_178), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_167), .B(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_167), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_167), .B(n_272), .Y(n_406) );
OR2x2_ASAP7_75t_L g422 ( .A(n_167), .B(n_325), .Y(n_422) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_176), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_174), .Y(n_168) );
INVx2_ASAP7_75t_SL g257 ( .A(n_174), .Y(n_257) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_174), .A2(n_505), .B(n_509), .Y(n_504) );
BUFx4f_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g198 ( .A(n_175), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_177), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g248 ( .A(n_177), .Y(n_248) );
AND2x2_ASAP7_75t_SL g355 ( .A(n_177), .B(n_239), .Y(n_355) );
AND2x4_ASAP7_75t_L g177 ( .A(n_178), .B(n_202), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_178), .B(n_203), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_178), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_178), .B(n_247), .Y(n_251) );
INVx3_ASAP7_75t_L g276 ( .A(n_178), .Y(n_276) );
INVx1_ASAP7_75t_L g309 ( .A(n_178), .Y(n_309) );
AND2x2_ASAP7_75t_L g389 ( .A(n_178), .B(n_253), .Y(n_389) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_194), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_182), .B1(n_187), .B2(n_192), .Y(n_179) );
INVx1_ASAP7_75t_L g477 ( .A(n_182), .Y(n_477) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_186), .Y(n_182) );
INVx1_ASAP7_75t_L g518 ( .A(n_183), .Y(n_518) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
OR2x6_ASAP7_75t_L g448 ( .A(n_184), .B(n_191), .Y(n_448) );
INVxp33_ASAP7_75t_L g494 ( .A(n_184), .Y(n_494) );
INVx1_ASAP7_75t_L g519 ( .A(n_186), .Y(n_519) );
INVxp67_ASAP7_75t_L g475 ( .A(n_187), .Y(n_475) );
NOR2x1p5_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVx1_ASAP7_75t_L g495 ( .A(n_190), .Y(n_495) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_197), .A2(n_464), .B1(n_469), .B2(n_470), .Y(n_463) );
INVx3_ASAP7_75t_L g470 ( .A(n_197), .Y(n_470) );
INVx4_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI21x1_ASAP7_75t_L g204 ( .A1(n_198), .A2(n_205), .B(n_211), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_198), .B(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_201), .B(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_201), .A2(n_448), .B1(n_530), .B2(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_203), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g274 ( .A(n_203), .Y(n_274) );
AND2x2_ASAP7_75t_L g299 ( .A(n_203), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g325 ( .A(n_203), .B(n_247), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_203), .B(n_276), .Y(n_342) );
INVx1_ASAP7_75t_L g348 ( .A(n_203), .Y(n_348) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_210), .Y(n_205) );
AOI222xp33_ASAP7_75t_SL g212 ( .A1(n_213), .A2(n_216), .B1(n_226), .B2(n_233), .C1(n_236), .C2(n_240), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_225), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_217), .B(n_286), .Y(n_337) );
AND2x4_ASAP7_75t_L g353 ( .A(n_217), .B(n_264), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_223), .Y(n_218) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_228), .B(n_230), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g278 ( .A(n_229), .B(n_279), .Y(n_278) );
AOI222xp33_ASAP7_75t_L g243 ( .A1(n_230), .A2(n_244), .B1(n_249), .B2(n_254), .C1(n_262), .C2(n_810), .Y(n_243) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g382 ( .A(n_231), .B(n_286), .Y(n_382) );
OR2x2_ASAP7_75t_L g425 ( .A(n_231), .B(n_331), .Y(n_425) );
AND2x2_ASAP7_75t_L g254 ( .A(n_232), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g315 ( .A(n_232), .Y(n_315) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_232), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_233), .A2(n_344), .B(n_349), .C(n_350), .Y(n_343) );
INVx1_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g371 ( .A(n_235), .Y(n_371) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g301 ( .A(n_240), .Y(n_301) );
AND2x2_ASAP7_75t_L g285 ( .A(n_241), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g294 ( .A(n_241), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OAI31xp33_ASAP7_75t_L g336 ( .A1(n_244), .A2(n_262), .A3(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_245), .A2(n_295), .B(n_339), .C(n_340), .Y(n_338) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
OR2x2_ASAP7_75t_L g327 ( .A(n_246), .B(n_276), .Y(n_327) );
INVx2_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
BUFx2_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
AND2x2_ASAP7_75t_L g304 ( .A(n_255), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_256), .Y(n_286) );
AOI21x1_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_261), .Y(n_256) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_257), .A2(n_489), .B(n_497), .Y(n_488) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_257), .A2(n_489), .B(n_497), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_264), .B(n_321), .Y(n_413) );
OAI211xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_277), .B(n_280), .C(n_302), .Y(n_265) );
INVxp33_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_268), .B(n_273), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g306 ( .A(n_270), .B(n_299), .Y(n_306) );
OR2x2_ASAP7_75t_L g282 ( .A(n_271), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g312 ( .A(n_271), .B(n_286), .Y(n_312) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g388 ( .A(n_272), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g411 ( .A(n_273), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_275), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_275), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g423 ( .A(n_275), .B(n_299), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_275), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g366 ( .A(n_276), .B(n_348), .Y(n_366) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AOI322xp5_ASAP7_75t_L g420 ( .A1(n_279), .A2(n_299), .A3(n_353), .B1(n_378), .B2(n_421), .C1(n_423), .C2(n_424), .Y(n_420) );
AOI211xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_285), .B(n_287), .C(n_296), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_283), .B(n_311), .Y(n_333) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g298 ( .A(n_284), .B(n_299), .Y(n_298) );
NOR2x1p5_ASAP7_75t_L g364 ( .A(n_284), .B(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_284), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_285), .A2(n_303), .B(n_306), .C(n_307), .Y(n_302) );
AND2x4_ASAP7_75t_L g321 ( .A(n_286), .B(n_305), .Y(n_321) );
INVx2_ASAP7_75t_L g331 ( .A(n_286), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_286), .B(n_320), .Y(n_351) );
AND2x2_ASAP7_75t_L g393 ( .A(n_286), .B(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_286), .B(n_410), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_286), .B(n_314), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_291), .B(n_293), .Y(n_287) );
AND2x2_ASAP7_75t_L g383 ( .A(n_289), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g311 ( .A(n_292), .Y(n_311) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_304), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g398 ( .A(n_304), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_310), .B(n_312), .C(n_313), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_311), .Y(n_395) );
INVx3_ASAP7_75t_SL g410 ( .A(n_314), .Y(n_410) );
NAND5xp2_ASAP7_75t_L g316 ( .A(n_317), .B(n_336), .C(n_343), .D(n_356), .E(n_367), .Y(n_316) );
AOI222xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_322), .B1(n_326), .B2(n_328), .C1(n_332), .C2(n_334), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_319), .A2(n_400), .B1(n_404), .B2(n_405), .Y(n_399) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g349 ( .A(n_320), .B(n_321), .Y(n_349) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_330), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_331), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g368 ( .A(n_331), .B(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g379 ( .A(n_331), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g409 ( .A(n_335), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g357 ( .A(n_342), .Y(n_357) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B(n_354), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_353), .A2(n_357), .B1(n_358), .B2(n_362), .Y(n_356) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
INVx2_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g370 ( .A(n_355), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g375 ( .A(n_357), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
INVx1_ASAP7_75t_SL g403 ( .A(n_366), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
NOR3xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_391), .C(n_414), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_374), .B(n_390), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_381), .B2(n_383), .C(n_386), .Y(n_374) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g415 ( .A(n_377), .B(n_403), .Y(n_415) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
OAI321xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .A3(n_396), .B1(n_398), .B2(n_399), .C(n_407), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_405), .A2(n_427), .B1(n_431), .B2(n_432), .Y(n_426) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI211xp5_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_416), .B(n_420), .C(n_426), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_434), .B(n_754), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_704), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_644), .B(n_703), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g754 ( .A(n_436), .B(n_705), .C(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g794 ( .A(n_436), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_608), .Y(n_436) );
NOR3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_549), .C(n_578), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_439), .B(n_538), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_459), .B1(n_498), .B2(n_510), .Y(n_439) );
NAND2x1_ASAP7_75t_L g740 ( .A(n_440), .B(n_539), .Y(n_740) );
INVx2_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_451), .Y(n_441) );
INVx2_ASAP7_75t_L g512 ( .A(n_442), .Y(n_512) );
INVx4_ASAP7_75t_L g554 ( .A(n_442), .Y(n_554) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_442), .Y(n_574) );
AND2x4_ASAP7_75t_L g585 ( .A(n_442), .B(n_553), .Y(n_585) );
AND2x2_ASAP7_75t_L g591 ( .A(n_442), .B(n_515), .Y(n_591) );
NOR2x1_ASAP7_75t_SL g664 ( .A(n_442), .B(n_526), .Y(n_664) );
OR2x6_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVxp67_ASAP7_75t_L g465 ( .A(n_448), .Y(n_465) );
INVx2_ASAP7_75t_L g525 ( .A(n_448), .Y(n_525) );
INVx2_ASAP7_75t_L g557 ( .A(n_451), .Y(n_557) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_451), .Y(n_571) );
INVx1_ASAP7_75t_L g582 ( .A(n_451), .Y(n_582) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_451), .Y(n_594) );
AND2x2_ASAP7_75t_L g626 ( .A(n_451), .B(n_526), .Y(n_626) );
INVx1_ASAP7_75t_L g652 ( .A(n_451), .Y(n_652) );
AND2x2_ASAP7_75t_L g714 ( .A(n_451), .B(n_542), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_478), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g607 ( .A(n_461), .B(n_546), .Y(n_607) );
INVx2_ASAP7_75t_L g649 ( .A(n_461), .Y(n_649) );
AND2x2_ASAP7_75t_L g751 ( .A(n_461), .B(n_478), .Y(n_751) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_462), .B(n_501), .Y(n_545) );
INVx2_ASAP7_75t_L g566 ( .A(n_462), .Y(n_566) );
AND2x4_ASAP7_75t_L g588 ( .A(n_462), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g623 ( .A(n_462), .Y(n_623) );
AND2x2_ASAP7_75t_L g747 ( .A(n_462), .B(n_504), .Y(n_747) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_471), .Y(n_462) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_470), .A2(n_480), .B(n_486), .Y(n_479) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_470), .A2(n_480), .B(n_486), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_475), .B1(n_476), .B2(n_477), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g721 ( .A(n_478), .Y(n_721) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_487), .Y(n_478) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_479), .B(n_566), .Y(n_596) );
AND2x2_ASAP7_75t_L g601 ( .A(n_479), .B(n_566), .Y(n_601) );
INVx2_ASAP7_75t_L g614 ( .A(n_479), .Y(n_614) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_479), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
AND2x4_ASAP7_75t_L g587 ( .A(n_487), .B(n_500), .Y(n_587) );
AND2x2_ASAP7_75t_L g602 ( .A(n_487), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g657 ( .A(n_487), .Y(n_657) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_488), .B(n_504), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_488), .B(n_501), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_490), .B(n_496), .Y(n_489) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVxp33_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
INVx3_ASAP7_75t_L g563 ( .A(n_500), .Y(n_563) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_501), .Y(n_561) );
AND2x2_ASAP7_75t_L g675 ( .A(n_501), .B(n_676), .Y(n_675) );
INVx3_ASAP7_75t_L g618 ( .A(n_502), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_502), .B(n_657), .Y(n_698) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g565 ( .A(n_503), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g546 ( .A(n_504), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g589 ( .A(n_504), .Y(n_589) );
INVxp67_ASAP7_75t_L g603 ( .A(n_504), .Y(n_603) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_504), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_504), .Y(n_680) );
INVx1_ASAP7_75t_L g658 ( .A(n_510), .Y(n_658) );
NOR2x1_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_511), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g700 ( .A(n_512), .B(n_541), .Y(n_700) );
OR2x2_ASAP7_75t_L g752 ( .A(n_513), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g651 ( .A(n_514), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g687 ( .A(n_514), .B(n_574), .Y(n_687) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_526), .Y(n_514) );
AND2x4_ASAP7_75t_L g541 ( .A(n_515), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g553 ( .A(n_515), .Y(n_553) );
INVx2_ASAP7_75t_L g570 ( .A(n_515), .Y(n_570) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_515), .Y(n_696) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_521), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .C(n_520), .Y(n_517) );
INVx3_ASAP7_75t_L g542 ( .A(n_526), .Y(n_542) );
INVx2_ASAP7_75t_L g636 ( .A(n_526), .Y(n_636) );
AND2x4_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_532), .B(n_537), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B1(n_535), .B2(n_536), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_540), .B(n_616), .Y(n_633) );
NOR2x1_ASAP7_75t_L g725 ( .A(n_540), .B(n_554), .Y(n_725) );
INVx4_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_541), .B(n_616), .Y(n_702) );
AND2x2_ASAP7_75t_L g569 ( .A(n_542), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g583 ( .A(n_542), .Y(n_583) );
AOI22xp5_ASAP7_75t_SL g631 ( .A1(n_543), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_631) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g628 ( .A(n_544), .B(n_602), .Y(n_628) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g736 ( .A(n_545), .B(n_577), .Y(n_736) );
AND2x2_ASAP7_75t_L g559 ( .A(n_546), .B(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g595 ( .A(n_546), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g738 ( .A(n_546), .B(n_649), .Y(n_738) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g613 ( .A(n_548), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g639 ( .A(n_548), .Y(n_639) );
AND2x2_ASAP7_75t_L g674 ( .A(n_548), .B(n_566), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_558), .B1(n_562), .B2(n_567), .C(n_572), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_L g630 ( .A(n_552), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_552), .B(n_626), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_552), .B(n_714), .Y(n_713) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NOR2xp67_ASAP7_75t_SL g598 ( .A(n_554), .B(n_599), .Y(n_598) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_554), .Y(n_611) );
AND2x4_ASAP7_75t_SL g695 ( .A(n_554), .B(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g742 ( .A(n_554), .B(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx3_ASAP7_75t_L g616 ( .A(n_556), .Y(n_616) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_557), .Y(n_753) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI221x1_ASAP7_75t_L g706 ( .A1(n_559), .A2(n_707), .B1(n_709), .B2(n_710), .C(n_712), .Y(n_706) );
AND2x2_ASAP7_75t_L g632 ( .A(n_560), .B(n_588), .Y(n_632) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AND2x2_ASAP7_75t_L g575 ( .A(n_563), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_563), .B(n_565), .Y(n_749) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND2x2_ASAP7_75t_SL g573 ( .A(n_569), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_569), .B(n_582), .Y(n_599) );
INVx2_ASAP7_75t_L g606 ( .A(n_569), .Y(n_606) );
INVx1_ASAP7_75t_L g668 ( .A(n_570), .Y(n_668) );
BUFx2_ASAP7_75t_L g688 ( .A(n_571), .Y(n_688) );
NAND2xp33_ASAP7_75t_SL g572 ( .A(n_573), .B(n_575), .Y(n_572) );
OR2x6_ASAP7_75t_L g605 ( .A(n_574), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g734 ( .A(n_574), .B(n_626), .Y(n_734) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_597), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_586), .B1(n_590), .B2(n_595), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_581), .B(n_585), .Y(n_643) );
AND2x4_ASAP7_75t_L g709 ( .A(n_581), .B(n_667), .Y(n_709) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_582), .B(n_583), .Y(n_581) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_582), .Y(n_724) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_585), .B(n_625), .Y(n_624) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_585), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_585), .B(n_616), .Y(n_708) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
AND2x2_ASAP7_75t_L g729 ( .A(n_587), .B(n_648), .Y(n_729) );
INVx3_ASAP7_75t_L g640 ( .A(n_588), .Y(n_640) );
AND2x2_ASAP7_75t_L g661 ( .A(n_588), .B(n_613), .Y(n_661) );
NAND2x1_ASAP7_75t_SL g732 ( .A(n_588), .B(n_639), .Y(n_732) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B1(n_604), .B2(n_607), .Y(n_597) );
BUFx2_ASAP7_75t_L g653 ( .A(n_599), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_600), .A2(n_691), .B1(n_700), .B2(n_701), .Y(n_699) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_601), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g621 ( .A(n_602), .B(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_606), .B(n_686), .C(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g641 ( .A(n_607), .Y(n_641) );
AOI211x1_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_617), .B(n_619), .C(n_637), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_612), .B(n_700), .Y(n_719) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_613), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g691 ( .A(n_613), .B(n_649), .Y(n_691) );
AND2x2_ASAP7_75t_L g746 ( .A(n_613), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g669 ( .A(n_616), .Y(n_669) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g711 ( .A(n_618), .B(n_656), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_631), .Y(n_619) );
AOI22xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_624), .B1(n_627), .B2(n_629), .Y(n_620) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g684 ( .A(n_623), .B(n_679), .Y(n_684) );
INVx1_ASAP7_75t_SL g726 ( .A(n_623), .Y(n_726) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_SL g694 ( .A(n_626), .B(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVxp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g730 ( .A(n_635), .B(n_652), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_641), .B(n_642), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_639), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g654 ( .A(n_640), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_644), .Y(n_796) );
NAND3x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_681), .C(n_689), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g755 ( .A(n_645), .B(n_681), .C(n_689), .D(n_756), .Y(n_755) );
NOR2x1_ASAP7_75t_L g645 ( .A(n_646), .B(n_659), .Y(n_645) );
OAI222xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_650), .B1(n_653), .B2(n_654), .C1(n_656), .C2(n_658), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI21xp5_ASAP7_75t_SL g733 ( .A1(n_651), .A2(n_734), .B(n_735), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_652), .B(n_667), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_655), .A2(n_713), .B1(n_715), .B2(n_716), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_670), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_663), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_667), .B(n_669), .Y(n_672) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .B1(n_677), .B2(n_678), .Y(n_670) );
AND2x4_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
AND2x2_ASAP7_75t_L g678 ( .A(n_674), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_682), .B(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g715 ( .A(n_684), .Y(n_715) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_699), .Y(n_689) );
AOI22xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_692), .B1(n_694), .B2(n_697), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp33_ASAP7_75t_L g704 ( .A(n_703), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g795 ( .A(n_705), .Y(n_795) );
NAND3x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_717), .C(n_737), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_709), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g743 ( .A(n_714), .Y(n_743) );
NOR2x1_ASAP7_75t_L g717 ( .A(n_718), .B(n_727), .Y(n_717) );
AOI21xp5_ASAP7_75t_SL g718 ( .A1(n_719), .A2(n_720), .B(n_726), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_733), .Y(n_727) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_732), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B1(n_741), .B2(n_744), .C(n_748), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVxp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B(n_752), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g762 ( .A(n_759), .Y(n_762) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx2_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
INVx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_781), .Y(n_774) );
INVxp67_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_777), .B(n_780), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OR2x2_ASAP7_75t_SL g799 ( .A(n_778), .B(n_780), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_778), .A2(n_804), .B(n_807), .Y(n_803) );
INVx1_ASAP7_75t_SL g786 ( .A(n_781), .Y(n_786) );
BUFx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
BUFx2_ASAP7_75t_L g808 ( .A(n_782), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_787), .B(n_797), .Y(n_783) );
CKINVDCx11_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B1(n_792), .B2(n_793), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AND3x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .C(n_796), .Y(n_793) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
CKINVDCx11_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
CKINVDCx8_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
endmodule