module fake_jpeg_32132_n_445 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_445);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_445;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_9),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_64),
.Y(n_103)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx2_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

NAND2x1_ASAP7_75t_SL g124 ( 
.A(n_70),
.B(n_81),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_72),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_76),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_24),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_80),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_82),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_30),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_84),
.Y(n_113)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_87),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_88),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_43),
.C(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_94),
.B(n_57),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_23),
.B1(n_27),
.B2(n_33),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_97),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_114),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_45),
.B(n_42),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_48),
.B(n_42),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_51),
.B(n_33),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_31),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_40),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_46),
.B(n_40),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_65),
.B(n_38),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_114),
.Y(n_158)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_56),
.Y(n_198)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_154),
.B1(n_168),
.B2(n_170),
.Y(n_176)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_25),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_155),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_97),
.A2(n_62),
.B1(n_68),
.B2(n_47),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_150),
.A2(n_96),
.B1(n_102),
.B2(n_101),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_109),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_157),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_81),
.B1(n_75),
.B2(n_85),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_104),
.B(n_26),
.Y(n_155)
);

CKINVDCx12_ASAP7_75t_R g157 ( 
.A(n_99),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_159),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_92),
.B(n_35),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_160),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_166),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_164),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_103),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_169),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_118),
.A2(n_88),
.B1(n_84),
.B2(n_52),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_67),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_124),
.A2(n_50),
.B1(n_44),
.B2(n_60),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_148),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_124),
.A2(n_61),
.B1(n_49),
.B2(n_31),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_53),
.B1(n_135),
.B2(n_121),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_141),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_109),
.B1(n_157),
.B2(n_135),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_94),
.B1(n_93),
.B2(n_131),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_192),
.A2(n_195),
.B1(n_202),
.B2(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_89),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_201),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_95),
.B1(n_108),
.B2(n_93),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_89),
.B(n_98),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_196),
.B(n_187),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_154),
.C(n_149),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_122),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_204),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_208),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_163),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_146),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_212),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_216),
.B1(n_181),
.B2(n_186),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_213),
.B(n_220),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_167),
.Y(n_214)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_215),
.A2(n_223),
.B1(n_227),
.B2(n_194),
.Y(n_249)
);

AO21x2_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_140),
.B(n_165),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_155),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_218),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_162),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_145),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_221),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_222),
.A2(n_199),
.B(n_174),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_196),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_164),
.C(n_152),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_102),
.C(n_101),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_188),
.B1(n_134),
.B2(n_110),
.Y(n_229)
);

NOR2x1_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_153),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_222),
.B(n_223),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_176),
.A3(n_188),
.B1(n_183),
.B2(n_122),
.Y(n_228)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_219),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_231),
.B(n_205),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_131),
.B1(n_95),
.B2(n_191),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_237),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_250),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_191),
.B1(n_143),
.B2(n_165),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_216),
.B(n_224),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_207),
.A2(n_143),
.B1(n_137),
.B2(n_140),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_181),
.B(n_184),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_216),
.B(n_204),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_99),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_205),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_137),
.B1(n_175),
.B2(n_178),
.Y(n_245)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_139),
.B1(n_178),
.B2(n_173),
.Y(n_246)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_139),
.B1(n_173),
.B2(n_175),
.Y(n_248)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_252),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_209),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_254),
.B(n_259),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_216),
.B1(n_227),
.B2(n_203),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_257),
.A2(n_251),
.B1(n_233),
.B2(n_173),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_247),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_258),
.Y(n_280)
);

NOR3xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_226),
.C(n_212),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_247),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_260),
.B(n_273),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_262),
.A2(n_268),
.B(n_189),
.Y(n_307)
);

AND2x6_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_208),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_264),
.Y(n_281)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_208),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_277),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_208),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_275),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_230),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_230),
.C(n_231),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_242),
.B(n_217),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_244),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_274),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_276),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_232),
.B(n_208),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_251),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_90),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_245),
.B1(n_240),
.B2(n_234),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_285),
.A2(n_296),
.B1(n_299),
.B2(n_227),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_289),
.C(n_293),
.Y(n_312)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_243),
.C(n_232),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_253),
.A2(n_246),
.B1(n_248),
.B2(n_237),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_292),
.A2(n_283),
.B1(n_294),
.B2(n_307),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_250),
.C(n_229),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_0),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_251),
.B1(n_238),
.B2(n_233),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_206),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_300),
.B(n_302),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_206),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_253),
.B(n_221),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_304),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_264),
.B(n_213),
.CI(n_99),
.CON(n_304),
.SN(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_279),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_306),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_252),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_261),
.B(n_270),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_262),
.C(n_252),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_265),
.C(n_261),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_215),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_263),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_329),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_315),
.A2(n_308),
.B(n_303),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_290),
.A2(n_270),
.B1(n_271),
.B2(n_255),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_316),
.A2(n_166),
.B1(n_136),
.B2(n_160),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_271),
.Y(n_318)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_256),
.Y(n_319)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_321),
.B(n_332),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_256),
.C(n_182),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_331),
.C(n_333),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_324),
.A2(n_285),
.B1(n_288),
.B2(n_282),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_287),
.B(n_194),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_330),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_292),
.B1(n_291),
.B2(n_299),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_301),
.A2(n_138),
.B(n_142),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_327),
.A2(n_328),
.B(n_147),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_301),
.A2(n_281),
.B(n_309),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_215),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_199),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_289),
.B(n_182),
.C(n_90),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_293),
.B(n_147),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_0),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_335),
.A2(n_344),
.B1(n_349),
.B2(n_353),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_311),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_332),
.Y(n_364)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_129),
.B(n_91),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_304),
.C(n_296),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_342),
.C(n_352),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_304),
.C(n_297),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_343),
.A2(n_347),
.B1(n_327),
.B2(n_329),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_320),
.A2(n_298),
.B1(n_282),
.B2(n_160),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_315),
.A2(n_100),
.B(n_96),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_345),
.A2(n_338),
.B(n_354),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_321),
.A2(n_328),
.B1(n_317),
.B2(n_323),
.Y(n_349)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_351),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_129),
.C(n_128),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_324),
.A2(n_106),
.B1(n_123),
.B2(n_121),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_311),
.A2(n_31),
.B1(n_43),
.B2(n_123),
.Y(n_355)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_147),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_0),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_333),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_314),
.B(n_16),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_358),
.B(n_10),
.Y(n_361)
);

NOR3xp33_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_318),
.C(n_313),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_359),
.Y(n_383)
);

BUFx12_ASAP7_75t_L g360 ( 
.A(n_357),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_373),
.Y(n_380)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_330),
.C(n_319),
.Y(n_362)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_363),
.B(n_375),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_364),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_368),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_370),
.Y(n_385)
);

NOR2x1_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_331),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_371),
.B(n_374),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_352),
.B(n_18),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_17),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_109),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_335),
.A2(n_31),
.B1(n_43),
.B2(n_128),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_378),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_350),
.B(n_340),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_SL g384 ( 
.A(n_379),
.B(n_350),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_375),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_379),
.A2(n_341),
.B(n_345),
.Y(n_386)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_367),
.B(n_336),
.C(n_346),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_389),
.C(n_366),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_336),
.C(n_343),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_344),
.B1(n_353),
.B2(n_43),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_394),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_14),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_383),
.B(n_372),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_401),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_392),
.A2(n_370),
.B(n_378),
.Y(n_397)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_397),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_405),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_403),
.C(n_393),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_381),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_389),
.B(n_365),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_402),
.B(n_404),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_369),
.C(n_363),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_360),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_371),
.C(n_374),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_368),
.C(n_91),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_380),
.C(n_382),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_388),
.B(n_12),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_408),
.B(n_17),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_403),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_410),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_415),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_401),
.A2(n_385),
.B1(n_381),
.B2(n_391),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_416),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_391),
.C(n_386),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_418),
.B(n_130),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_400),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_419),
.A2(n_420),
.B1(n_69),
.B2(n_79),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_407),
.A2(n_66),
.B(n_82),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_424),
.Y(n_431)
);

AOI322xp5_ASAP7_75t_L g425 ( 
.A1(n_417),
.A2(n_130),
.A3(n_15),
.B1(n_14),
.B2(n_11),
.C1(n_8),
.C2(n_63),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_425),
.B(n_429),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_409),
.A2(n_14),
.B(n_11),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_426),
.A2(n_414),
.B(n_413),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_11),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_428),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_1),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_430),
.B(n_434),
.C(n_7),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_423),
.B(n_411),
.Y(n_433)
);

AO21x1_ASAP7_75t_L g439 ( 
.A1(n_433),
.A2(n_432),
.B(n_5),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_422),
.A2(n_1),
.B(n_3),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g436 ( 
.A1(n_431),
.A2(n_425),
.B(n_3),
.C(n_4),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_436),
.A2(n_4),
.B(n_5),
.Y(n_440)
);

NOR3xp33_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_438),
.C(n_439),
.Y(n_441)
);

O2A1O1Ixp33_ASAP7_75t_SL g438 ( 
.A1(n_435),
.A2(n_1),
.B(n_4),
.C(n_5),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_440),
.B(n_5),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_442),
.A2(n_441),
.B1(n_6),
.B2(n_7),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_443),
.B(n_6),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_6),
.Y(n_445)
);


endmodule