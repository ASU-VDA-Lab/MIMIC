module fake_jpeg_27957_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_2),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_26),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_16),
.B1(n_25),
.B2(n_20),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_61),
.B1(n_72),
.B2(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_31),
.B1(n_25),
.B2(n_16),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_63),
.B1(n_44),
.B2(n_34),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_51),
.B(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_26),
.C(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_60),
.B(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_19),
.B1(n_29),
.B2(n_32),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_71),
.Y(n_77)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_22),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_22),
.B1(n_15),
.B2(n_6),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_36),
.B(n_15),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_9),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_78),
.Y(n_109)
);

INVx5_ASAP7_75t_SL g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_81),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_73),
.B1(n_52),
.B2(n_48),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_34),
.B1(n_44),
.B2(n_6),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_86),
.Y(n_118)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_35),
.B1(n_40),
.B2(n_7),
.Y(n_88)
);

OAI21x1_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_68),
.B(n_52),
.Y(n_121)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_10),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_93),
.Y(n_105)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_9),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_40),
.B1(n_4),
.B2(n_7),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_51),
.B1(n_59),
.B2(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_48),
.Y(n_115)
);

NAND2x1_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_57),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_115),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_56),
.C(n_59),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_122),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_116),
.B1(n_89),
.B2(n_88),
.Y(n_146)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_77),
.B(n_50),
.CI(n_51),
.CON(n_113),
.SN(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_126),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_101),
.B1(n_103),
.B2(n_102),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_69),
.C(n_68),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_3),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_129),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_94),
.C(n_14),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_92),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_138),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_144),
.B1(n_146),
.B2(n_110),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_105),
.B(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_145),
.Y(n_150)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_139),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_92),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_140),
.A2(n_91),
.B1(n_117),
.B2(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_143),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_114),
.A2(n_88),
.B1(n_79),
.B2(n_86),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_123),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_141),
.A2(n_125),
.B1(n_114),
.B2(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_149),
.A2(n_154),
.B1(n_142),
.B2(n_127),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_88),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_156),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_106),
.CI(n_113),
.CON(n_156),
.SN(n_156)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_144),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_130),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_130),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_161),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_170),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_163),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_130),
.C(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_171),
.C(n_172),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_169),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_131),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_104),
.C(n_109),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_182),
.Y(n_187)
);

AOI21x1_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_170),
.B(n_172),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_179),
.Y(n_185)
);

AOI321xp33_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_150),
.A3(n_156),
.B1(n_147),
.B2(n_160),
.C(n_149),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_151),
.C(n_161),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_174),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_184),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_170),
.B1(n_162),
.B2(n_147),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_155),
.B(n_156),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_188),
.Y(n_189)
);

NOR2xp67_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_148),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_191),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_187),
.B(n_178),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_175),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_13),
.B(n_83),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_183),
.B1(n_104),
.B2(n_109),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_194),
.A2(n_196),
.B(n_100),
.C(n_83),
.Y(n_198)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_13),
.B(n_78),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_96),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_195),
.B(n_194),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_199),
.Y(n_202)
);


endmodule