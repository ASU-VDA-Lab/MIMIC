module fake_jpeg_17228_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_260;
wire n_112;
wire n_199;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_23),
.C(n_19),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_40),
.C(n_19),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_38),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_38),
.B1(n_39),
.B2(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_20),
.B1(n_17),
.B2(n_24),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_76),
.B1(n_28),
.B2(n_24),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_68),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_37),
.B1(n_38),
.B2(n_33),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_80),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_20),
.B1(n_17),
.B2(n_22),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

CKINVDCx12_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_48),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_35),
.B1(n_37),
.B2(n_36),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_35),
.B1(n_20),
.B2(n_58),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_47),
.B(n_48),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_22),
.B(n_29),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_94),
.Y(n_114)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_20),
.B1(n_33),
.B2(n_47),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_104),
.B1(n_61),
.B2(n_59),
.Y(n_116)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_33),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_39),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_106),
.Y(n_122)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_68),
.B1(n_71),
.B2(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_105),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_110),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_23),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_82),
.C(n_74),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_73),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_74),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_120),
.B(n_95),
.Y(n_151)
);

OAI22x1_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_124),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_126),
.B1(n_129),
.B2(n_136),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_114),
.C(n_124),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_28),
.B(n_24),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_84),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_66),
.B1(n_71),
.B2(n_65),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_65),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_86),
.A2(n_78),
.B1(n_34),
.B2(n_56),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_57),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_72),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_23),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_105),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_60),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_93),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_34),
.B1(n_22),
.B2(n_31),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_86),
.B1(n_98),
.B2(n_107),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_138),
.A2(n_121),
.B1(n_135),
.B2(n_111),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_98),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_155),
.C(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_143),
.A2(n_149),
.B(n_25),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_161),
.B1(n_89),
.B2(n_135),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_30),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_153),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_90),
.B1(n_96),
.B2(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_99),
.B1(n_101),
.B2(n_90),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_156),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_165),
.B(n_29),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_96),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_159),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_103),
.A3(n_29),
.B1(n_30),
.B2(n_16),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_162),
.B(n_125),
.Y(n_174)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_106),
.C(n_34),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_110),
.B1(n_108),
.B2(n_89),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_113),
.B(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_112),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_134),
.C(n_120),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_166),
.C(n_34),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_26),
.B1(n_31),
.B2(n_30),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_34),
.C(n_56),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_27),
.C(n_25),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_27),
.Y(n_190)
);

AND2x4_ASAP7_75t_SL g168 ( 
.A(n_148),
.B(n_137),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_168),
.A2(n_49),
.B(n_1),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_118),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_192),
.C(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_115),
.B1(n_112),
.B2(n_128),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_177),
.B1(n_182),
.B2(n_184),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_176),
.B(n_193),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_144),
.B1(n_150),
.B2(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_128),
.B(n_111),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_185),
.B(n_190),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_111),
.Y(n_187)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_25),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_189),
.B(n_191),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_25),
.Y(n_191)
);

CKINVDCx12_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_49),
.B1(n_43),
.B2(n_31),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_194),
.A2(n_196),
.B1(n_165),
.B2(n_16),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_R g195 ( 
.A(n_157),
.B(n_27),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_195),
.B(n_21),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_143),
.A2(n_16),
.B1(n_26),
.B2(n_21),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_204),
.C(n_194),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_207),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_205),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_138),
.A3(n_153),
.B1(n_154),
.B2(n_26),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_203),
.B(n_190),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_49),
.C(n_21),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_172),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_215),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_0),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_209),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_217),
.B1(n_218),
.B2(n_8),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_181),
.B1(n_168),
.B2(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_181),
.B1(n_192),
.B2(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_174),
.C(n_183),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_222),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_182),
.B1(n_180),
.B2(n_185),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_227),
.C(n_236),
.Y(n_242)
);

OA21x2_ASAP7_75t_SL g225 ( 
.A1(n_219),
.A2(n_175),
.B(n_176),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_201),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_175),
.C(n_196),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_216),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_235),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_238),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_2),
.C(n_3),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_9),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_226),
.C(n_236),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_251),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_211),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_246),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_214),
.C(n_216),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_234),
.C(n_209),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_223),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_251),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_259),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_205),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_221),
.C(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_242),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_231),
.B1(n_200),
.B2(n_222),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_261),
.A2(n_252),
.B1(n_248),
.B2(n_246),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_266),
.Y(n_271)
);

AO221x1_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_213),
.B1(n_229),
.B2(n_220),
.C(n_199),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_264),
.Y(n_276)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_267),
.B(n_274),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_240),
.C(n_237),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_271),
.B(n_268),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_277),
.C(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_257),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_262),
.A2(n_199),
.B(n_235),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_256),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_203),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_283),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_284),
.B(n_11),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_282),
.C(n_285),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_265),
.C(n_198),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_258),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_208),
.B(n_228),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_208),
.B1(n_210),
.B2(n_7),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_11),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_281),
.A2(n_267),
.B1(n_275),
.B2(n_7),
.Y(n_287)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_289),
.A2(n_292),
.B1(n_8),
.B2(n_9),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_8),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_11),
.C(n_6),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_293),
.A2(n_295),
.B(n_292),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_296),
.B(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_288),
.C(n_291),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_293),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_12),
.B(n_13),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_14),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_4),
.Y(n_302)
);


endmodule