module fake_jpeg_587_n_542 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_542);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_50),
.Y(n_140)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_52),
.Y(n_125)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_56),
.B(n_59),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_0),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_60),
.Y(n_131)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_62),
.Y(n_154)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_69),
.B(n_78),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_13),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_16),
.B(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_97),
.Y(n_106)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_95),
.Y(n_151)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_96),
.Y(n_134)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_13),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_102),
.Y(n_152)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_17),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_104),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_42),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_56),
.A2(n_59),
.B1(n_22),
.B2(n_32),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_113),
.A2(n_160),
.B1(n_161),
.B2(n_27),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_32),
.B1(n_22),
.B2(n_46),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_121),
.A2(n_157),
.B1(n_48),
.B2(n_30),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_55),
.A2(n_36),
.B1(n_47),
.B2(n_46),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_123),
.A2(n_147),
.B1(n_150),
.B2(n_164),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_54),
.A2(n_19),
.B1(n_14),
.B2(n_26),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_138),
.A2(n_139),
.B1(n_28),
.B2(n_65),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_54),
.A2(n_19),
.B1(n_14),
.B2(n_26),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_64),
.A2(n_36),
.B1(n_47),
.B2(n_19),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_67),
.A2(n_14),
.B1(n_45),
.B2(n_43),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_76),
.A2(n_79),
.B1(n_88),
.B2(n_86),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_94),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_74),
.A2(n_17),
.B1(n_45),
.B2(n_43),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_58),
.A2(n_20),
.B1(n_45),
.B2(n_43),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_162),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_90),
.A2(n_20),
.B1(n_42),
.B2(n_39),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_82),
.A2(n_20),
.B1(n_42),
.B2(n_39),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_39),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_170),
.B(n_172),
.Y(n_243)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_171),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_57),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_113),
.A2(n_105),
.B1(n_73),
.B2(n_85),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_176),
.A2(n_177),
.B1(n_187),
.B2(n_213),
.Y(n_221)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_57),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_194),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_81),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_129),
.Y(n_184)
);

BUFx24_ASAP7_75t_L g255 ( 
.A(n_184),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_101),
.B1(n_98),
.B2(n_62),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_185),
.A2(n_173),
.B1(n_196),
.B2(n_189),
.Y(n_253)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_75),
.B1(n_77),
.B2(n_66),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_188),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_139),
.B1(n_140),
.B2(n_149),
.Y(n_226)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_SL g191 ( 
.A1(n_156),
.A2(n_27),
.B(n_28),
.C(n_35),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_191),
.A2(n_197),
.B1(n_215),
.B2(n_216),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_124),
.B(n_35),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_134),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_104),
.C(n_77),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_195),
.C(n_201),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_141),
.B(n_66),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_151),
.B(n_65),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_129),
.A2(n_145),
.B1(n_151),
.B2(n_137),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_209),
.Y(n_228)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_198),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_131),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_115),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_2),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_203),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_204),
.Y(n_238)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_206),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_135),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

NAND2x1_ASAP7_75t_L g210 ( 
.A(n_136),
.B(n_48),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_149),
.B(n_132),
.Y(n_230)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_111),
.B(n_2),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_214),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_135),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_166),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_145),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_136),
.B(n_48),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_144),
.C(n_146),
.Y(n_251)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_142),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_219),
.B(n_254),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_180),
.A2(n_165),
.B1(n_109),
.B2(n_146),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_206),
.B1(n_211),
.B2(n_183),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_230),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_153),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_248),
.C(n_250),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_246),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_182),
.B(n_208),
.C(n_172),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_117),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_217),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_182),
.B(n_143),
.C(n_140),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_210),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_183),
.A2(n_126),
.B1(n_155),
.B2(n_130),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_253),
.B1(n_176),
.B2(n_217),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_170),
.B(n_144),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_257),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_258),
.B(n_254),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_230),
.A2(n_217),
.B(n_177),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_259),
.A2(n_274),
.B(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_261),
.A2(n_267),
.B1(n_273),
.B2(n_278),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_188),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_241),
.Y(n_297)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_203),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_221),
.A2(n_192),
.B1(n_195),
.B2(n_191),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_284),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_221),
.A2(n_195),
.B1(n_191),
.B2(n_174),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_185),
.B1(n_217),
.B2(n_187),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_276),
.B1(n_285),
.B2(n_233),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_195),
.B1(n_165),
.B2(n_194),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_193),
.B1(n_201),
.B2(n_155),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_220),
.A2(n_225),
.B(n_228),
.Y(n_274)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_201),
.B1(n_207),
.B2(n_205),
.Y(n_276)
);

OAI21x1_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_251),
.B(n_245),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_224),
.A2(n_130),
.B1(n_128),
.B2(n_126),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_236),
.A2(n_214),
.B1(n_218),
.B2(n_184),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_228),
.A2(n_210),
.B(n_199),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_282),
.Y(n_293)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

AOI32xp33_ASAP7_75t_L g282 ( 
.A1(n_220),
.A2(n_202),
.A3(n_179),
.B1(n_209),
.B2(n_133),
.Y(n_282)
);

AO22x1_ASAP7_75t_L g283 ( 
.A1(n_237),
.A2(n_199),
.B1(n_171),
.B2(n_214),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_251),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_228),
.A2(n_128),
.B1(n_186),
.B2(n_190),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_224),
.A2(n_175),
.B1(n_178),
.B2(n_143),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_219),
.B1(n_245),
.B2(n_243),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_289),
.A2(n_281),
.B1(n_287),
.B2(n_261),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g350 ( 
.A1(n_290),
.A2(n_276),
.B(n_278),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_243),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_291),
.B(n_299),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_296),
.A2(n_313),
.B1(n_268),
.B2(n_269),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_297),
.B(n_272),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_298),
.A2(n_315),
.B(n_259),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_262),
.Y(n_299)
);

CKINVDCx12_ASAP7_75t_R g300 ( 
.A(n_282),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_300),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_301),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_250),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_311),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_248),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_317),
.C(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_280),
.Y(n_329)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_285),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_261),
.A2(n_229),
.B1(n_242),
.B2(n_244),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_265),
.B(n_242),
.C(n_238),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_286),
.C(n_277),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_264),
.A2(n_274),
.B(n_280),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_265),
.B(n_246),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_234),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_257),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_320),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_327),
.C(n_334),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_277),
.C(n_258),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_331),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_330),
.B(n_342),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_271),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_271),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_332),
.B(n_339),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_317),
.C(n_313),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_288),
.A2(n_270),
.B1(n_277),
.B2(n_275),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_336),
.A2(n_345),
.B1(n_310),
.B2(n_294),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_337),
.A2(n_347),
.B(n_304),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_288),
.A2(n_270),
.B1(n_264),
.B2(n_275),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_338),
.A2(n_296),
.B1(n_305),
.B2(n_301),
.Y(n_353)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_315),
.A2(n_264),
.B(n_268),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_318),
.B(n_273),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_351),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_284),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_302),
.B(n_260),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_346),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_264),
.B1(n_276),
.B2(n_263),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_292),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_302),
.B(n_238),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_350),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_304),
.A2(n_279),
.B(n_284),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_349),
.A2(n_293),
.B(n_303),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_298),
.B(n_227),
.C(n_222),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_297),
.B(n_283),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_352),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_353),
.A2(n_354),
.B1(n_363),
.B2(n_367),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_330),
.A2(n_301),
.B1(n_305),
.B2(n_289),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_356),
.A2(n_381),
.B(n_380),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_344),
.Y(n_357)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_358),
.A2(n_366),
.B1(n_369),
.B2(n_372),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_359),
.A2(n_375),
.B(n_380),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_338),
.A2(n_293),
.B1(n_316),
.B2(n_294),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_320),
.A2(n_316),
.B1(n_303),
.B2(n_312),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_336),
.A2(n_316),
.B1(n_319),
.B2(n_283),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_345),
.A2(n_247),
.B1(n_231),
.B2(n_222),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_368),
.A2(n_376),
.B1(n_382),
.B2(n_383),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_344),
.A2(n_247),
.B1(n_231),
.B2(n_222),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_331),
.A2(n_247),
.B1(n_231),
.B2(n_235),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_347),
.A2(n_227),
.B(n_232),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_332),
.A2(n_235),
.B1(n_232),
.B2(n_239),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_322),
.B(n_144),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_384),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_342),
.A2(n_235),
.B1(n_198),
.B2(n_239),
.Y(n_379)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_379),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_337),
.A2(n_232),
.B(n_239),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_120),
.B(n_142),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_352),
.A2(n_132),
.B1(n_154),
.B2(n_255),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_349),
.A2(n_255),
.B1(n_108),
.B2(n_133),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_322),
.B(n_255),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_334),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_394),
.Y(n_422)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_361),
.Y(n_386)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_386),
.Y(n_417)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_354),
.B(n_323),
.Y(n_391)
);

XNOR2x1_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_402),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_362),
.B(n_323),
.C(n_340),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_406),
.C(n_353),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_341),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_327),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_400),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_365),
.B(n_333),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_396),
.B(n_397),
.Y(n_431)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_327),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_399),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_351),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_329),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_405),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_355),
.B(n_333),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_404),
.A2(n_381),
.B(n_374),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_371),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_355),
.B(n_351),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_360),
.A2(n_326),
.B1(n_328),
.B2(n_321),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_407),
.A2(n_390),
.B1(n_360),
.B2(n_358),
.Y(n_415)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_408),
.A2(n_369),
.B1(n_379),
.B2(n_382),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_357),
.B(n_348),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_409),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_373),
.B(n_343),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_411),
.Y(n_439)
);

INVx3_ASAP7_75t_SL g413 ( 
.A(n_375),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_413),
.B(n_414),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_373),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_415),
.A2(n_419),
.B1(n_420),
.B2(n_433),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_390),
.A2(n_364),
.B1(n_363),
.B2(n_378),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_394),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_403),
.Y(n_424)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

FAx1_ASAP7_75t_SL g425 ( 
.A(n_393),
.B(n_378),
.CI(n_326),
.CON(n_425),
.SN(n_425)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_427),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_395),
.B(n_356),
.C(n_359),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_404),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_335),
.Y(n_429)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_429),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_387),
.A2(n_367),
.B1(n_374),
.B2(n_368),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_430),
.A2(n_387),
.B1(n_392),
.B2(n_410),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_407),
.A2(n_366),
.B1(n_339),
.B2(n_383),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_412),
.A2(n_339),
.B(n_325),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_437),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_385),
.B(n_346),
.C(n_325),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_391),
.B(n_324),
.C(n_376),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_402),
.C(n_400),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_440),
.A2(n_462),
.B1(n_430),
.B2(n_392),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_449),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_416),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_406),
.C(n_398),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_446),
.B(n_448),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_434),
.C(n_438),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_429),
.Y(n_450)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_434),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_452),
.B(n_456),
.Y(n_475)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_417),
.Y(n_453)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_418),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_458),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_399),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_388),
.C(n_413),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_457),
.B(n_460),
.C(n_426),
.Y(n_464)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_432),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_431),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_424),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_388),
.C(n_426),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_416),
.B(n_412),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_428),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_324),
.Y(n_462)
);

INVx11_ASAP7_75t_L g463 ( 
.A(n_461),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_463),
.A2(n_480),
.B1(n_425),
.B2(n_456),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_473),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_448),
.C(n_449),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_467),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_440),
.A2(n_421),
.B1(n_415),
.B2(n_419),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_441),
.Y(n_468)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_477),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_435),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_321),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_444),
.A2(n_442),
.B(n_445),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_454),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_451),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_443),
.A2(n_425),
.B(n_433),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_482),
.A2(n_255),
.B(n_133),
.Y(n_494)
);

XNOR2x1_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_473),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_470),
.B(n_452),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_489),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_500),
.Y(n_505)
);

INVx6_ASAP7_75t_L g487 ( 
.A(n_481),
.Y(n_487)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_487),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_372),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_478),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_491),
.B(n_495),
.Y(n_514)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_492),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_494),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_471),
.A2(n_108),
.B1(n_5),
.B2(n_6),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g496 ( 
.A(n_480),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_496),
.B(n_475),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_468),
.B(n_2),
.Y(n_497)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_469),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_499)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_499),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_477),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_500)
);

INVxp33_ASAP7_75t_L g516 ( 
.A(n_502),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_474),
.Y(n_503)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_503),
.Y(n_521)
);

XNOR2x1_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_464),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_504),
.A2(n_510),
.B(n_483),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_493),
.A2(n_463),
.B(n_474),
.Y(n_509)
);

AOI31xp33_ASAP7_75t_L g524 ( 
.A1(n_509),
.A2(n_512),
.A3(n_10),
.B(n_11),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_488),
.A2(n_475),
.B(n_476),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_483),
.B(n_7),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_498),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_487),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_517),
.B(n_518),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_493),
.Y(n_518)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_519),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_520),
.A2(n_522),
.B1(n_524),
.B2(n_525),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_495),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_513),
.B(n_500),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_526),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_10),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_10),
.Y(n_526)
);

AOI21x1_ASAP7_75t_L g527 ( 
.A1(n_521),
.A2(n_509),
.B(n_505),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_531),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_516),
.A2(n_505),
.B(n_507),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_502),
.C(n_511),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_10),
.Y(n_537)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_533),
.A2(n_508),
.B(n_11),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_536),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_529),
.B(n_528),
.C(n_530),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_12),
.C(n_10),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_538),
.A2(n_535),
.B(n_534),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_539),
.B1(n_11),
.B2(n_12),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_12),
.B(n_535),
.Y(n_542)
);


endmodule