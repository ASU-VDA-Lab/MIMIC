module fake_jpeg_14549_n_360 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_360);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_14),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_0),
.B(n_1),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_33),
.B(n_43),
.C(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_56),
.Y(n_75)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_38),
.B1(n_30),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_69),
.A2(n_96),
.B1(n_94),
.B2(n_74),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_30),
.B1(n_38),
.B2(n_41),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_87),
.B1(n_33),
.B2(n_26),
.Y(n_115)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_72),
.Y(n_118)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_26),
.B(n_27),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_91),
.Y(n_116)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_41),
.B1(n_30),
.B2(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_100),
.Y(n_124)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_42),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_48),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_101),
.A2(n_102),
.B(n_109),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_0),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_58),
.C(n_45),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_98),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_0),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_46),
.B1(n_57),
.B2(n_43),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_61),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_126),
.Y(n_138)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_80),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_139)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_120),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_65),
.B1(n_21),
.B2(n_31),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_93),
.A2(n_63),
.B1(n_53),
.B2(n_66),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_21),
.B1(n_31),
.B2(n_42),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_0),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_45),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_68),
.B1(n_82),
.B2(n_86),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_45),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_132),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_73),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_85),
.A2(n_40),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_137),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_119),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_143),
.C(n_123),
.Y(n_173)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_112),
.B(n_81),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_150),
.B1(n_154),
.B2(n_129),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_79),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

CKINVDCx12_ASAP7_75t_R g154 ( 
.A(n_108),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_156),
.A2(n_158),
.B1(n_85),
.B2(n_67),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_22),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_102),
.Y(n_180)
);

OAI22x1_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_101),
.B1(n_110),
.B2(n_130),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_155),
.B1(n_143),
.B2(n_109),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_106),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_172),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_98),
.B1(n_103),
.B2(n_107),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_167),
.A2(n_96),
.B1(n_68),
.B2(n_160),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_102),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_180),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_103),
.B1(n_86),
.B2(n_111),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_179),
.B1(n_145),
.B2(n_159),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_163),
.A2(n_107),
.B1(n_67),
.B2(n_132),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_126),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_147),
.A2(n_109),
.B1(n_126),
.B2(n_40),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_155),
.B(n_138),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_197),
.B1(n_180),
.B2(n_139),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_193),
.B(n_202),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_196),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_136),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_171),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_198),
.B1(n_175),
.B2(n_158),
.Y(n_223)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_162),
.A3(n_163),
.B1(n_158),
.B2(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_135),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_164),
.A2(n_182),
.B1(n_174),
.B2(n_165),
.Y(n_197)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_134),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_162),
.B(n_156),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_217),
.B1(n_188),
.B2(n_149),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_207),
.B(n_153),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_172),
.C(n_166),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_189),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_213),
.A2(n_221),
.B(n_222),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_169),
.C(n_137),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_167),
.B1(n_177),
.B2(n_179),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_215),
.A2(n_224),
.B1(n_198),
.B2(n_202),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_190),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_216),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_184),
.B1(n_193),
.B2(n_199),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_134),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_175),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_168),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_221),
.B1(n_206),
.B2(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_186),
.A2(n_158),
.B1(n_176),
.B2(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_236),
.B1(n_241),
.B2(n_209),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_186),
.B(n_185),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_244),
.B(n_219),
.Y(n_261)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_234),
.A2(n_237),
.B(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_235),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_220),
.B(n_204),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_144),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_214),
.C(n_224),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_178),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_242),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_206),
.A2(n_142),
.B1(n_140),
.B2(n_104),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_178),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_205),
.Y(n_243)
);

XNOR2x2_ASAP7_75t_SL g244 ( 
.A(n_203),
.B(n_128),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_134),
.B1(n_118),
.B2(n_178),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_245),
.A2(n_49),
.B1(n_128),
.B2(n_34),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_247),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_207),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_251),
.B(n_271),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_256),
.C(n_259),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_225),
.C(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_215),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_245),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_268),
.B1(n_237),
.B2(n_240),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_153),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_269),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_231),
.B(n_34),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_241),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_266),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_227),
.A2(n_34),
.B1(n_2),
.B2(n_3),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_242),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_236),
.B(n_35),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_287),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_226),
.C(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_285),
.C(n_290),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_259),
.B(n_248),
.CI(n_229),
.CON(n_280),
.SN(n_280)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_280),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_281),
.Y(n_300)
);

AO22x1_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_249),
.B1(n_244),
.B2(n_247),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_283),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_254),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_266),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_269),
.C(n_255),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_244),
.B1(n_243),
.B2(n_234),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_267),
.B(n_240),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_262),
.B(n_270),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_233),
.C(n_45),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_264),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_298),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_289),
.A2(n_262),
.B(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_294),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_257),
.B1(n_268),
.B2(n_252),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_303),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_252),
.B(n_233),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_277),
.B1(n_290),
.B2(n_9),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_267),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_306),
.C(n_280),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_272),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_275),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_274),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_35),
.C(n_23),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_302),
.B(n_278),
.CI(n_286),
.CON(n_307),
.SN(n_307)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_309),
.C(n_310),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_280),
.C(n_283),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_284),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_320),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_35),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_298),
.B1(n_291),
.B2(n_11),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_316),
.A2(n_305),
.B1(n_296),
.B2(n_300),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_325),
.B(n_326),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_312),
.B(n_299),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_314),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_307),
.A2(n_8),
.B(n_10),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_11),
.B(n_13),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_35),
.C(n_23),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_317),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_321),
.B(n_310),
.Y(n_332)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_332),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_334),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_322),
.B(n_308),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_335),
.A2(n_336),
.B(n_338),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_317),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_327),
.Y(n_347)
);

INVx11_ASAP7_75t_L g338 ( 
.A(n_323),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_340),
.A2(n_16),
.B(n_17),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_13),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_328),
.C(n_330),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_343),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_324),
.C(n_329),
.Y(n_343)
);

AOI21x1_ASAP7_75t_SL g352 ( 
.A1(n_347),
.A2(n_348),
.B(n_16),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_345),
.B(n_338),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_349),
.A2(n_350),
.B(n_352),
.Y(n_354)
);

NAND3xp33_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_334),
.C(n_18),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_344),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_353),
.A2(n_346),
.B(n_354),
.Y(n_355)
);

AO21x1_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_18),
.B(n_19),
.Y(n_356)
);

AOI311xp33_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_18),
.A3(n_19),
.B(n_20),
.C(n_22),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_19),
.B(n_20),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_22),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_359),
.B(n_36),
.Y(n_360)
);


endmodule