module real_aes_7904_n_15 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_15);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_15;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR2xp33_ASAP7_75t_R g22 ( .A(n_0), .B(n_23), .Y(n_22) );
NAND2xp33_ASAP7_75t_SL g36 ( .A(n_0), .B(n_37), .Y(n_36) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_1), .B(n_19), .Y(n_18) );
NOR2xp33_ASAP7_75t_R g42 ( .A(n_1), .B(n_14), .Y(n_42) );
AOI322xp5_ASAP7_75t_SL g43 ( .A1(n_1), .A2(n_5), .A3(n_8), .B1(n_11), .B2(n_20), .C1(n_44), .C2(n_48), .Y(n_43) );
CKINVDCx20_ASAP7_75t_R g47 ( .A(n_1), .Y(n_47) );
NAND2xp33_ASAP7_75t_SL g49 ( .A(n_1), .B(n_46), .Y(n_49) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_2), .Y(n_28) );
NOR3xp33_ASAP7_75t_SL g26 ( .A(n_3), .B(n_9), .C(n_27), .Y(n_26) );
NOR2xp33_ASAP7_75t_R g20 ( .A(n_4), .B(n_21), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g41 ( .A(n_4), .Y(n_41) );
CKINVDCx20_ASAP7_75t_R g31 ( .A(n_6), .Y(n_31) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_7), .Y(n_27) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_10), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_12), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_12), .B(n_34), .Y(n_33) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_13), .Y(n_23) );
NAND4xp25_ASAP7_75t_SL g21 ( .A(n_14), .B(n_22), .C(n_24), .D(n_25), .Y(n_21) );
OAI221xp5_ASAP7_75t_R g15 ( .A1(n_16), .A2(n_17), .B1(n_29), .B2(n_32), .C(n_43), .Y(n_15) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
CKINVDCx16_ASAP7_75t_R g19 ( .A(n_20), .Y(n_19) );
NOR2xp33_ASAP7_75t_R g46 ( .A(n_21), .B(n_41), .Y(n_46) );
NAND2xp33_ASAP7_75t_SL g40 ( .A(n_23), .B(n_25), .Y(n_40) );
AND2x2_ASAP7_75t_L g25 ( .A(n_26), .B(n_28), .Y(n_25) );
INVx1_ASAP7_75t_L g29 ( .A(n_30), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
CKINVDCx16_ASAP7_75t_R g32 ( .A(n_33), .Y(n_32) );
NAND2xp33_ASAP7_75t_SL g34 ( .A(n_35), .B(n_42), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_36), .Y(n_35) );
CKINVDCx20_ASAP7_75t_R g37 ( .A(n_38), .Y(n_37) );
NAND2xp33_ASAP7_75t_SL g38 ( .A(n_39), .B(n_41), .Y(n_38) );
CKINVDCx20_ASAP7_75t_R g39 ( .A(n_40), .Y(n_39) );
INVx1_ASAP7_75t_SL g44 ( .A(n_45), .Y(n_44) );
NAND2xp33_ASAP7_75t_SL g45 ( .A(n_46), .B(n_47), .Y(n_45) );
CKINVDCx14_ASAP7_75t_R g48 ( .A(n_49), .Y(n_48) );
endmodule