module real_jpeg_21562_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_52),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_52),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_2),
.A2(n_35),
.B1(n_43),
.B2(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_2),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_3),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_133),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_133),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_3),
.A2(n_43),
.B1(n_51),
.B2(n_133),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_4),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_165),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_4),
.A2(n_43),
.B1(n_51),
.B2(n_165),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_165),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_6),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_6),
.A2(n_124),
.B(n_172),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_6),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_201)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_8),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_159),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_159),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_8),
.A2(n_43),
.B1(n_51),
.B2(n_159),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_9),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_9),
.A2(n_14),
.B(n_47),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_9),
.A2(n_43),
.B1(n_51),
.B2(n_163),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_9),
.A2(n_79),
.B1(n_218),
.B2(n_219),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_9),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_9),
.B(n_27),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_9),
.A2(n_27),
.B(n_245),
.Y(n_249)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_11),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_11),
.A2(n_43),
.B1(n_51),
.B2(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_63),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_13),
.A2(n_32),
.B1(n_43),
.B2(n_51),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_32),
.B1(n_46),
.B2(n_47),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_14),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_43),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_15),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_111),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_109),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_92),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_19),
.B(n_92),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_66),
.C(n_75),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_20),
.B(n_66),
.CI(n_75),
.CON(n_137),
.SN(n_137)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_38),
.B2(n_39),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_21),
.A2(n_22),
.B1(n_94),
.B2(n_107),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_22),
.B(n_40),
.C(n_54),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_33),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_23),
.A2(n_28),
.B1(n_88),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_23),
.A2(n_88),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_23),
.B(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_23),
.A2(n_88),
.B1(n_132),
.B2(n_178),
.Y(n_289)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_25),
.B(n_30),
.C(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_24),
.B(n_90),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_24),
.A2(n_36),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_25),
.B(n_27),
.Y(n_169)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_26),
.A2(n_37),
.B1(n_162),
.B2(n_169),
.Y(n_168)
);

AOI32xp33_ASAP7_75t_L g244 ( 
.A1(n_26),
.A2(n_43),
.A3(n_58),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_27),
.A2(n_57),
.B(n_59),
.C(n_60),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_57),
.Y(n_59)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g162 ( 
.A(n_30),
.B(n_163),
.CON(n_162),
.SN(n_162)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_53),
.B2(n_54),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_40),
.A2(n_41),
.B1(n_99),
.B2(n_105),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_49),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_42),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_42),
.A2(n_45),
.B1(n_84),
.B2(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_42),
.A2(n_49),
.B(n_85),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_42),
.A2(n_45),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_42),
.A2(n_45),
.B1(n_214),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_42),
.A2(n_45),
.B1(n_236),
.B2(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_42),
.A2(n_70),
.B(n_252),
.Y(n_267)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_45),
.A2(n_72),
.B(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_45),
.B(n_163),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_46),
.B(n_224),
.Y(n_223)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_80),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_48),
.A2(n_51),
.B(n_163),
.C(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_71),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g246 ( 
.A(n_51),
.B(n_57),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B(n_64),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_55),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_55),
.A2(n_101),
.B(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_55),
.A2(n_64),
.B(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_60),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_56),
.A2(n_60),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_56),
.A2(n_60),
.B1(n_158),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_56),
.A2(n_60),
.B1(n_190),
.B2(n_249),
.Y(n_248)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_60),
.A2(n_68),
.B(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_60),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_65),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_86),
.B(n_87),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_77),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_86),
.B1(n_87),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_78),
.A2(n_83),
.B1(n_86),
.B2(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B(n_81),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_79),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_79),
.A2(n_148),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_79),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_79),
.A2(n_204),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_79),
.A2(n_126),
.B(n_206),
.Y(n_237)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_80),
.B(n_125),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_80),
.B(n_163),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_82),
.A2(n_150),
.B(n_202),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_83),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_91),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_132),
.B(n_134),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_108),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B1(n_98),
.B2(n_106),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_102),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_138),
.B(n_315),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_137),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_113),
.B(n_137),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_119),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_114),
.B(n_118),
.Y(n_313)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_119),
.A2(n_120),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_130),
.C(n_135),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_121),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_128),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_122),
.B(n_128),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_130),
.A2(n_131),
.B1(n_135),
.B2(n_136),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_137),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_309),
.B(n_314),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_297),
.B(n_308),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_194),
.B(n_276),
.C(n_296),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_183),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_142),
.B(n_183),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_166),
.B2(n_182),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_145),
.B(n_153),
.C(n_182),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_146),
.B(n_152),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_151),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_161),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_161),
.B(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_167),
.B(n_175),
.C(n_180),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_170),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_184),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_188),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_192),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_189),
.B(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_191),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_275),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_269),
.B(n_274),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_257),
.B(n_268),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_239),
.B(n_256),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_227),
.B(n_238),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_215),
.B(n_226),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_207),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_211),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_221),
.B(n_225),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_229),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_235),
.C(n_237),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_241),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_247),
.B1(n_254),
.B2(n_255),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_242),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_248),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_253),
.C(n_254),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_266),
.C(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_278),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_294),
.B2(n_295),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_284),
.C(n_295),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_293),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_291),
.C(n_293),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_307),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_305),
.C(n_307),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);


endmodule