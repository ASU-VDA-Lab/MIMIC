module fake_ariane_544_n_1781 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1781);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1781;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g155 ( 
.A(n_15),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_29),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_8),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_91),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_76),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_20),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_100),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_7),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_52),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_38),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_85),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_8),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_110),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_4),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_45),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_132),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_34),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_82),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_35),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_37),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_5),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_101),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_77),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_13),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_14),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_29),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_41),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_10),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_45),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_19),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_11),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_65),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_80),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_20),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_60),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_149),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_49),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_4),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_51),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_135),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_87),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_96),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_84),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_58),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_38),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_6),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_10),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_56),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_66),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_55),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_30),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_147),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_22),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_34),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_92),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_61),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_126),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_63),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_108),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_114),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_30),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_112),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_41),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_59),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_48),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_130),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_74),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_31),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_106),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_116),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_28),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_121),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_1),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_99),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_136),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_103),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_26),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_28),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_105),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_42),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_151),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_19),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_98),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_128),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_107),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_17),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_89),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_62),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_129),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_12),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_64),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_113),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_72),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_24),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_18),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_68),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_36),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_51),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_32),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_15),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_26),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_21),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_90),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_54),
.Y(n_276)
);

BUFx8_ASAP7_75t_SL g277 ( 
.A(n_40),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_146),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_83),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_111),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_3),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_145),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_18),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_134),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_46),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_123),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_102),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_22),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_53),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_69),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_75),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_88),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_115),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_25),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_37),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_125),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_16),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_94),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_17),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_139),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_52),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_12),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_1),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_50),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_0),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_32),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_277),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_267),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_159),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_178),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_157),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_225),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_160),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_165),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_159),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_213),
.B(n_2),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_165),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_225),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_233),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_225),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_163),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_225),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_181),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_170),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_249),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_191),
.B(n_2),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_225),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_190),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_191),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_233),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_209),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_170),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_209),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_210),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_192),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_210),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_263),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_193),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_263),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_259),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_259),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_291),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_155),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_166),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_195),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_249),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_291),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_156),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_170),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_198),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_204),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_236),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_175),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_182),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_156),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_164),
.B(n_3),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_206),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_183),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_184),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_215),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_187),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_289),
.B(n_6),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_196),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_270),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_174),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_270),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_166),
.B(n_7),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_197),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_201),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_297),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_236),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_289),
.B(n_9),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_207),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_217),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_222),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_221),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_251),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_262),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_281),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_283),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_297),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_309),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_313),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_320),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_322),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_275),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_327),
.B(n_162),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_318),
.A2(n_306),
.B1(n_374),
.B2(n_364),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_335),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_336),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_338),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_339),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_339),
.B(n_167),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_341),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_341),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_312),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_348),
.B(n_168),
.Y(n_413)
);

AND2x6_ASAP7_75t_L g414 ( 
.A(n_358),
.B(n_174),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_355),
.B(n_162),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_355),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_360),
.B(n_205),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_361),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_314),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_365),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_323),
.B(n_162),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_325),
.B(n_296),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_370),
.B(n_173),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_370),
.A2(n_179),
.B(n_176),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_375),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_375),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_378),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_330),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_378),
.B(n_186),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_379),
.B(n_231),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_379),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_380),
.B(n_218),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_380),
.B(n_202),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_381),
.B(n_218),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_337),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_316),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_328),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_369),
.Y(n_452)
);

AO21x2_ASAP7_75t_L g453 ( 
.A1(n_433),
.A2(n_230),
.B(n_219),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_386),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_400),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_386),
.Y(n_456)
);

AO22x2_ASAP7_75t_L g457 ( 
.A1(n_417),
.A2(n_351),
.B1(n_326),
.B2(n_334),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_340),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_347),
.Y(n_460)
);

AO21x2_ASAP7_75t_L g461 ( 
.A1(n_433),
.A2(n_252),
.B(n_238),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_385),
.Y(n_463)
);

OAI22xp33_ASAP7_75t_L g464 ( 
.A1(n_399),
.A2(n_306),
.B1(n_373),
.B2(n_354),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_427),
.B(n_352),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_385),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_385),
.Y(n_467)
);

OAI21xp33_ASAP7_75t_SL g468 ( 
.A1(n_399),
.A2(n_301),
.B(n_288),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_399),
.A2(n_315),
.B1(n_311),
.B2(n_319),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_427),
.B(n_353),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_409),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_427),
.B(n_359),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_423),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_385),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_417),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_427),
.B(n_362),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_387),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_427),
.B(n_429),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_389),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_443),
.B(n_376),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_SL g485 ( 
.A(n_411),
.B(n_377),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_439),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_441),
.A2(n_445),
.B1(n_443),
.B2(n_414),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_439),
.B(n_449),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_428),
.B(n_303),
.C(n_261),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_394),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_441),
.A2(n_315),
.B1(n_346),
.B2(n_214),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_443),
.B(n_236),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_394),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_387),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_445),
.B(n_172),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_445),
.B(n_218),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_450),
.B(n_308),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_396),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_396),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_393),
.B(n_177),
.Y(n_504)
);

BUFx10_ASAP7_75t_L g505 ( 
.A(n_430),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_393),
.B(n_227),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_429),
.B(n_254),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_398),
.B(n_256),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_400),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_387),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_423),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_450),
.A2(n_234),
.B1(n_172),
.B2(n_244),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_449),
.B(n_430),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_411),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_449),
.B(n_169),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_422),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_387),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_R g521 ( 
.A(n_449),
.B(n_310),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_449),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_390),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_423),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_398),
.B(n_441),
.Y(n_525)
);

NOR3xp33_ASAP7_75t_L g526 ( 
.A(n_449),
.B(n_294),
.C(n_244),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_423),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_390),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_398),
.B(n_280),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_423),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_428),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_441),
.B(n_169),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_423),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_423),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_441),
.B(n_205),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_390),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_390),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_395),
.Y(n_540)
);

OR2x6_ASAP7_75t_L g541 ( 
.A(n_441),
.B(n_231),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_418),
.B(n_229),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_423),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_450),
.B(n_264),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_426),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_452),
.B(n_171),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_391),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_428),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_426),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_391),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_426),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_452),
.B(n_171),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_426),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_426),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_450),
.B(n_452),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_418),
.B(n_229),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_428),
.B(n_180),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_413),
.B(n_180),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_428),
.B(n_293),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_426),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_391),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_392),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_414),
.A2(n_245),
.B1(n_243),
.B2(n_229),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_426),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_438),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_384),
.B(n_294),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_428),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_392),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_422),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_413),
.B(n_282),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_395),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_418),
.B(n_293),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_451),
.B(n_300),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_419),
.B(n_420),
.Y(n_577)
);

XNOR2x2_ASAP7_75t_L g578 ( 
.A(n_384),
.B(n_317),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_409),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_438),
.Y(n_580)
);

NAND3xp33_ASAP7_75t_L g581 ( 
.A(n_438),
.B(n_292),
.C(n_284),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_419),
.B(n_300),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_395),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_419),
.B(n_255),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_451),
.B(n_295),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_438),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_438),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_420),
.B(n_243),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_395),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_420),
.B(n_255),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_438),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_392),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_392),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_438),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_409),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_421),
.B(n_434),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_451),
.B(n_295),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_395),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_409),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_414),
.A2(n_245),
.B1(n_243),
.B2(n_232),
.Y(n_601)
);

BUFx12f_ASAP7_75t_SL g602 ( 
.A(n_497),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_486),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_522),
.B(n_414),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_599),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_455),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_493),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_513),
.A2(n_433),
.B(n_448),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_515),
.B(n_448),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_508),
.A2(n_414),
.B1(n_447),
.B2(n_435),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_463),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_486),
.B(n_438),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_466),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_454),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_502),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_466),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_577),
.A2(n_433),
.B(n_432),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_481),
.A2(n_414),
.B1(n_447),
.B2(n_434),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_467),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_454),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_460),
.B(n_448),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_459),
.B(n_421),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_456),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_456),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_477),
.B(n_421),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_455),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_483),
.B(n_447),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_493),
.B(n_321),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_477),
.B(n_434),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_488),
.B(n_435),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_458),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_533),
.B(n_446),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_574),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_542),
.B(n_557),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_505),
.B(n_435),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_533),
.B(n_446),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_467),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_542),
.B(n_436),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_505),
.B(n_446),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_574),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_505),
.B(n_446),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_458),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_497),
.B(n_332),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_505),
.B(n_446),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_583),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_455),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_557),
.B(n_436),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_588),
.B(n_436),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_510),
.B(n_432),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_588),
.B(n_395),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_531),
.B(n_440),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_462),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_516),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_533),
.B(n_549),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_462),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_473),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_573),
.B(n_446),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_533),
.B(n_446),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_473),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_525),
.B(n_446),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_544),
.B(n_446),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_475),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_464),
.A2(n_414),
.B1(n_442),
.B2(n_415),
.Y(n_664)
);

INVx5_ASAP7_75t_L g665 ( 
.A(n_537),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_468),
.A2(n_414),
.B1(n_442),
.B2(n_415),
.Y(n_666)
);

AOI22x1_ASAP7_75t_L g667 ( 
.A1(n_549),
.A2(n_415),
.B1(n_442),
.B2(n_437),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_476),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_475),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_480),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_496),
.B(n_440),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_549),
.B(n_415),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_487),
.B(n_444),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_549),
.B(n_416),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_SL g675 ( 
.A(n_468),
.B(n_342),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_570),
.B(n_416),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_480),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_482),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_570),
.B(n_416),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_570),
.B(n_416),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_496),
.B(n_444),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_482),
.Y(n_682)
);

OAI221xp5_ASAP7_75t_L g683 ( 
.A1(n_469),
.A2(n_299),
.B1(n_302),
.B2(n_304),
.C(n_305),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_496),
.B(n_424),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_496),
.B(n_424),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_578),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_541),
.A2(n_414),
.B1(n_442),
.B2(n_431),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_565),
.A2(n_414),
.B1(n_431),
.B2(n_425),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_511),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_514),
.B(n_305),
.C(n_299),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_476),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_504),
.B(n_424),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_506),
.B(n_424),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_484),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_583),
.B(n_425),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_589),
.B(n_425),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_569),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_SL g698 ( 
.A(n_465),
.B(n_302),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_499),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_583),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_484),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_540),
.B(n_425),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_490),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_479),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_540),
.B(n_559),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_570),
.B(n_431),
.Y(n_706)
);

NOR2xp67_ASAP7_75t_L g707 ( 
.A(n_499),
.B(n_431),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_589),
.B(n_437),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_556),
.B(n_437),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_575),
.B(n_437),
.Y(n_710)
);

BUFx5_ASAP7_75t_L g711 ( 
.A(n_513),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_569),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_578),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_582),
.B(n_397),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_534),
.B(n_397),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_470),
.B(n_397),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_521),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_546),
.B(n_403),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_541),
.B(n_407),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_490),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_541),
.A2(n_414),
.B1(n_403),
.B2(n_404),
.Y(n_721)
);

OR2x6_ASAP7_75t_SL g722 ( 
.A(n_485),
.B(n_304),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_511),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_479),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_601),
.A2(n_414),
.B1(n_406),
.B2(n_401),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_553),
.B(n_403),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_472),
.B(n_404),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_526),
.B(n_274),
.C(n_272),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_541),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_507),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_541),
.A2(n_404),
.B1(n_407),
.B2(n_410),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_495),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_478),
.B(n_410),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_491),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_517),
.B(n_224),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_491),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_494),
.Y(n_737)
);

INVx8_ASAP7_75t_L g738 ( 
.A(n_537),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_495),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_494),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_512),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_596),
.B(n_507),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_576),
.B(n_410),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_512),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_585),
.B(n_401),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_511),
.B(n_401),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_514),
.B(n_492),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_600),
.B(n_409),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_457),
.A2(n_298),
.B1(n_401),
.B2(n_402),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_598),
.B(n_343),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_558),
.A2(n_402),
.B(n_408),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_457),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_528),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_457),
.Y(n_754)
);

AO22x2_ASAP7_75t_L g755 ( 
.A1(n_457),
.A2(n_349),
.B1(n_344),
.B2(n_383),
.Y(n_755)
);

NAND2x1_ASAP7_75t_L g756 ( 
.A(n_500),
.B(n_402),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_528),
.B(n_402),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_528),
.B(n_412),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_500),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_471),
.B(n_600),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_560),
.B(n_405),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_501),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_584),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_501),
.B(n_405),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_503),
.A2(n_405),
.B(n_408),
.C(n_406),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_503),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_471),
.B(n_409),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_519),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_537),
.A2(n_405),
.B1(n_406),
.B2(n_408),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_590),
.B(n_406),
.Y(n_770)
);

OA21x2_ASAP7_75t_L g771 ( 
.A1(n_524),
.A2(n_408),
.B(n_412),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_537),
.B(n_412),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_650),
.B(n_537),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_609),
.A2(n_527),
.B(n_524),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_609),
.A2(n_532),
.B1(n_535),
.B2(n_552),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_661),
.A2(n_529),
.B(n_527),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_672),
.A2(n_536),
.B(n_529),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_617),
.A2(n_543),
.B(n_536),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_672),
.A2(n_545),
.B(n_543),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_603),
.B(n_738),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_717),
.B(n_489),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_707),
.B(n_537),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_618),
.B(n_242),
.C(n_239),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_602),
.B(n_350),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_606),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_635),
.A2(n_580),
.B(n_597),
.C(n_563),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_614),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_697),
.B(n_357),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_674),
.A2(n_679),
.B(n_676),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_615),
.B(n_366),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_650),
.B(n_537),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_652),
.B(n_519),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_652),
.B(n_523),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_674),
.A2(n_679),
.B(n_676),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_671),
.B(n_523),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_655),
.A2(n_550),
.B(n_545),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_654),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_690),
.B(n_253),
.C(n_248),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_655),
.A2(n_554),
.B(n_550),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_646),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_680),
.A2(n_563),
.B(n_554),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_671),
.B(n_530),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_760),
.A2(n_568),
.B(n_567),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_680),
.A2(n_568),
.B(n_567),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_695),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_622),
.B(n_530),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_760),
.A2(n_587),
.B(n_597),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_706),
.A2(n_587),
.B(n_594),
.Y(n_808)
);

BUFx4f_ASAP7_75t_L g809 ( 
.A(n_646),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_699),
.B(n_368),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_706),
.A2(n_580),
.B(n_594),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_747),
.A2(n_489),
.B1(n_591),
.B2(n_552),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_621),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_622),
.B(n_538),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_L g815 ( 
.A1(n_636),
.A2(n_257),
.B(n_266),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_624),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_623),
.A2(n_591),
.B(n_561),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_628),
.B(n_681),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_628),
.B(n_538),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_629),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_633),
.A2(n_535),
.B(n_566),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_644),
.B(n_372),
.Y(n_822)
);

O2A1O1Ixp5_ASAP7_75t_L g823 ( 
.A1(n_636),
.A2(n_561),
.B(n_532),
.C(n_535),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_630),
.B(n_539),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_630),
.B(n_539),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_633),
.A2(n_474),
.B(n_561),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_738),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_639),
.B(n_547),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_648),
.B(n_547),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_712),
.B(n_474),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_634),
.A2(n_555),
.B1(n_552),
.B2(n_474),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_608),
.A2(n_595),
.B(n_532),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_683),
.B(n_269),
.C(n_271),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_607),
.B(n_555),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_649),
.B(n_548),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_637),
.A2(n_555),
.B(n_566),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_695),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_634),
.A2(n_586),
.B1(n_566),
.B2(n_595),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_606),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_646),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_637),
.A2(n_586),
.B(n_593),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_659),
.A2(n_742),
.B(n_746),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_607),
.A2(n_586),
.B(n_593),
.C(n_564),
.Y(n_843)
);

BUFx4f_ASAP7_75t_L g844 ( 
.A(n_646),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_659),
.A2(n_461),
.B(n_453),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_685),
.A2(n_684),
.B(n_626),
.C(n_641),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_631),
.A2(n_548),
.B(n_592),
.C(n_551),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_611),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_700),
.B(n_471),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_700),
.B(n_471),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_700),
.B(n_729),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_651),
.B(n_551),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_605),
.B(n_412),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_641),
.B(n_562),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_619),
.A2(n_562),
.B(n_592),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_757),
.A2(n_461),
.B(n_453),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_627),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_750),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_702),
.B(n_564),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_763),
.B(n_471),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_631),
.A2(n_571),
.B(n_581),
.C(n_579),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_702),
.B(n_571),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_700),
.B(n_498),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_710),
.A2(n_600),
.B(n_579),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_658),
.A2(n_761),
.B(n_714),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_675),
.Y(n_866)
);

AOI22xp5_ASAP7_75t_L g867 ( 
.A1(n_705),
.A2(n_600),
.B1(n_579),
.B2(n_520),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_761),
.A2(n_581),
.B(n_422),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_715),
.A2(n_453),
.B(n_461),
.C(n_285),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_718),
.A2(n_600),
.B(n_579),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_755),
.B(n_409),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_673),
.B(n_692),
.Y(n_872)
);

BUFx12f_ASAP7_75t_L g873 ( 
.A(n_719),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_729),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_613),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_730),
.B(n_498),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_664),
.B(n_498),
.Y(n_877)
);

AOI33xp33_ASAP7_75t_L g878 ( 
.A1(n_749),
.A2(n_307),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.B3(n_21),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_647),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_625),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_705),
.A2(n_579),
.B(n_520),
.C(n_498),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_752),
.B(n_509),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_743),
.A2(n_498),
.B(n_520),
.C(n_161),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_632),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_738),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_664),
.A2(n_520),
.B1(n_158),
.B2(n_241),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_693),
.B(n_520),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_665),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_726),
.B(n_245),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_751),
.A2(n_572),
.B(n_518),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_748),
.A2(n_572),
.B(n_518),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_643),
.A2(n_737),
.B(n_678),
.C(n_694),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_765),
.A2(n_422),
.B(n_518),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_653),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_743),
.A2(n_240),
.B(n_188),
.C(n_189),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_748),
.A2(n_572),
.B(n_518),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_656),
.A2(n_9),
.B(n_23),
.C(n_24),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_657),
.A2(n_23),
.B(n_25),
.C(n_27),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_767),
.A2(n_572),
.B(n_518),
.Y(n_899)
);

O2A1O1Ixp5_ASAP7_75t_L g900 ( 
.A1(n_698),
.A2(n_422),
.B(n_31),
.C(n_33),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_660),
.B(n_185),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_722),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_754),
.B(n_199),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_758),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_627),
.B(n_509),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_663),
.A2(n_572),
.B1(n_518),
.B2(n_509),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_616),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_758),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_665),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_669),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_620),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_755),
.B(n_27),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_745),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_670),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_677),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_767),
.A2(n_572),
.B(n_509),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_612),
.B(n_268),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_682),
.A2(n_33),
.B(n_35),
.C(n_39),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_701),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_719),
.B(n_265),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_703),
.B(n_276),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_720),
.A2(n_39),
.B(n_40),
.C(n_42),
.Y(n_922)
);

BUFx4f_ASAP7_75t_L g923 ( 
.A(n_719),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_758),
.Y(n_924)
);

AOI33xp33_ASAP7_75t_L g925 ( 
.A1(n_734),
.A2(n_43),
.A3(n_44),
.B1(n_46),
.B2(n_47),
.B3(n_48),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_736),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_764),
.A2(n_509),
.B(n_237),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_740),
.A2(n_509),
.B1(n_290),
.B2(n_287),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_745),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_755),
.B(n_43),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_716),
.A2(n_226),
.B1(n_286),
.B2(n_279),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_638),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_759),
.B(n_247),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_686),
.B(n_44),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_770),
.A2(n_223),
.B(n_278),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_640),
.A2(n_228),
.B(n_260),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_762),
.B(n_246),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_647),
.B(n_235),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_668),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_766),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_731),
.B(n_250),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_689),
.B(n_723),
.Y(n_942)
);

CKINVDCx10_ASAP7_75t_R g943 ( 
.A(n_728),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_R g944 ( 
.A(n_735),
.B(n_200),
.Y(n_944)
);

NOR2xp67_ASAP7_75t_L g945 ( 
.A(n_716),
.B(n_203),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_727),
.B(n_258),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_662),
.A2(n_211),
.B(n_212),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_727),
.B(n_208),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_733),
.A2(n_205),
.B(n_216),
.C(n_50),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_733),
.B(n_47),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_604),
.A2(n_216),
.B(n_205),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_L g952 ( 
.A(n_728),
.B(n_49),
.C(n_53),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_610),
.A2(n_216),
.B(n_205),
.C(n_220),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_665),
.B(n_723),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_756),
.A2(n_696),
.B(n_708),
.Y(n_955)
);

NAND3xp33_ASAP7_75t_L g956 ( 
.A(n_666),
.B(n_216),
.C(n_422),
.Y(n_956)
);

AO21x1_ASAP7_75t_L g957 ( 
.A1(n_642),
.A2(n_220),
.B(n_194),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_691),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_665),
.B(n_422),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_704),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_645),
.A2(n_216),
.B(n_422),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_689),
.B(n_422),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_818),
.A2(n_753),
.B(n_667),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_810),
.B(n_713),
.Y(n_964)
);

OAI22x1_ASAP7_75t_L g965 ( 
.A1(n_912),
.A2(n_721),
.B1(n_687),
.B2(n_666),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_797),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_820),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_SL g968 ( 
.A(n_790),
.B(n_772),
.Y(n_968)
);

AO21x2_ASAP7_75t_L g969 ( 
.A1(n_856),
.A2(n_709),
.B(n_768),
.Y(n_969)
);

AND3x1_ASAP7_75t_SL g970 ( 
.A(n_943),
.B(n_422),
.C(n_220),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_788),
.B(n_753),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_929),
.B(n_739),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_865),
.A2(n_771),
.B(n_732),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_787),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_913),
.B(n_724),
.Y(n_975)
);

INVx5_ASAP7_75t_L g976 ( 
.A(n_780),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_SL g977 ( 
.A(n_902),
.B(n_422),
.C(n_711),
.Y(n_977)
);

CKINVDCx11_ASAP7_75t_R g978 ( 
.A(n_873),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_813),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_792),
.B(n_744),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_822),
.B(n_741),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_806),
.A2(n_771),
.B(n_688),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_950),
.A2(n_688),
.B(n_725),
.C(n_769),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_793),
.B(n_711),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_949),
.A2(n_725),
.B(n_771),
.C(n_711),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_858),
.B(n_784),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_814),
.A2(n_711),
.B(n_70),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_809),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_848),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_819),
.A2(n_711),
.B(n_71),
.Y(n_990)
);

OA22x2_ASAP7_75t_L g991 ( 
.A1(n_930),
.A2(n_711),
.B1(n_220),
.B2(n_194),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_809),
.Y(n_992)
);

AOI221xp5_ASAP7_75t_L g993 ( 
.A1(n_833),
.A2(n_220),
.B1(n_194),
.B2(n_78),
.C(n_79),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_844),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_795),
.A2(n_57),
.B(n_73),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_874),
.B(n_220),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_904),
.B(n_81),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_816),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_773),
.A2(n_220),
.B(n_194),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_923),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_946),
.A2(n_194),
.B1(n_97),
.B2(n_104),
.Y(n_1001)
);

OR2x6_ASAP7_75t_L g1002 ( 
.A(n_904),
.B(n_95),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_923),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_934),
.B(n_194),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_802),
.A2(n_117),
.B(n_119),
.Y(n_1005)
);

INVx6_ASAP7_75t_L g1006 ( 
.A(n_780),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_791),
.A2(n_194),
.B(n_124),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_948),
.A2(n_919),
.B1(n_940),
.B2(n_926),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_952),
.A2(n_120),
.B1(n_137),
.B2(n_141),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_SL g1010 ( 
.A1(n_878),
.A2(n_142),
.B(n_143),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_774),
.A2(n_144),
.B(n_153),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_866),
.B(n_889),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_844),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_892),
.A2(n_846),
.B(n_815),
.C(n_872),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_875),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_897),
.A2(n_898),
.B(n_922),
.C(n_918),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_924),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_R g1018 ( 
.A(n_885),
.B(n_800),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_885),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_885),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_920),
.B(n_853),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_805),
.B(n_837),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_780),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_800),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_907),
.Y(n_1025)
);

AOI221xp5_ASAP7_75t_L g1026 ( 
.A1(n_783),
.A2(n_798),
.B1(n_894),
.B2(n_880),
.C(n_884),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_800),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_910),
.B(n_914),
.Y(n_1028)
);

OAI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_941),
.A2(n_915),
.B1(n_931),
.B2(n_886),
.Y(n_1029)
);

BUFx4f_ASAP7_75t_L g1030 ( 
.A(n_908),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_840),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_774),
.A2(n_887),
.B(n_859),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_895),
.A2(n_921),
.B(n_937),
.C(n_933),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_827),
.B(n_908),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_840),
.B(n_888),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_944),
.Y(n_1036)
);

NOR2xp67_ASAP7_75t_L g1037 ( 
.A(n_827),
.B(n_785),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_911),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_834),
.B(n_830),
.Y(n_1039)
);

INVx6_ASAP7_75t_L g1040 ( 
.A(n_871),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_932),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_824),
.B(n_825),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_939),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_945),
.B(n_781),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_901),
.A2(n_786),
.B(n_843),
.C(n_883),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_851),
.B(n_959),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_888),
.Y(n_1047)
);

INVx5_ASAP7_75t_L g1048 ( 
.A(n_888),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_958),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_879),
.A2(n_828),
.B1(n_829),
.B2(n_835),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_862),
.A2(n_842),
.B(n_864),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_960),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_854),
.A2(n_938),
.B1(n_852),
.B2(n_860),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_876),
.Y(n_1054)
);

NOR2x1_ASAP7_75t_R g1055 ( 
.A(n_959),
.B(n_782),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_909),
.B(n_782),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_909),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_842),
.A2(n_776),
.B(n_817),
.Y(n_1058)
);

AOI21xp33_ASAP7_75t_L g1059 ( 
.A1(n_903),
.A2(n_917),
.B(n_869),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_849),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_785),
.B(n_839),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_839),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_956),
.A2(n_877),
.B1(n_882),
.B2(n_812),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_863),
.Y(n_1064)
);

AOI21x1_ASAP7_75t_L g1065 ( 
.A1(n_856),
.A2(n_845),
.B(n_776),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_909),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_900),
.A2(n_881),
.B(n_847),
.C(n_823),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_789),
.A2(n_794),
.B(n_868),
.C(n_951),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_850),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_R g1070 ( 
.A(n_857),
.B(n_942),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_775),
.A2(n_953),
.B(n_789),
.C(n_794),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_954),
.B(n_951),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_857),
.B(n_867),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_817),
.A2(n_870),
.B(n_832),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_925),
.B(n_855),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_936),
.Y(n_1076)
);

BUFx12f_ASAP7_75t_L g1077 ( 
.A(n_954),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_893),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_935),
.B(n_947),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_R g1080 ( 
.A(n_962),
.B(n_957),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_838),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_955),
.B(n_831),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_947),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_779),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_928),
.A2(n_841),
.B1(n_811),
.B2(n_804),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_801),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_808),
.A2(n_861),
.B1(n_845),
.B2(n_955),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_905),
.Y(n_1088)
);

O2A1O1Ixp5_ASAP7_75t_SL g1089 ( 
.A1(n_778),
.A2(n_906),
.B(n_927),
.C(n_803),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_796),
.A2(n_799),
.B(n_807),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_777),
.A2(n_821),
.B1(n_826),
.B2(n_836),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_821),
.Y(n_1092)
);

AND3x1_ASAP7_75t_SL g1093 ( 
.A(n_826),
.B(n_836),
.C(n_777),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_961),
.B(n_927),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_R g1095 ( 
.A(n_961),
.B(n_891),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_891),
.B(n_896),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_896),
.B(n_899),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_899),
.B(n_916),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_916),
.B(n_890),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_890),
.B(n_486),
.Y(n_1100)
);

AND2x2_ASAP7_75t_SL g1101 ( 
.A(n_923),
.B(n_912),
.Y(n_1101)
);

NOR2xp67_ASAP7_75t_L g1102 ( 
.A(n_827),
.B(n_913),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_818),
.A2(n_609),
.B(n_865),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_818),
.A2(n_609),
.B(n_865),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_820),
.Y(n_1105)
);

INVx5_ASAP7_75t_L g1106 ( 
.A(n_780),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_818),
.A2(n_609),
.B(n_865),
.Y(n_1107)
);

BUFx4f_ASAP7_75t_L g1108 ( 
.A(n_780),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_810),
.B(n_486),
.Y(n_1109)
);

INVx6_ASAP7_75t_L g1110 ( 
.A(n_988),
.Y(n_1110)
);

AO32x2_ASAP7_75t_L g1111 ( 
.A1(n_1091),
.A2(n_1008),
.A3(n_1050),
.B1(n_1053),
.B2(n_1001),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_988),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1094),
.A2(n_1096),
.A3(n_1098),
.B(n_1058),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1105),
.B(n_986),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1109),
.B(n_964),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_989),
.Y(n_1117)
);

BUFx2_ASAP7_75t_R g1118 ( 
.A(n_1013),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_984),
.A2(n_1082),
.B(n_1032),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1012),
.B(n_1021),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_974),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_967),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_978),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1014),
.A2(n_1039),
.B(n_1100),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1051),
.A2(n_1074),
.B(n_1068),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_971),
.B(n_966),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_SL g1127 ( 
.A1(n_1010),
.A2(n_1016),
.B1(n_1075),
.B2(n_1029),
.C(n_1033),
.Y(n_1127)
);

AO32x2_ASAP7_75t_L g1128 ( 
.A1(n_1023),
.A2(n_1093),
.A3(n_1088),
.B1(n_1065),
.B2(n_1000),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1071),
.A2(n_1087),
.B(n_985),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_979),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_998),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_SL g1132 ( 
.A1(n_1045),
.A2(n_1067),
.B(n_1081),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_981),
.B(n_1101),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_1099),
.A2(n_1087),
.B(n_1090),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1036),
.Y(n_1135)
);

AO32x2_ASAP7_75t_L g1136 ( 
.A1(n_1003),
.A2(n_991),
.A3(n_969),
.B1(n_1092),
.B2(n_1010),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_987),
.A2(n_990),
.B(n_963),
.Y(n_1137)
);

INVx5_ASAP7_75t_L g1138 ( 
.A(n_988),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1038),
.Y(n_1139)
);

AOI21x1_ASAP7_75t_L g1140 ( 
.A1(n_973),
.A2(n_982),
.B(n_1097),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1059),
.A2(n_1044),
.B(n_1026),
.C(n_1007),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_1030),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1017),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1079),
.A2(n_983),
.B(n_1011),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1089),
.A2(n_999),
.B(n_1005),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1041),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_993),
.A2(n_1064),
.B(n_975),
.C(n_1084),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_992),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_994),
.B(n_976),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_972),
.B(n_968),
.Y(n_1150)
);

AO21x2_ASAP7_75t_L g1151 ( 
.A1(n_969),
.A2(n_1095),
.B(n_1080),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1049),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1086),
.A2(n_1061),
.B(n_996),
.C(n_1060),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_994),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1052),
.B(n_1022),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1030),
.B(n_1042),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_992),
.B(n_1004),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_980),
.A2(n_1072),
.B(n_1085),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_965),
.A2(n_1078),
.A3(n_1069),
.B(n_1054),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_995),
.A2(n_1063),
.B(n_1085),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1048),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1015),
.A2(n_1025),
.A3(n_1043),
.B(n_1062),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_997),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_992),
.B(n_1102),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_SL g1165 ( 
.A(n_1002),
.B(n_1108),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1040),
.A2(n_1083),
.B1(n_1002),
.B2(n_1073),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1057),
.A2(n_1037),
.B(n_1009),
.Y(n_1167)
);

AOI221x1_ASAP7_75t_L g1168 ( 
.A1(n_1057),
.A2(n_1031),
.B1(n_1027),
.B2(n_1066),
.C(n_1047),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1072),
.A2(n_1037),
.B(n_1108),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_SL g1170 ( 
.A1(n_1009),
.A2(n_1070),
.B(n_1102),
.C(n_1076),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_1072),
.A2(n_1040),
.A3(n_1019),
.B(n_977),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_1024),
.Y(n_1172)
);

CKINVDCx11_ASAP7_75t_R g1173 ( 
.A(n_1077),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_976),
.A2(n_1106),
.B(n_1006),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1056),
.A2(n_1034),
.B(n_1002),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_976),
.A2(n_1106),
.B(n_1048),
.C(n_1066),
.Y(n_1176)
);

O2A1O1Ixp5_ASAP7_75t_L g1177 ( 
.A1(n_1019),
.A2(n_970),
.B(n_1106),
.C(n_1006),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1027),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1056),
.A2(n_1034),
.B(n_1048),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_1020),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1055),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1034),
.A2(n_1056),
.B1(n_1046),
.B2(n_1020),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_1018),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_1035),
.A2(n_1046),
.B(n_1055),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_SL g1185 ( 
.A1(n_1047),
.A2(n_1066),
.B(n_1027),
.C(n_1031),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1020),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1031),
.A2(n_818),
.B1(n_515),
.B2(n_399),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1047),
.A2(n_1104),
.B(n_1103),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_966),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1014),
.A2(n_515),
.B(n_636),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1058),
.A2(n_1051),
.B(n_973),
.Y(n_1191)
);

AOI221x1_ASAP7_75t_L g1192 ( 
.A1(n_1059),
.A2(n_952),
.B1(n_1001),
.B2(n_755),
.C(n_1100),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1028),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1100),
.A2(n_515),
.B(n_1059),
.C(n_481),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_994),
.Y(n_1195)
);

NOR2xp67_ASAP7_75t_L g1196 ( 
.A(n_1048),
.B(n_1057),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1013),
.B(n_994),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1109),
.B(n_486),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1065),
.A2(n_1074),
.B(n_1058),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1109),
.A2(n_818),
.B1(n_515),
.B2(n_399),
.Y(n_1200)
);

OAI22x1_ASAP7_75t_L g1201 ( 
.A1(n_1109),
.A2(n_399),
.B1(n_930),
.B2(n_912),
.Y(n_1201)
);

CKINVDCx11_ASAP7_75t_R g1202 ( 
.A(n_966),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1203)
);

OR2x6_ASAP7_75t_L g1204 ( 
.A(n_1002),
.B(n_1056),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1109),
.B(n_486),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1109),
.B(n_486),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1058),
.A2(n_1051),
.B(n_973),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1100),
.A2(n_515),
.B(n_1059),
.C(n_481),
.Y(n_1209)
);

OR2x6_ASAP7_75t_L g1210 ( 
.A(n_1002),
.B(n_1056),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1109),
.Y(n_1211)
);

NAND2x1_ASAP7_75t_L g1212 ( 
.A(n_1034),
.B(n_785),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_994),
.Y(n_1215)
);

INVxp67_ASAP7_75t_SL g1216 ( 
.A(n_1064),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1100),
.A2(n_515),
.B(n_1059),
.C(n_481),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1218)
);

OAI22x1_ASAP7_75t_L g1219 ( 
.A1(n_1109),
.A2(n_399),
.B1(n_930),
.B2(n_912),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_966),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1014),
.A2(n_515),
.B(n_636),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1048),
.B(n_1057),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_966),
.Y(n_1223)
);

AO22x1_ASAP7_75t_L g1224 ( 
.A1(n_1109),
.A2(n_486),
.B1(n_747),
.B2(n_964),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1109),
.A2(n_818),
.B1(n_515),
.B2(n_399),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_967),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1058),
.A2(n_1051),
.B(n_973),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1058),
.A2(n_1051),
.B(n_973),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1014),
.A2(n_515),
.B(n_636),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_967),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1100),
.A2(n_515),
.B(n_1059),
.C(n_481),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_1048),
.B(n_1057),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1028),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1109),
.B(n_486),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_1109),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1028),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1109),
.B(n_486),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_1048),
.B(n_1057),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_966),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_1105),
.B(n_615),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1109),
.A2(n_464),
.B1(n_486),
.B2(n_747),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1109),
.A2(n_818),
.B1(n_515),
.B2(n_399),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1094),
.A2(n_1096),
.A3(n_1098),
.B(n_1091),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1058),
.A2(n_1051),
.B(n_973),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_986),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1109),
.A2(n_464),
.B1(n_486),
.B2(n_747),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1100),
.A2(n_515),
.B(n_1059),
.C(n_481),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1103),
.A2(n_1107),
.B(n_1104),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1200),
.A2(n_1246),
.B1(n_1225),
.B2(n_1165),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1121),
.Y(n_1254)
);

CKINVDCx6p67_ASAP7_75t_R g1255 ( 
.A(n_1123),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1171),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1201),
.A2(n_1219),
.B1(n_1250),
.B2(n_1243),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_1202),
.Y(n_1258)
);

INVx6_ASAP7_75t_L g1259 ( 
.A(n_1183),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1173),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1189),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1243),
.A2(n_1250),
.B1(n_1116),
.B2(n_1124),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1133),
.A2(n_1187),
.B1(n_1165),
.B2(n_1235),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1220),
.Y(n_1264)
);

BUFx12f_ASAP7_75t_L g1265 ( 
.A(n_1223),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1241),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1190),
.A2(n_1230),
.B1(n_1221),
.B2(n_1129),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1130),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1131),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1237),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1192),
.A2(n_1120),
.B1(n_1211),
.B2(n_1206),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1135),
.Y(n_1272)
);

INVx6_ASAP7_75t_SL g1273 ( 
.A(n_1204),
.Y(n_1273)
);

BUFx4f_ASAP7_75t_SL g1274 ( 
.A(n_1148),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1207),
.A2(n_1239),
.B(n_1141),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1224),
.B(n_1249),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1166),
.A2(n_1132),
.B1(n_1129),
.B2(n_1238),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1139),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1146),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1152),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1193),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1122),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1234),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1198),
.A2(n_1204),
.B1(n_1210),
.B2(n_1249),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1210),
.A2(n_1163),
.B1(n_1216),
.B2(n_1175),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1194),
.A2(n_1232),
.B1(n_1251),
.B2(n_1217),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1210),
.A2(n_1150),
.B1(n_1184),
.B2(n_1156),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1226),
.Y(n_1288)
);

AOI21xp33_ASAP7_75t_L g1289 ( 
.A1(n_1127),
.A2(n_1147),
.B(n_1209),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1115),
.A2(n_1144),
.B1(n_1242),
.B2(n_1175),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1155),
.Y(n_1291)
);

CKINVDCx11_ASAP7_75t_R g1292 ( 
.A(n_1237),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1126),
.A2(n_1231),
.B1(n_1181),
.B2(n_1157),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1162),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1158),
.A2(n_1143),
.B1(n_1151),
.B2(n_1160),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1162),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1174),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1113),
.Y(n_1298)
);

INVx6_ASAP7_75t_L g1299 ( 
.A(n_1113),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1118),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1151),
.A2(n_1142),
.B1(n_1149),
.B2(n_1182),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1159),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1159),
.Y(n_1303)
);

BUFx8_ASAP7_75t_L g1304 ( 
.A(n_1186),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1128),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1110),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1136),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1149),
.A2(n_1169),
.B1(n_1179),
.B2(n_1110),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1247),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1136),
.Y(n_1310)
);

AND2x2_ASAP7_75t_SL g1311 ( 
.A(n_1134),
.B(n_1111),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1134),
.A2(n_1127),
.B1(n_1179),
.B2(n_1172),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1178),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1195),
.A2(n_1215),
.B1(n_1154),
.B2(n_1164),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_SL g1315 ( 
.A(n_1195),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1170),
.A2(n_1215),
.B1(n_1154),
.B2(n_1197),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1136),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1128),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1168),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1128),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1113),
.A2(n_1138),
.B1(n_1240),
.B2(n_1233),
.Y(n_1321)
);

BUFx10_ASAP7_75t_L g1322 ( 
.A(n_1186),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1138),
.A2(n_1167),
.B1(n_1196),
.B2(n_1222),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1138),
.A2(n_1240),
.B1(n_1233),
.B2(n_1222),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1247),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1247),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1153),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1196),
.A2(n_1180),
.B1(n_1161),
.B2(n_1188),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1112),
.A2(n_1252),
.B1(n_1203),
.B2(n_1205),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1111),
.A2(n_1244),
.B1(n_1214),
.B2(n_1218),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1212),
.A2(n_1213),
.B1(n_1229),
.B2(n_1236),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1119),
.A2(n_1145),
.B1(n_1245),
.B2(n_1125),
.Y(n_1332)
);

INVx6_ASAP7_75t_L g1333 ( 
.A(n_1176),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1177),
.B(n_1114),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1111),
.A2(n_1137),
.B1(n_1114),
.B2(n_1248),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1191),
.A2(n_1208),
.B1(n_1228),
.B2(n_1227),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1185),
.Y(n_1337)
);

INVx3_ASAP7_75t_L g1338 ( 
.A(n_1114),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1199),
.A2(n_1200),
.B1(n_1246),
.B2(n_1225),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1140),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1183),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1200),
.A2(n_1246),
.B1(n_1225),
.B2(n_1211),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1200),
.A2(n_930),
.B1(n_912),
.B2(n_755),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1200),
.A2(n_930),
.B1(n_912),
.B2(n_755),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1121),
.Y(n_1345)
);

BUFx8_ASAP7_75t_L g1346 ( 
.A(n_1123),
.Y(n_1346)
);

BUFx2_ASAP7_75t_SL g1347 ( 
.A(n_1189),
.Y(n_1347)
);

CKINVDCx11_ASAP7_75t_R g1348 ( 
.A(n_1123),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1223),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1189),
.Y(n_1350)
);

BUFx12f_ASAP7_75t_L g1351 ( 
.A(n_1202),
.Y(n_1351)
);

INVx6_ASAP7_75t_L g1352 ( 
.A(n_1183),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1189),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1174),
.B(n_976),
.Y(n_1354)
);

INVx6_ASAP7_75t_L g1355 ( 
.A(n_1183),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1121),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1121),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1200),
.A2(n_1246),
.B1(n_1225),
.B2(n_1211),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1202),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1200),
.A2(n_1246),
.B1(n_1225),
.B2(n_1211),
.Y(n_1360)
);

INVx4_ASAP7_75t_L g1361 ( 
.A(n_1223),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1201),
.A2(n_755),
.B1(n_1219),
.B2(n_930),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1200),
.A2(n_1225),
.B1(n_1246),
.B2(n_1243),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1201),
.A2(n_755),
.B1(n_1219),
.B2(n_930),
.Y(n_1364)
);

BUFx12f_ASAP7_75t_L g1365 ( 
.A(n_1202),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1201),
.A2(n_755),
.B1(n_1219),
.B2(n_930),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1121),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1247),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1121),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1201),
.A2(n_755),
.B1(n_1219),
.B2(n_930),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1121),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1117),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1116),
.B(n_1224),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1121),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1200),
.A2(n_1225),
.B1(n_1246),
.B2(n_1243),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1202),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1200),
.A2(n_930),
.B1(n_912),
.B2(n_755),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1201),
.A2(n_755),
.B1(n_1219),
.B2(n_930),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1200),
.A2(n_930),
.B1(n_912),
.B2(n_755),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1254),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1331),
.A2(n_1332),
.B(n_1336),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1325),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1326),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1309),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1294),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1268),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1311),
.B(n_1309),
.Y(n_1387)
);

AOI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1339),
.A2(n_1286),
.B(n_1340),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1363),
.B(n_1375),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1296),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1368),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1329),
.A2(n_1338),
.B(n_1295),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1368),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1373),
.B(n_1275),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1259),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1334),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1329),
.A2(n_1338),
.B(n_1312),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1363),
.B(n_1375),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_SL g1399 ( 
.A1(n_1342),
.A2(n_1358),
.B(n_1360),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1311),
.Y(n_1400)
);

CKINVDCx16_ASAP7_75t_R g1401 ( 
.A(n_1260),
.Y(n_1401)
);

AOI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1327),
.A2(n_1314),
.B(n_1305),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1269),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1320),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1318),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1312),
.A2(n_1256),
.B(n_1323),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1345),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1356),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1256),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1267),
.A2(n_1330),
.B(n_1289),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1253),
.A2(n_1267),
.B(n_1262),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1343),
.A2(n_1379),
.B1(n_1344),
.B2(n_1377),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1357),
.Y(n_1413)
);

BUFx2_ASAP7_75t_SL g1414 ( 
.A(n_1315),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1253),
.A2(n_1271),
.B(n_1290),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1303),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1259),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1343),
.A2(n_1379),
.B1(n_1344),
.B2(n_1377),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1367),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1369),
.B(n_1371),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1374),
.B(n_1307),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1278),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1279),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1280),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1257),
.A2(n_1271),
.B1(n_1277),
.B2(n_1263),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1378),
.A2(n_1364),
.B1(n_1362),
.B2(n_1370),
.Y(n_1426)
);

AOI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1276),
.A2(n_1317),
.B(n_1310),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1259),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1302),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1290),
.A2(n_1319),
.B(n_1281),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1335),
.B(n_1277),
.Y(n_1431)
);

AOI222xp33_ASAP7_75t_L g1432 ( 
.A1(n_1257),
.A2(n_1378),
.B1(n_1364),
.B2(n_1366),
.C1(n_1370),
.C2(n_1362),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1328),
.A2(n_1301),
.B(n_1287),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1319),
.A2(n_1283),
.B(n_1291),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1335),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1372),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1330),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1297),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1313),
.Y(n_1439)
);

NAND3xp33_ASAP7_75t_L g1440 ( 
.A(n_1293),
.B(n_1284),
.C(n_1366),
.Y(n_1440)
);

CKINVDCx16_ASAP7_75t_R g1441 ( 
.A(n_1351),
.Y(n_1441)
);

AO21x2_ASAP7_75t_L g1442 ( 
.A1(n_1316),
.A2(n_1321),
.B(n_1285),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1297),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1354),
.A2(n_1308),
.B(n_1324),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1297),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1273),
.A2(n_1337),
.B(n_1285),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1333),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1333),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1333),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1299),
.A2(n_1322),
.B(n_1298),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1348),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1347),
.B(n_1261),
.Y(n_1452)
);

AO21x2_ASAP7_75t_L g1453 ( 
.A1(n_1299),
.A2(n_1304),
.B(n_1306),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1341),
.B(n_1352),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1304),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1270),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1341),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1352),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1352),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1355),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_1282),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1355),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1264),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1396),
.B(n_1353),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1396),
.B(n_1350),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1400),
.B(n_1292),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_SL g1467 ( 
.A1(n_1389),
.A2(n_1376),
.B(n_1258),
.C(n_1266),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1421),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1380),
.B(n_1272),
.Y(n_1469)
);

AOI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1394),
.A2(n_1415),
.B1(n_1411),
.B2(n_1435),
.C(n_1410),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1461),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1398),
.A2(n_1349),
.B(n_1361),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1386),
.B(n_1349),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1400),
.B(n_1288),
.Y(n_1474)
);

AND2x6_ASAP7_75t_L g1475 ( 
.A(n_1448),
.B(n_1274),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1381),
.A2(n_1300),
.B(n_1359),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1387),
.B(n_1255),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1381),
.A2(n_1274),
.B(n_1265),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1387),
.B(n_1365),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1405),
.B(n_1346),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1403),
.Y(n_1481)
);

A2O1A1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1425),
.A2(n_1346),
.B(n_1418),
.C(n_1412),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1420),
.B(n_1437),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1397),
.A2(n_1392),
.B(n_1406),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1420),
.B(n_1437),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1425),
.A2(n_1431),
.B(n_1433),
.C(n_1435),
.Y(n_1486)
);

AOI221xp5_ASAP7_75t_L g1487 ( 
.A1(n_1431),
.A2(n_1426),
.B1(n_1399),
.B2(n_1440),
.C(n_1405),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1433),
.A2(n_1446),
.B(n_1406),
.C(n_1444),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1407),
.B(n_1408),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1404),
.B(n_1413),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1407),
.B(n_1408),
.Y(n_1491)
);

O2A1O1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1399),
.A2(n_1463),
.B(n_1430),
.C(n_1449),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1460),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1419),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1422),
.B(n_1423),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1404),
.B(n_1434),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1463),
.A2(n_1430),
.B(n_1447),
.C(n_1449),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1446),
.B(n_1444),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_L g1499 ( 
.A(n_1384),
.B(n_1391),
.C(n_1393),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1424),
.Y(n_1500)
);

AO32x2_ASAP7_75t_L g1501 ( 
.A1(n_1395),
.A2(n_1417),
.A3(n_1428),
.B1(n_1427),
.B2(n_1434),
.Y(n_1501)
);

AO32x1_ASAP7_75t_L g1502 ( 
.A1(n_1384),
.A2(n_1391),
.A3(n_1393),
.B1(n_1382),
.B2(n_1383),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1388),
.A2(n_1402),
.B(n_1450),
.Y(n_1503)
);

NAND4xp25_ASAP7_75t_L g1504 ( 
.A(n_1432),
.B(n_1452),
.C(n_1455),
.D(n_1459),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1430),
.B(n_1438),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1430),
.A2(n_1382),
.B1(n_1383),
.B2(n_1429),
.C(n_1434),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1438),
.B(n_1443),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1443),
.B(n_1388),
.Y(n_1508)
);

NOR2x1_ASAP7_75t_R g1509 ( 
.A(n_1451),
.B(n_1461),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1452),
.Y(n_1510)
);

NOR2x1_ASAP7_75t_SL g1511 ( 
.A(n_1442),
.B(n_1453),
.Y(n_1511)
);

AO32x2_ASAP7_75t_L g1512 ( 
.A1(n_1402),
.A2(n_1436),
.A3(n_1390),
.B1(n_1385),
.B2(n_1416),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1481),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1505),
.B(n_1443),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1490),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1475),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1512),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1508),
.B(n_1468),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1512),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1470),
.A2(n_1442),
.B1(n_1458),
.B2(n_1457),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1489),
.B(n_1409),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1507),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1512),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1508),
.B(n_1445),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1512),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1490),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1489),
.B(n_1491),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1487),
.A2(n_1504),
.B1(n_1506),
.B2(n_1442),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1480),
.B(n_1462),
.Y(n_1529)
);

NAND2x1p5_ASAP7_75t_SL g1530 ( 
.A(n_1466),
.B(n_1454),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1483),
.B(n_1485),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1466),
.A2(n_1442),
.B1(n_1457),
.B2(n_1401),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1499),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1512),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1494),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1500),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1496),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1495),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1528),
.A2(n_1486),
.B1(n_1482),
.B2(n_1480),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1517),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1531),
.B(n_1510),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1533),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_1533),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1517),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1517),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1535),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1528),
.A2(n_1520),
.B1(n_1532),
.B2(n_1517),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1535),
.B(n_1495),
.Y(n_1548)
);

INVxp67_ASAP7_75t_SL g1549 ( 
.A(n_1519),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1518),
.B(n_1464),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1518),
.B(n_1465),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1531),
.B(n_1476),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1516),
.Y(n_1553)
);

INVx5_ASAP7_75t_L g1554 ( 
.A(n_1516),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1529),
.Y(n_1555)
);

OAI31xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1529),
.A2(n_1472),
.A3(n_1479),
.B(n_1477),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_L g1557 ( 
.A1(n_1520),
.A2(n_1492),
.B(n_1488),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1530),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1513),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1514),
.B(n_1476),
.Y(n_1560)
);

AO21x2_ASAP7_75t_L g1561 ( 
.A1(n_1519),
.A2(n_1503),
.B(n_1497),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1513),
.Y(n_1562)
);

OAI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1532),
.A2(n_1498),
.B1(n_1523),
.B2(n_1534),
.C(n_1519),
.Y(n_1563)
);

NAND3xp33_ASAP7_75t_L g1564 ( 
.A(n_1523),
.B(n_1476),
.C(n_1478),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1514),
.B(n_1501),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1523),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1523),
.A2(n_1474),
.B1(n_1498),
.B2(n_1484),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1537),
.A2(n_1502),
.B(n_1511),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_SL g1569 ( 
.A1(n_1516),
.A2(n_1478),
.B(n_1511),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1531),
.B(n_1493),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1515),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1525),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1515),
.A2(n_1473),
.B1(n_1469),
.B2(n_1477),
.C(n_1479),
.Y(n_1573)
);

NAND3xp33_ASAP7_75t_L g1574 ( 
.A(n_1525),
.B(n_1478),
.C(n_1467),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1543),
.B(n_1542),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1542),
.B(n_1525),
.C(n_1534),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1543),
.B(n_1526),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1559),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1558),
.B(n_1526),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1541),
.B(n_1548),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1540),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1541),
.B(n_1527),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1571),
.B(n_1536),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1540),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_SL g1585 ( 
.A(n_1555),
.B(n_1471),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1559),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1571),
.B(n_1536),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1541),
.B(n_1527),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1565),
.B(n_1524),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1565),
.B(n_1524),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1546),
.B(n_1536),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1548),
.B(n_1521),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1555),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1550),
.B(n_1522),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1553),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1554),
.B(n_1516),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1554),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1553),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1570),
.B(n_1521),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1565),
.B(n_1538),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1559),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1546),
.B(n_1573),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1570),
.B(n_1441),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1562),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1546),
.B(n_1525),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1573),
.B(n_1534),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1578),
.Y(n_1607)
);

OR2x2_ASAP7_75t_SL g1608 ( 
.A(n_1575),
.B(n_1401),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1581),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1578),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1603),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1575),
.B(n_1556),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1581),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1583),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1606),
.A2(n_1556),
.B(n_1557),
.Y(n_1615)
);

AND2x4_ASAP7_75t_SL g1616 ( 
.A(n_1596),
.B(n_1456),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1583),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1587),
.Y(n_1618)
);

INVx2_ASAP7_75t_SL g1619 ( 
.A(n_1595),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1581),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1587),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1580),
.B(n_1570),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1595),
.B(n_1551),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1595),
.B(n_1551),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1580),
.B(n_1552),
.Y(n_1625)
);

OR2x6_ASAP7_75t_L g1626 ( 
.A(n_1597),
.B(n_1569),
.Y(n_1626)
);

OAI21xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1602),
.A2(n_1544),
.B(n_1549),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1602),
.B(n_1561),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1598),
.B(n_1553),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1582),
.B(n_1547),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1598),
.B(n_1551),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1586),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1596),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1586),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1593),
.B(n_1561),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1593),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1582),
.B(n_1588),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1606),
.B(n_1552),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1601),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1577),
.B(n_1561),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1589),
.B(n_1551),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1601),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1604),
.Y(n_1643)
);

AND2x4_ASAP7_75t_SL g1644 ( 
.A(n_1596),
.B(n_1456),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1584),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1599),
.B(n_1552),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1599),
.B(n_1540),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1604),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1615),
.B(n_1576),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1636),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1632),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1609),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1634),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1616),
.B(n_1589),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1616),
.B(n_1589),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1644),
.B(n_1590),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1614),
.B(n_1577),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1617),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1618),
.B(n_1576),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1621),
.B(n_1600),
.Y(n_1660)
);

AND2x2_ASAP7_75t_SL g1661 ( 
.A(n_1612),
.B(n_1547),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1609),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1639),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1644),
.B(n_1590),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1623),
.B(n_1590),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1637),
.B(n_1600),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1607),
.B(n_1600),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1642),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1629),
.B(n_1585),
.Y(n_1669)
);

NAND2x1_ASAP7_75t_L g1670 ( 
.A(n_1626),
.B(n_1579),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1622),
.B(n_1592),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1629),
.B(n_1574),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1629),
.B(n_1574),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1623),
.B(n_1594),
.Y(n_1674)
);

OAI31xp33_ASAP7_75t_L g1675 ( 
.A1(n_1630),
.A2(n_1557),
.A3(n_1539),
.B(n_1563),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1619),
.B(n_1579),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1610),
.B(n_1591),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1643),
.Y(n_1678)
);

OAI322xp33_ASAP7_75t_L g1679 ( 
.A1(n_1628),
.A2(n_1539),
.A3(n_1605),
.B1(n_1568),
.B2(n_1549),
.C1(n_1544),
.C2(n_1563),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1648),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1638),
.B(n_1592),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1624),
.B(n_1641),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1613),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1651),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1649),
.A2(n_1608),
.B1(n_1611),
.B2(n_1574),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1650),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1649),
.A2(n_1627),
.B(n_1635),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1650),
.B(n_1619),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1676),
.Y(n_1689)
);

NAND4xp25_ASAP7_75t_L g1690 ( 
.A(n_1672),
.B(n_1633),
.C(n_1624),
.D(n_1638),
.Y(n_1690)
);

INVxp67_ASAP7_75t_SL g1691 ( 
.A(n_1670),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1651),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1661),
.A2(n_1557),
.B(n_1640),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1679),
.A2(n_1564),
.B1(n_1568),
.B2(n_1572),
.C(n_1540),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1682),
.B(n_1631),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1682),
.Y(n_1696)
);

OAI211xp5_ASAP7_75t_L g1697 ( 
.A1(n_1673),
.A2(n_1633),
.B(n_1631),
.C(n_1597),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1661),
.A2(n_1564),
.B(n_1626),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1653),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1661),
.B(n_1456),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1653),
.Y(n_1701)
);

INVxp67_ASAP7_75t_SL g1702 ( 
.A(n_1670),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1675),
.A2(n_1564),
.B1(n_1567),
.B2(n_1626),
.C(n_1534),
.Y(n_1703)
);

A2O1A1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1675),
.A2(n_1567),
.B(n_1560),
.C(n_1625),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1679),
.B(n_1441),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1663),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1671),
.B(n_1456),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1669),
.B(n_1456),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1686),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1696),
.B(n_1671),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1689),
.B(n_1665),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1684),
.Y(n_1713)
);

OAI32xp33_ASAP7_75t_L g1714 ( 
.A1(n_1705),
.A2(n_1659),
.A3(n_1681),
.B1(n_1657),
.B2(n_1667),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1692),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1695),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1700),
.B(n_1688),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1700),
.B(n_1665),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1705),
.A2(n_1561),
.B1(n_1659),
.B2(n_1683),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1708),
.B(n_1674),
.Y(n_1720)
);

INVxp33_ASAP7_75t_L g1721 ( 
.A(n_1707),
.Y(n_1721)
);

INVxp67_ASAP7_75t_SL g1722 ( 
.A(n_1691),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1704),
.A2(n_1666),
.B1(n_1626),
.B2(n_1681),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1707),
.B(n_1674),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_SL g1725 ( 
.A1(n_1698),
.A2(n_1703),
.B1(n_1693),
.B2(n_1685),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1699),
.Y(n_1726)
);

AOI322xp5_ASAP7_75t_L g1727 ( 
.A1(n_1704),
.A2(n_1666),
.A3(n_1660),
.B1(n_1683),
.B2(n_1652),
.C1(n_1662),
.C2(n_1667),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1711),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1709),
.Y(n_1729)
);

XOR2x2_ASAP7_75t_L g1730 ( 
.A(n_1723),
.B(n_1687),
.Y(n_1730)
);

AOI21xp33_ASAP7_75t_L g1731 ( 
.A1(n_1714),
.A2(n_1702),
.B(n_1701),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1725),
.A2(n_1690),
.B1(n_1694),
.B2(n_1652),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1724),
.B(n_1716),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1727),
.A2(n_1697),
.B(n_1706),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1716),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1710),
.Y(n_1736)
);

NOR2xp67_ASAP7_75t_L g1737 ( 
.A(n_1712),
.B(n_1633),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1722),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1719),
.A2(n_1668),
.B(n_1663),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1733),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1732),
.A2(n_1717),
.B(n_1721),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1733),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1738),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1735),
.Y(n_1744)
);

NOR3xp33_ASAP7_75t_SL g1745 ( 
.A(n_1734),
.B(n_1717),
.C(n_1715),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1728),
.B(n_1721),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1729),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1732),
.A2(n_1720),
.B(n_1718),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1736),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1745),
.A2(n_1739),
.B1(n_1731),
.B2(n_1726),
.C(n_1713),
.Y(n_1750)
);

O2A1O1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1745),
.A2(n_1730),
.B(n_1737),
.C(n_1720),
.Y(n_1751)
);

NAND4xp25_ASAP7_75t_L g1752 ( 
.A(n_1748),
.B(n_1730),
.C(n_1654),
.D(n_1664),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1741),
.A2(n_1683),
.B1(n_1652),
.B2(n_1662),
.Y(n_1753)
);

AOI22x1_ASAP7_75t_L g1754 ( 
.A1(n_1740),
.A2(n_1456),
.B1(n_1678),
.B2(n_1668),
.Y(n_1754)
);

OAI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1753),
.A2(n_1746),
.B1(n_1742),
.B2(n_1744),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_L g1756 ( 
.A(n_1750),
.B(n_1749),
.C(n_1743),
.Y(n_1756)
);

OAI211xp5_ASAP7_75t_L g1757 ( 
.A1(n_1751),
.A2(n_1749),
.B(n_1747),
.C(n_1680),
.Y(n_1757)
);

AOI32xp33_ASAP7_75t_L g1758 ( 
.A1(n_1752),
.A2(n_1680),
.A3(n_1678),
.B1(n_1654),
.B2(n_1664),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1754),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1750),
.A2(n_1662),
.B1(n_1656),
.B2(n_1655),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1757),
.Y(n_1761)
);

NOR2x1_ASAP7_75t_L g1762 ( 
.A(n_1755),
.B(n_1677),
.Y(n_1762)
);

NOR3xp33_ASAP7_75t_L g1763 ( 
.A(n_1756),
.B(n_1509),
.C(n_1439),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1759),
.B(n_1655),
.Y(n_1764)
);

NOR2x1_ASAP7_75t_L g1765 ( 
.A(n_1758),
.B(n_1677),
.Y(n_1765)
);

NOR3xp33_ASAP7_75t_L g1766 ( 
.A(n_1761),
.B(n_1760),
.C(n_1613),
.Y(n_1766)
);

A2O1A1Ixp33_ASAP7_75t_SL g1767 ( 
.A1(n_1763),
.A2(n_1660),
.B(n_1656),
.C(n_1645),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1764),
.B(n_1579),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1768),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1769),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1766),
.B1(n_1762),
.B2(n_1765),
.Y(n_1771)
);

XNOR2xp5_ASAP7_75t_L g1772 ( 
.A(n_1770),
.B(n_1767),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1772),
.Y(n_1773)
);

OAI22x1_ASAP7_75t_SL g1774 ( 
.A1(n_1771),
.A2(n_1471),
.B1(n_1455),
.B2(n_1645),
.Y(n_1774)
);

AOI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1773),
.A2(n_1620),
.B1(n_1572),
.B2(n_1545),
.C(n_1566),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1774),
.Y(n_1776)
);

AOI21xp33_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1620),
.B(n_1625),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1777),
.A2(n_1775),
.B(n_1646),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1778),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1414),
.B1(n_1605),
.B2(n_1584),
.C(n_1646),
.Y(n_1780)
);

AOI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1780),
.A2(n_1454),
.B(n_1647),
.C(n_1414),
.Y(n_1781)
);


endmodule