module fake_netlist_1_1947_n_1809 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_407, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_383, n_6, n_400, n_296, n_157, n_79, n_202, n_386, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_389, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_387, n_163, n_105, n_227, n_384, n_231, n_298, n_411, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_401, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_392, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_393, n_24, n_247, n_381, n_304, n_399, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_402, n_32, n_413, n_391, n_235, n_243, n_415, n_394, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_404, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_412, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_403, n_254, n_262, n_10, n_239, n_87, n_379, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_388, n_193, n_273, n_390, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_416, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_409, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_396, n_168, n_398, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_397, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_410, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_380, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_382, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_332, n_414, n_350, n_164, n_175, n_145, n_408, n_290, n_405, n_280, n_21, n_99, n_109, n_132, n_395, n_406, n_151, n_385, n_257, n_269, n_1809);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_407;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_383;
input n_6;
input n_400;
input n_296;
input n_157;
input n_79;
input n_202;
input n_386;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_389;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_387;
input n_163;
input n_105;
input n_227;
input n_384;
input n_231;
input n_298;
input n_411;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_401;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_392;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_393;
input n_24;
input n_247;
input n_381;
input n_304;
input n_399;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_402;
input n_32;
input n_413;
input n_391;
input n_235;
input n_243;
input n_415;
input n_394;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_404;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_412;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_403;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_379;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_388;
input n_193;
input n_273;
input n_390;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_416;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_409;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_396;
input n_168;
input n_398;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_397;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_410;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_380;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_382;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_414;
input n_350;
input n_164;
input n_175;
input n_145;
input n_408;
input n_290;
input n_405;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_395;
input n_406;
input n_151;
input n_385;
input n_257;
input n_269;
output n_1809;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_1671;
wire n_646;
wire n_1334;
wire n_1627;
wire n_1698;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_1785;
wire n_965;
wire n_1646;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_1667;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_1782;
wire n_877;
wire n_1663;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1743;
wire n_1019;
wire n_1714;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_452;
wire n_518;
wire n_1336;
wire n_1341;
wire n_1381;
wire n_1760;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1672;
wire n_1342;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_1631;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_1661;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1683;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_533;
wire n_1010;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_1656;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_1744;
wire n_501;
wire n_699;
wire n_1654;
wire n_551;
wire n_1061;
wire n_509;
wire n_849;
wire n_1732;
wire n_864;
wire n_1772;
wire n_961;
wire n_1525;
wire n_1718;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1739;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1775;
wire n_1620;
wire n_537;
wire n_1764;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1758;
wire n_1406;
wire n_1789;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_1623;
wire n_556;
wire n_1214;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_1707;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_1731;
wire n_514;
wire n_1693;
wire n_1690;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1790;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1703;
wire n_1377;
wire n_1079;
wire n_1582;
wire n_1321;
wire n_1801;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1728;
wire n_1385;
wire n_1711;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_1716;
wire n_1662;
wire n_790;
wire n_761;
wire n_1660;
wire n_1287;
wire n_472;
wire n_1100;
wire n_1648;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_1695;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1788;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1682;
wire n_1740;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_1639;
wire n_1730;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_1768;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1802;
wire n_1164;
wire n_1628;
wire n_1533;
wire n_1611;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1694;
wire n_1563;
wire n_1642;
wire n_824;
wire n_793;
wire n_1792;
wire n_753;
wire n_1753;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_992;
wire n_1748;
wire n_1754;
wire n_1077;
wire n_838;
wire n_705;
wire n_1741;
wire n_964;
wire n_590;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1681;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1602;
wire n_1769;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_1733;
wire n_911;
wire n_980;
wire n_1675;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1709;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1625;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_1725;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_1787;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_1629;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1670;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1807;
wire n_1791;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_1643;
wire n_1687;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_550;
wire n_826;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1537;
wire n_634;
wire n_1271;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_478;
wire n_482;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1777;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1778;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_1710;
wire n_1781;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1765;
wire n_1050;
wire n_1593;
wire n_1763;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_1647;
wire n_1621;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1668;
wire n_1692;
wire n_1153;
wire n_1797;
wire n_1657;
wire n_1655;
wire n_1771;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_1762;
wire n_942;
wire n_1029;
wire n_1665;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1766;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1696;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_1796;
wire n_734;
wire n_919;
wire n_763;
wire n_1724;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_1638;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1752;
wire n_1645;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_1633;
wire n_1784;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1626;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_1800;
wire n_515;
wire n_1577;
wire n_1719;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1641;
wire n_1798;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_1705;
wire n_457;
wire n_1799;
wire n_1757;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1729;
wire n_1585;
wire n_1425;
wire n_1292;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_1697;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_1720;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1679;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_1688;
wire n_1767;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_1634;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_1455;
wire n_659;
wire n_432;
wire n_1329;
wire n_1750;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_436;
wire n_1653;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1640;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1658;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_1761;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_1795;
wire n_1659;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1734;
wire n_1701;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_1272;
wire n_928;
wire n_882;
wire n_1635;
wire n_871;
wire n_803;
wire n_1704;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1759;
wire n_1774;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_516;
wire n_549;
wire n_1576;
wire n_1609;
wire n_832;
wire n_996;
wire n_1578;
wire n_1794;
wire n_420;
wire n_1684;
wire n_1089;
wire n_1717;
wire n_1434;
wire n_1058;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_1706;
wire n_1473;
wire n_1678;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1674;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1622;
wire n_1755;
wire n_1804;
wire n_1773;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1712;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1779;
wire n_1170;
wire n_1523;
wire n_1700;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1636;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1722;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_1726;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1735;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1689;
wire n_1756;
wire n_1805;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_1624;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_1699;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_1713;
wire n_913;
wire n_845;
wire n_1776;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_1780;
wire n_934;
wire n_425;
wire n_1737;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1749;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_1786;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_1806;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_1676;
wire n_678;
wire n_1200;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_1708;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_1666;
wire n_1169;
wire n_975;
wire n_1721;
wire n_1081;
wire n_1680;
wire n_1644;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_1669;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1673;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1742;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1736;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_1630;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1808;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1793;
wire n_1041;
wire n_1745;
wire n_1080;
wire n_1727;
wire n_1637;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1632;
wire n_1738;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_1664;
wire n_682;
wire n_1607;
wire n_906;
wire n_1650;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1702;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1685;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1335;
wire n_1239;
wire n_924;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1677;
wire n_1296;
wire n_1751;
wire n_1428;
wire n_766;
wire n_602;
wire n_1649;
wire n_1143;
wire n_629;
wire n_1723;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1783;
wire n_1390;
wire n_1691;
wire n_1715;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_1747;
wire n_418;
wire n_1686;
wire n_600;
wire n_1531;
wire n_1548;
wire n_1651;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_1770;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_1652;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_1803;
wire n_1398;
wire n_491;
wire n_1746;
wire n_1291;
INVx1_ASAP7_75t_L g417 ( .A(n_68), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_272), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_295), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_68), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_70), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_121), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_328), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_118), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_298), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_258), .Y(n_426) );
XNOR2x1_ASAP7_75t_L g427 ( .A(n_287), .B(n_184), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_86), .Y(n_428) );
INVxp33_ASAP7_75t_L g429 ( .A(n_58), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_139), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_383), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_412), .Y(n_432) );
INVx1_ASAP7_75t_SL g433 ( .A(n_41), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_90), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_278), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_360), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_100), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_326), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_372), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_189), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_172), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_183), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_376), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_39), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_27), .Y(n_445) );
INVxp33_ASAP7_75t_L g446 ( .A(n_270), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_155), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_345), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_315), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_361), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_358), .Y(n_451) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_367), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_329), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_143), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_282), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_364), .Y(n_456) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_279), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_1), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_408), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_192), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_133), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_120), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_181), .B(n_53), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_373), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_164), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_108), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_144), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_220), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_55), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_378), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_99), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_236), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_232), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_151), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_9), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_406), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_355), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_352), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_255), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_238), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_75), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_407), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_362), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_179), .Y(n_484) );
INVxp67_ASAP7_75t_L g485 ( .A(n_413), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_229), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_370), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_400), .B(n_70), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_45), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_350), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_349), .B(n_381), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_108), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_40), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_296), .B(n_174), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_114), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_318), .Y(n_496) );
BUFx5_ASAP7_75t_L g497 ( .A(n_226), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_347), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_103), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_216), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_18), .Y(n_501) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_233), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_75), .Y(n_503) );
CKINVDCx14_ASAP7_75t_R g504 ( .A(n_176), .Y(n_504) );
INVxp33_ASAP7_75t_L g505 ( .A(n_416), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_203), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_163), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_14), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_401), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_132), .Y(n_510) );
NOR2xp67_ASAP7_75t_L g511 ( .A(n_138), .B(n_180), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_260), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_377), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_250), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_185), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_81), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_147), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_379), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_193), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_266), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_121), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_330), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_346), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_139), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_154), .Y(n_525) );
NOR2xp67_ASAP7_75t_L g526 ( .A(n_19), .B(n_223), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_210), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_262), .Y(n_528) );
BUFx2_ASAP7_75t_L g529 ( .A(n_304), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_138), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_291), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_399), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_392), .Y(n_533) );
CKINVDCx14_ASAP7_75t_R g534 ( .A(n_132), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_249), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_175), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_134), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_197), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_199), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_375), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_227), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_101), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_88), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_277), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_222), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_252), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_177), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_152), .Y(n_548) );
INVxp67_ASAP7_75t_L g549 ( .A(n_32), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_363), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_60), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_297), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_331), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_23), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_90), .B(n_237), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_110), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_267), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_327), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_28), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_5), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_137), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_273), .Y(n_562) );
NOR2xp67_ASAP7_75t_L g563 ( .A(n_71), .B(n_385), .Y(n_563) );
INVxp67_ASAP7_75t_SL g564 ( .A(n_72), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_72), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_411), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_202), .Y(n_567) );
BUFx8_ASAP7_75t_SL g568 ( .A(n_308), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_3), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_112), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_382), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_81), .Y(n_572) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_322), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_170), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_182), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_388), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_224), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_312), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_305), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_234), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_112), .Y(n_581) );
INVxp33_ASAP7_75t_SL g582 ( .A(n_374), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_64), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_317), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_228), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_274), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_285), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_194), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_169), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_115), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_245), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_4), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_371), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_254), .Y(n_594) );
BUFx10_ASAP7_75t_L g595 ( .A(n_141), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_167), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_88), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_195), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_235), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_332), .Y(n_600) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_178), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g602 ( .A(n_196), .B(n_61), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_414), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_264), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_248), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_256), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_92), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_230), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_86), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_316), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_303), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_42), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_149), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_288), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_40), .Y(n_615) );
BUFx10_ASAP7_75t_L g616 ( .A(n_294), .Y(n_616) );
BUFx10_ASAP7_75t_L g617 ( .A(n_158), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_300), .Y(n_618) );
CKINVDCx14_ASAP7_75t_R g619 ( .A(n_191), .Y(n_619) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_134), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_309), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_359), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_231), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_221), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_84), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_103), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_356), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_53), .Y(n_628) );
BUFx8_ASAP7_75t_SL g629 ( .A(n_42), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_208), .Y(n_630) );
INVx3_ASAP7_75t_L g631 ( .A(n_289), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_499), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_631), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_499), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_429), .B(n_0), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_542), .Y(n_636) );
BUFx2_ASAP7_75t_L g637 ( .A(n_534), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_568), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_542), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_418), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_631), .B(n_0), .Y(n_641) );
OA21x2_ASAP7_75t_L g642 ( .A1(n_460), .A2(n_142), .B(n_140), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_419), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_497), .Y(n_644) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_450), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_497), .Y(n_646) );
OAI22xp5_ASAP7_75t_SL g647 ( .A1(n_462), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_423), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_495), .Y(n_649) );
INVx3_ASAP7_75t_L g650 ( .A(n_595), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_497), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_534), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_432), .Y(n_653) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_450), .Y(n_654) );
INVx5_ASAP7_75t_L g655 ( .A(n_450), .Y(n_655) );
INVx3_ASAP7_75t_L g656 ( .A(n_595), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_495), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_429), .A2(n_5), .B1(n_2), .B2(n_4), .Y(n_658) );
INVx3_ASAP7_75t_L g659 ( .A(n_616), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_564), .A2(n_8), .B1(n_6), .B2(n_7), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_497), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_436), .B(n_6), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_435), .Y(n_663) );
INVx6_ASAP7_75t_L g664 ( .A(n_616), .Y(n_664) );
OA21x2_ASAP7_75t_L g665 ( .A1(n_460), .A2(n_146), .B(n_145), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_439), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_497), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_568), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_448), .B(n_7), .Y(n_669) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_450), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_440), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_650), .B(n_446), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_645), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_644), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_644), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_644), .Y(n_676) );
BUFx3_ASAP7_75t_L g677 ( .A(n_642), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_646), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_640), .B(n_532), .Y(n_679) );
INVx4_ASAP7_75t_L g680 ( .A(n_642), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_646), .Y(n_681) );
INVx2_ASAP7_75t_SL g682 ( .A(n_633), .Y(n_682) );
BUFx3_ASAP7_75t_L g683 ( .A(n_642), .Y(n_683) );
INVx3_ASAP7_75t_L g684 ( .A(n_646), .Y(n_684) );
BUFx3_ASAP7_75t_L g685 ( .A(n_642), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_650), .B(n_446), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_651), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_640), .B(n_571), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_645), .Y(n_689) );
INVx3_ASAP7_75t_L g690 ( .A(n_651), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_643), .A2(n_420), .B1(n_444), .B2(n_417), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_645), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_658), .B(n_564), .C(n_560), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_645), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_645), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_643), .B(n_447), .C(n_442), .Y(n_696) );
INVx2_ASAP7_75t_SL g697 ( .A(n_633), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_645), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_648), .A2(n_458), .B1(n_466), .B2(n_445), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_637), .Y(n_700) );
AO22x2_ASAP7_75t_L g701 ( .A1(n_635), .A2(n_427), .B1(n_502), .B2(n_457), .Y(n_701) );
INVx4_ASAP7_75t_L g702 ( .A(n_665), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_660), .A2(n_524), .B1(n_441), .B2(n_451), .Y(n_703) );
INVx3_ASAP7_75t_L g704 ( .A(n_651), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_661), .Y(n_705) );
NAND2xp33_ASAP7_75t_L g706 ( .A(n_648), .B(n_497), .Y(n_706) );
BUFx3_ASAP7_75t_L g707 ( .A(n_665), .Y(n_707) );
OR2x6_ASAP7_75t_L g708 ( .A(n_647), .B(n_529), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_682), .Y(n_709) );
BUFx2_ASAP7_75t_L g710 ( .A(n_700), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_682), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_697), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_693), .A2(n_641), .B(n_634), .C(n_636), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_697), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_697), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_672), .B(n_637), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_672), .B(n_652), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_686), .B(n_652), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_686), .B(n_649), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_688), .B(n_650), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_677), .A2(n_665), .B(n_661), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_688), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_693), .A2(n_653), .B1(n_666), .B2(n_663), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_680), .A2(n_653), .B1(n_666), .B2(n_663), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_700), .B(n_650), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_679), .B(n_656), .Y(n_726) );
NAND2xp33_ASAP7_75t_L g727 ( .A(n_674), .B(n_635), .Y(n_727) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_708), .A2(n_647), .B1(n_660), .B2(n_638), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g729 ( .A(n_703), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_679), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_677), .A2(n_665), .B(n_667), .Y(n_731) );
INVx2_ASAP7_75t_SL g732 ( .A(n_701), .Y(n_732) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_677), .Y(n_733) );
NOR3x1_ASAP7_75t_L g734 ( .A(n_703), .B(n_502), .C(n_457), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_680), .A2(n_671), .B1(n_667), .B2(n_634), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_674), .B(n_656), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_675), .B(n_656), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_696), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_675), .B(n_656), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_676), .B(n_671), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_684), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_701), .A2(n_453), .B1(n_515), .B2(n_438), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_676), .B(n_659), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_678), .B(n_659), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_680), .A2(n_636), .B1(n_639), .B2(n_632), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_678), .B(n_659), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_681), .B(n_659), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_691), .B(n_669), .C(n_662), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_701), .B(n_657), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_684), .Y(n_750) );
INVx4_ASAP7_75t_L g751 ( .A(n_684), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_681), .B(n_664), .Y(n_752) );
INVx2_ASAP7_75t_SL g753 ( .A(n_701), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_687), .B(n_443), .Y(n_754) );
BUFx3_ASAP7_75t_L g755 ( .A(n_684), .Y(n_755) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_683), .Y(n_756) );
A2O1A1Ixp33_ASAP7_75t_L g757 ( .A1(n_687), .A2(n_505), .B(n_639), .C(n_632), .Y(n_757) );
INVx3_ASAP7_75t_L g758 ( .A(n_690), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_683), .A2(n_491), .B(n_505), .Y(n_759) );
AND2x6_ASAP7_75t_SL g760 ( .A(n_708), .B(n_471), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_680), .A2(n_475), .B1(n_501), .B2(n_492), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_702), .B(n_664), .Y(n_762) );
O2A1O1Ixp33_ASAP7_75t_L g763 ( .A1(n_691), .A2(n_560), .B(n_549), .C(n_508), .Y(n_763) );
AND2x2_ASAP7_75t_SL g764 ( .A(n_706), .B(n_452), .Y(n_764) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_683), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_699), .B(n_664), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_685), .A2(n_538), .B(n_532), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_702), .B(n_479), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_699), .B(n_664), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_690), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_702), .B(n_514), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_705), .B(n_546), .Y(n_772) );
NOR3xp33_ASAP7_75t_L g773 ( .A(n_701), .B(n_668), .C(n_549), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_690), .Y(n_774) );
INVxp67_ASAP7_75t_L g775 ( .A(n_708), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_705), .B(n_504), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_702), .B(n_582), .Y(n_777) );
BUFx6f_ASAP7_75t_L g778 ( .A(n_685), .Y(n_778) );
NAND2xp5_ASAP7_75t_SL g779 ( .A(n_690), .B(n_455), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_708), .A2(n_528), .B1(n_588), .B2(n_527), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_704), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_704), .B(n_504), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_704), .B(n_619), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_685), .B(n_621), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_721), .A2(n_707), .B(n_704), .Y(n_785) );
O2A1O1Ixp5_ASAP7_75t_L g786 ( .A1(n_768), .A2(n_463), .B(n_480), .C(n_425), .Y(n_786) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_749), .A2(n_503), .B1(n_543), .B2(n_530), .C(n_521), .Y(n_787) );
AOI21x1_ASAP7_75t_L g788 ( .A1(n_731), .A2(n_759), .B(n_768), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_736), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_737), .Y(n_790) );
OAI21x1_ASAP7_75t_L g791 ( .A1(n_767), .A2(n_689), .B(n_673), .Y(n_791) );
O2A1O1Ixp33_ASAP7_75t_L g792 ( .A1(n_713), .A2(n_708), .B(n_556), .C(n_565), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_733), .A2(n_707), .B(n_494), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_733), .A2(n_707), .B(n_459), .Y(n_794) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_710), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g796 ( .A1(n_771), .A2(n_464), .B(n_456), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_760), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_719), .B(n_708), .Y(n_798) );
INVx3_ASAP7_75t_L g799 ( .A(n_751), .Y(n_799) );
AOI21x1_ASAP7_75t_L g800 ( .A1(n_771), .A2(n_689), .B(n_673), .Y(n_800) );
BUFx2_ASAP7_75t_L g801 ( .A(n_784), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_724), .A2(n_485), .B(n_468), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_739), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_777), .A2(n_472), .B(n_465), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_722), .B(n_433), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_751), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_777), .A2(n_762), .B(n_776), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g808 ( .A1(n_762), .A2(n_474), .B(n_473), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_725), .B(n_629), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_723), .B(n_421), .Y(n_810) );
NAND2xp5_ASAP7_75t_SL g811 ( .A(n_756), .B(n_426), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_775), .B(n_629), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_723), .B(n_422), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_772), .B(n_424), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_758), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_720), .B(n_428), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g817 ( .A(n_773), .B(n_761), .C(n_724), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_780), .B(n_784), .Y(n_818) );
INVxp67_ASAP7_75t_L g819 ( .A(n_754), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_716), .B(n_434), .Y(n_820) );
NAND2x1p5_ASAP7_75t_L g821 ( .A(n_756), .B(n_488), .Y(n_821) );
AO21x1_ASAP7_75t_L g822 ( .A1(n_782), .A2(n_483), .B(n_476), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_717), .B(n_437), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_758), .Y(n_824) );
OAI22x1_ASAP7_75t_L g825 ( .A1(n_729), .A2(n_481), .B1(n_489), .B2(n_469), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_742), .B(n_461), .Y(n_826) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_755), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_732), .A2(n_624), .B1(n_493), .B2(n_537), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_718), .B(n_510), .Y(n_829) );
BUFx2_ASAP7_75t_L g830 ( .A(n_753), .Y(n_830) );
NAND3xp33_ASAP7_75t_SL g831 ( .A(n_763), .B(n_516), .C(n_559), .Y(n_831) );
NOR2xp33_ASAP7_75t_R g832 ( .A(n_764), .B(n_619), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_783), .A2(n_487), .B(n_484), .Y(n_833) );
O2A1O1Ixp33_ASAP7_75t_L g834 ( .A1(n_713), .A2(n_569), .B(n_583), .C(n_551), .Y(n_834) );
AND2x4_ASAP7_75t_L g835 ( .A(n_748), .B(n_592), .Y(n_835) );
O2A1O1Ixp33_ASAP7_75t_L g836 ( .A1(n_757), .A2(n_612), .B(n_615), .C(n_609), .Y(n_836) );
NAND2xp5_ASAP7_75t_SL g837 ( .A(n_765), .B(n_449), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_727), .B(n_561), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_715), .A2(n_498), .B(n_490), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_766), .B(n_570), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_764), .A2(n_572), .B1(n_590), .B2(n_581), .Y(n_841) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_765), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_769), .B(n_597), .Y(n_843) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_743), .A2(n_512), .B(n_500), .Y(n_844) );
AOI21xp5_ASAP7_75t_L g845 ( .A1(n_744), .A2(n_517), .B(n_513), .Y(n_845) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_746), .A2(n_519), .B(n_518), .Y(n_846) );
BUFx3_ASAP7_75t_L g847 ( .A(n_750), .Y(n_847) );
O2A1O1Ixp33_ASAP7_75t_L g848 ( .A1(n_754), .A2(n_626), .B(n_628), .C(n_625), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_770), .Y(n_849) );
OAI21xp5_ASAP7_75t_L g850 ( .A1(n_735), .A2(n_485), .B(n_522), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_761), .B(n_620), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_741), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_747), .A2(n_539), .B(n_536), .Y(n_853) );
AO21x1_ASAP7_75t_L g854 ( .A1(n_779), .A2(n_541), .B(n_540), .Y(n_854) );
O2A1O1Ixp33_ASAP7_75t_SL g855 ( .A1(n_738), .A2(n_547), .B(n_548), .C(n_544), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_745), .B(n_607), .Y(n_856) );
BUFx8_ASAP7_75t_L g857 ( .A(n_730), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g858 ( .A(n_728), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_740), .Y(n_859) );
OAI22xp5_ASAP7_75t_SL g860 ( .A1(n_734), .A2(n_463), .B1(n_555), .B2(n_467), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g861 ( .A1(n_709), .A2(n_557), .B(n_553), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_726), .A2(n_562), .B1(n_566), .B2(n_558), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_774), .Y(n_863) );
INVxp67_ASAP7_75t_L g864 ( .A(n_752), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_711), .A2(n_574), .B(n_567), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_745), .B(n_454), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_735), .B(n_470), .Y(n_867) );
AOI21xp5_ASAP7_75t_L g868 ( .A1(n_712), .A2(n_578), .B(n_575), .Y(n_868) );
INVxp67_ASAP7_75t_L g869 ( .A(n_726), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g870 ( .A1(n_714), .A2(n_778), .B(n_781), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_778), .B(n_617), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_778), .B(n_617), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_723), .A2(n_511), .B1(n_563), .B2(n_526), .Y(n_873) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_756), .Y(n_874) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_721), .A2(n_580), .B(n_579), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g876 ( .A1(n_721), .A2(n_586), .B(n_584), .Y(n_876) );
INVx3_ASAP7_75t_L g877 ( .A(n_751), .Y(n_877) );
NAND3xp33_ASAP7_75t_L g878 ( .A(n_773), .B(n_593), .C(n_587), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_722), .B(n_594), .Y(n_879) );
AOI21xp5_ASAP7_75t_L g880 ( .A1(n_721), .A2(n_600), .B(n_599), .Y(n_880) );
OR2x2_ASAP7_75t_L g881 ( .A(n_710), .B(n_8), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_742), .A2(n_554), .B1(n_430), .B2(n_477), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_719), .B(n_552), .Y(n_883) );
INVx3_ASAP7_75t_L g884 ( .A(n_751), .Y(n_884) );
OAI22xp5_ASAP7_75t_SL g885 ( .A1(n_728), .A2(n_482), .B1(n_496), .B2(n_486), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_722), .B(n_603), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_751), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_722), .B(n_604), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_722), .B(n_605), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_722), .B(n_610), .Y(n_890) );
AOI21xp5_ASAP7_75t_L g891 ( .A1(n_721), .A2(n_614), .B(n_611), .Y(n_891) );
INVx4_ASAP7_75t_L g892 ( .A(n_751), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_710), .B(n_430), .Y(n_893) );
BUFx2_ASAP7_75t_L g894 ( .A(n_710), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_710), .B(n_430), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_736), .Y(n_896) );
OAI21x1_ASAP7_75t_L g897 ( .A1(n_721), .A2(n_694), .B(n_692), .Y(n_897) );
INVxp67_ASAP7_75t_SL g898 ( .A(n_733), .Y(n_898) );
OAI21xp5_ASAP7_75t_L g899 ( .A1(n_721), .A2(n_627), .B(n_623), .Y(n_899) );
NAND2x1p5_ASAP7_75t_L g900 ( .A(n_751), .B(n_602), .Y(n_900) );
INVx4_ASAP7_75t_L g901 ( .A(n_892), .Y(n_901) );
AOI21xp5_ASAP7_75t_L g902 ( .A1(n_785), .A2(n_698), .B(n_694), .Y(n_902) );
OAI21x1_ASAP7_75t_L g903 ( .A1(n_897), .A2(n_694), .B(n_692), .Y(n_903) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_879), .A2(n_591), .B1(n_506), .B2(n_509), .Y(n_904) );
OAI21xp5_ASAP7_75t_L g905 ( .A1(n_793), .A2(n_698), .B(n_695), .Y(n_905) );
BUFx6f_ASAP7_75t_L g906 ( .A(n_842), .Y(n_906) );
AND2x4_ASAP7_75t_L g907 ( .A(n_892), .B(n_431), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g908 ( .A1(n_794), .A2(n_698), .B(n_695), .Y(n_908) );
AO31x2_ASAP7_75t_L g909 ( .A1(n_822), .A2(n_670), .A3(n_654), .B(n_478), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_805), .B(n_798), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_792), .B(n_430), .Y(n_911) );
AOI21xp5_ASAP7_75t_L g912 ( .A1(n_899), .A2(n_576), .B(n_431), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_795), .Y(n_913) );
OAI21xp5_ASAP7_75t_L g914 ( .A1(n_875), .A2(n_520), .B(n_507), .Y(n_914) );
NAND2xp5_ASAP7_75t_SL g915 ( .A(n_894), .B(n_523), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_818), .A2(n_554), .B1(n_525), .B2(n_533), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_787), .B(n_554), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g918 ( .A1(n_870), .A2(n_545), .B(n_531), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g919 ( .A1(n_876), .A2(n_577), .B(n_550), .Y(n_919) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_880), .A2(n_589), .B(n_585), .Y(n_920) );
BUFx2_ASAP7_75t_L g921 ( .A(n_801), .Y(n_921) );
BUFx3_ASAP7_75t_L g922 ( .A(n_857), .Y(n_922) );
OA21x2_ASAP7_75t_L g923 ( .A1(n_791), .A2(n_598), .B(n_596), .Y(n_923) );
AOI21xp5_ASAP7_75t_L g924 ( .A1(n_891), .A2(n_608), .B(n_606), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_881), .B(n_9), .Y(n_925) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_821), .Y(n_926) );
A2O1A1Ixp33_ASAP7_75t_L g927 ( .A1(n_804), .A2(n_554), .B(n_535), .C(n_478), .Y(n_927) );
AOI221x1_ASAP7_75t_L g928 ( .A1(n_873), .A2(n_670), .B1(n_654), .B2(n_573), .C(n_601), .Y(n_928) );
BUFx2_ASAP7_75t_SL g929 ( .A(n_827), .Y(n_929) );
O2A1O1Ixp33_ASAP7_75t_L g930 ( .A1(n_834), .A2(n_12), .B(n_10), .C(n_11), .Y(n_930) );
AO32x2_ASAP7_75t_L g931 ( .A1(n_873), .A2(n_670), .A3(n_654), .B1(n_573), .B2(n_601), .Y(n_931) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_833), .A2(n_618), .B(n_613), .Y(n_932) );
NOR4xp25_ASAP7_75t_L g933 ( .A(n_836), .B(n_12), .C(n_10), .D(n_11), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_826), .B(n_13), .Y(n_934) );
CKINVDCx5p33_ASAP7_75t_R g935 ( .A(n_797), .Y(n_935) );
AO22x2_ASAP7_75t_L g936 ( .A1(n_878), .A2(n_15), .B1(n_13), .B2(n_14), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_879), .A2(n_630), .B1(n_622), .B2(n_535), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_788), .A2(n_796), .B(n_808), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_849), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_819), .B(n_15), .Y(n_940) );
NAND2x1p5_ASAP7_75t_L g941 ( .A(n_799), .B(n_573), .Y(n_941) );
OAI21xp5_ASAP7_75t_L g942 ( .A1(n_786), .A2(n_655), .B(n_654), .Y(n_942) );
BUFx2_ASAP7_75t_L g943 ( .A(n_857), .Y(n_943) );
AO31x2_ASAP7_75t_L g944 ( .A1(n_854), .A2(n_670), .A3(n_601), .B(n_573), .Y(n_944) );
BUFx3_ASAP7_75t_L g945 ( .A(n_893), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_886), .B(n_16), .Y(n_946) );
INVx2_ASAP7_75t_SL g947 ( .A(n_895), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_886), .B(n_16), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_888), .Y(n_949) );
AND2x4_ASAP7_75t_L g950 ( .A(n_898), .B(n_17), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g951 ( .A1(n_888), .A2(n_601), .B(n_655), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_889), .B(n_17), .Y(n_952) );
AOI21xp5_ASAP7_75t_SL g953 ( .A1(n_842), .A2(n_150), .B(n_148), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_852), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_889), .B(n_18), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_890), .A2(n_655), .B(n_156), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_858), .B(n_19), .Y(n_957) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_832), .Y(n_958) );
AOI21xp5_ASAP7_75t_L g959 ( .A1(n_890), .A2(n_843), .B(n_840), .Y(n_959) );
NOR2xp67_ASAP7_75t_L g960 ( .A(n_825), .B(n_20), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_835), .B(n_20), .Y(n_961) );
NOR2xp33_ASAP7_75t_L g962 ( .A(n_812), .B(n_21), .Y(n_962) );
AOI21xp5_ASAP7_75t_L g963 ( .A1(n_789), .A2(n_655), .B(n_157), .Y(n_963) );
A2O1A1Ixp33_ASAP7_75t_L g964 ( .A1(n_848), .A2(n_655), .B(n_23), .C(n_21), .Y(n_964) );
INVx2_ASAP7_75t_SL g965 ( .A(n_835), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g966 ( .A(n_809), .B(n_22), .Y(n_966) );
NAND3xp33_ASAP7_75t_L g967 ( .A(n_883), .B(n_817), .C(n_882), .Y(n_967) );
OAI21x1_ASAP7_75t_L g968 ( .A1(n_800), .A2(n_159), .B(n_153), .Y(n_968) );
AOI21xp5_ASAP7_75t_L g969 ( .A1(n_790), .A2(n_161), .B(n_160), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_859), .Y(n_970) );
BUFx6f_ASAP7_75t_L g971 ( .A(n_874), .Y(n_971) );
BUFx4f_ASAP7_75t_SL g972 ( .A(n_811), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_885), .Y(n_973) );
NAND2x1_ASAP7_75t_SL g974 ( .A(n_828), .B(n_22), .Y(n_974) );
INVx2_ASAP7_75t_SL g975 ( .A(n_900), .Y(n_975) );
AOI221xp5_ASAP7_75t_L g976 ( .A1(n_860), .A2(n_24), .B1(n_25), .B2(n_26), .C(n_27), .Y(n_976) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_814), .B(n_24), .Y(n_977) );
OAI21xp5_ASAP7_75t_L g978 ( .A1(n_869), .A2(n_165), .B(n_162), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_803), .A2(n_168), .B(n_166), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_896), .Y(n_980) );
AND3x4_ASAP7_75t_L g981 ( .A(n_847), .B(n_25), .C(n_26), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_831), .A2(n_30), .B1(n_28), .B2(n_29), .Y(n_982) );
AOI21xp5_ASAP7_75t_L g983 ( .A1(n_867), .A2(n_173), .B(n_171), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_841), .B(n_29), .Y(n_984) );
AOI221x1_ASAP7_75t_L g985 ( .A1(n_850), .A2(n_30), .B1(n_31), .B2(n_32), .C(n_33), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_851), .A2(n_34), .B1(n_31), .B2(n_33), .Y(n_986) );
HB1xp67_ASAP7_75t_L g987 ( .A(n_821), .Y(n_987) );
INVx3_ASAP7_75t_L g988 ( .A(n_799), .Y(n_988) );
OR2x2_ASAP7_75t_L g989 ( .A(n_820), .B(n_34), .Y(n_989) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_862), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_823), .B(n_35), .Y(n_991) );
CKINVDCx5p33_ASAP7_75t_R g992 ( .A(n_810), .Y(n_992) );
BUFx2_ASAP7_75t_L g993 ( .A(n_864), .Y(n_993) );
INVx6_ASAP7_75t_L g994 ( .A(n_874), .Y(n_994) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_829), .B(n_35), .Y(n_995) );
AOI21xp5_ASAP7_75t_L g996 ( .A1(n_837), .A2(n_187), .B(n_186), .Y(n_996) );
AO21x2_ASAP7_75t_L g997 ( .A1(n_855), .A2(n_190), .B(n_188), .Y(n_997) );
AO21x1_ASAP7_75t_L g998 ( .A1(n_900), .A2(n_200), .B(n_198), .Y(n_998) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_813), .B(n_36), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_802), .B(n_36), .Y(n_1000) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_802), .Y(n_1001) );
AOI21xp5_ASAP7_75t_L g1002 ( .A1(n_816), .A2(n_204), .B(n_201), .Y(n_1002) );
AO31x2_ASAP7_75t_L g1003 ( .A1(n_856), .A2(n_39), .A3(n_37), .B(n_38), .Y(n_1003) );
OAI21x1_ASAP7_75t_SL g1004 ( .A1(n_839), .A2(n_37), .B(n_38), .Y(n_1004) );
AOI21x1_ASAP7_75t_L g1005 ( .A1(n_844), .A2(n_846), .B(n_845), .Y(n_1005) );
BUFx3_ASAP7_75t_L g1006 ( .A(n_877), .Y(n_1006) );
AO31x2_ASAP7_75t_L g1007 ( .A1(n_830), .A2(n_44), .A3(n_41), .B(n_43), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g1008 ( .A(n_877), .Y(n_1008) );
AND2x2_ASAP7_75t_SL g1009 ( .A(n_874), .B(n_43), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_838), .B(n_44), .Y(n_1010) );
BUFx2_ASAP7_75t_L g1011 ( .A(n_884), .Y(n_1011) );
INVxp67_ASAP7_75t_SL g1012 ( .A(n_884), .Y(n_1012) );
OAI21xp5_ASAP7_75t_L g1013 ( .A1(n_853), .A2(n_206), .B(n_205), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_871), .B(n_45), .Y(n_1014) );
AOI21xp5_ASAP7_75t_L g1015 ( .A1(n_866), .A2(n_209), .B(n_207), .Y(n_1015) );
OA21x2_ASAP7_75t_L g1016 ( .A1(n_861), .A2(n_212), .B(n_211), .Y(n_1016) );
O2A1O1Ixp33_ASAP7_75t_L g1017 ( .A1(n_865), .A2(n_48), .B(n_46), .C(n_47), .Y(n_1017) );
BUFx6f_ASAP7_75t_L g1018 ( .A(n_806), .Y(n_1018) );
BUFx10_ASAP7_75t_L g1019 ( .A(n_872), .Y(n_1019) );
AOI31xp67_ASAP7_75t_L g1020 ( .A1(n_863), .A2(n_214), .A3(n_215), .B(n_213), .Y(n_1020) );
OAI21x1_ASAP7_75t_L g1021 ( .A1(n_868), .A2(n_218), .B(n_217), .Y(n_1021) );
A2O1A1Ixp33_ASAP7_75t_L g1022 ( .A1(n_815), .A2(n_46), .B(n_47), .C(n_48), .Y(n_1022) );
NOR2xp67_ASAP7_75t_L g1023 ( .A(n_887), .B(n_49), .Y(n_1023) );
AOI21xp5_ASAP7_75t_L g1024 ( .A1(n_824), .A2(n_225), .B(n_219), .Y(n_1024) );
BUFx8_ASAP7_75t_SL g1025 ( .A(n_894), .Y(n_1025) );
AO22x1_ASAP7_75t_SL g1026 ( .A1(n_832), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_1026) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_894), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_798), .B(n_50), .Y(n_1028) );
INVx3_ASAP7_75t_L g1029 ( .A(n_892), .Y(n_1029) );
OA21x2_ASAP7_75t_L g1030 ( .A1(n_899), .A2(n_240), .B(n_239), .Y(n_1030) );
AOI21xp5_ASAP7_75t_L g1031 ( .A1(n_785), .A2(n_242), .B(n_241), .Y(n_1031) );
A2O1A1Ixp33_ASAP7_75t_L g1032 ( .A1(n_807), .A2(n_51), .B(n_52), .C(n_54), .Y(n_1032) );
NOR2xp33_ASAP7_75t_L g1033 ( .A(n_798), .B(n_52), .Y(n_1033) );
AOI21xp5_ASAP7_75t_L g1034 ( .A1(n_785), .A2(n_244), .B(n_243), .Y(n_1034) );
A2O1A1Ixp33_ASAP7_75t_L g1035 ( .A1(n_807), .A2(n_54), .B(n_55), .C(n_56), .Y(n_1035) );
AND2x4_ASAP7_75t_L g1036 ( .A(n_892), .B(n_56), .Y(n_1036) );
INVx5_ASAP7_75t_L g1037 ( .A(n_892), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_805), .B(n_57), .Y(n_1038) );
OAI21x1_ASAP7_75t_L g1039 ( .A1(n_897), .A2(n_247), .B(n_246), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_849), .Y(n_1040) );
OAI22x1_ASAP7_75t_L g1041 ( .A1(n_894), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_1041) );
INVxp67_ASAP7_75t_L g1042 ( .A(n_993), .Y(n_1042) );
NAND2x1p5_ASAP7_75t_L g1043 ( .A(n_1037), .B(n_59), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_980), .Y(n_1044) );
OAI21xp5_ASAP7_75t_L g1045 ( .A1(n_959), .A2(n_60), .B(n_61), .Y(n_1045) );
AO31x2_ASAP7_75t_L g1046 ( .A1(n_928), .A2(n_62), .A3(n_63), .B(n_64), .Y(n_1046) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_922), .Y(n_1047) );
INVx2_ASAP7_75t_L g1048 ( .A(n_939), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1049 ( .A(n_1027), .Y(n_1049) );
OAI21x1_ASAP7_75t_L g1050 ( .A1(n_903), .A2(n_253), .B(n_251), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_970), .Y(n_1051) );
INVx3_ASAP7_75t_L g1052 ( .A(n_1037), .Y(n_1052) );
OAI21xp5_ASAP7_75t_L g1053 ( .A1(n_967), .A2(n_62), .B(n_63), .Y(n_1053) );
A2O1A1Ixp33_ASAP7_75t_L g1054 ( .A1(n_949), .A2(n_65), .B(n_66), .C(n_67), .Y(n_1054) );
AOI21xp33_ASAP7_75t_SL g1055 ( .A1(n_981), .A2(n_65), .B(n_66), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_910), .B(n_67), .Y(n_1056) );
NAND2xp5_ASAP7_75t_SL g1057 ( .A(n_1037), .B(n_69), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_950), .Y(n_1058) );
AOI21xp5_ASAP7_75t_L g1059 ( .A1(n_938), .A2(n_259), .B(n_257), .Y(n_1059) );
AOI21xp5_ASAP7_75t_L g1060 ( .A1(n_902), .A2(n_263), .B(n_261), .Y(n_1060) );
AND2x4_ASAP7_75t_L g1061 ( .A(n_901), .B(n_69), .Y(n_1061) );
AOI21xp5_ASAP7_75t_L g1062 ( .A1(n_905), .A2(n_268), .B(n_265), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_950), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_913), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1001), .B(n_71), .Y(n_1065) );
INVx3_ASAP7_75t_L g1066 ( .A(n_901), .Y(n_1066) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_1025), .Y(n_1067) );
OAI21x1_ASAP7_75t_L g1068 ( .A1(n_1039), .A2(n_271), .B(n_269), .Y(n_1068) );
OA21x2_ASAP7_75t_L g1069 ( .A1(n_968), .A2(n_276), .B(n_275), .Y(n_1069) );
OAI21x1_ASAP7_75t_SL g1070 ( .A1(n_978), .A2(n_73), .B(n_74), .Y(n_1070) );
BUFx6f_ASAP7_75t_L g1071 ( .A(n_906), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1038), .B(n_73), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1036), .Y(n_1073) );
OAI21xp5_ASAP7_75t_L g1074 ( .A1(n_999), .A2(n_74), .B(n_76), .Y(n_1074) );
AOI21xp5_ASAP7_75t_L g1075 ( .A1(n_951), .A2(n_281), .B(n_280), .Y(n_1075) );
OAI21x1_ASAP7_75t_L g1076 ( .A1(n_908), .A2(n_310), .B(n_410), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1036), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1078 ( .A1(n_990), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_965), .B(n_77), .Y(n_1079) );
INVx4_ASAP7_75t_L g1080 ( .A(n_1009), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1040), .Y(n_1081) );
INVx3_ASAP7_75t_L g1082 ( .A(n_1029), .Y(n_1082) );
CKINVDCx20_ASAP7_75t_R g1083 ( .A(n_943), .Y(n_1083) );
NOR2x1_ASAP7_75t_R g1084 ( .A(n_935), .B(n_78), .Y(n_1084) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_926), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_1033), .A2(n_992), .B1(n_984), .B2(n_934), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_987), .Y(n_1087) );
OR2x6_ASAP7_75t_L g1088 ( .A(n_929), .B(n_79), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_961), .Y(n_1089) );
OAI21xp5_ASAP7_75t_L g1090 ( .A1(n_991), .A2(n_80), .B(n_82), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_957), .B(n_80), .Y(n_1091) );
NAND4xp25_ASAP7_75t_L g1092 ( .A(n_960), .B(n_82), .C(n_83), .D(n_84), .Y(n_1092) );
NOR3xp33_ASAP7_75t_L g1093 ( .A(n_966), .B(n_83), .C(n_85), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_995), .B(n_85), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_954), .Y(n_1095) );
INVx2_ASAP7_75t_L g1096 ( .A(n_941), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1097 ( .A(n_921), .B(n_87), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_977), .A2(n_87), .B1(n_89), .B2(n_91), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_925), .B(n_89), .Y(n_1099) );
BUFx10_ASAP7_75t_L g1100 ( .A(n_907), .Y(n_1100) );
AO21x2_ASAP7_75t_L g1101 ( .A1(n_912), .A2(n_314), .B(n_409), .Y(n_1101) );
AND2x4_ASAP7_75t_L g1102 ( .A(n_1029), .B(n_1006), .Y(n_1102) );
AOI21xp5_ASAP7_75t_L g1103 ( .A1(n_942), .A2(n_313), .B(n_405), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_946), .Y(n_1104) );
AOI21xp5_ASAP7_75t_L g1105 ( .A1(n_956), .A2(n_311), .B(n_404), .Y(n_1105) );
OA21x2_ASAP7_75t_L g1106 ( .A1(n_985), .A2(n_307), .B(n_403), .Y(n_1106) );
OAI21x1_ASAP7_75t_L g1107 ( .A1(n_1031), .A2(n_306), .B(n_402), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_989), .B(n_91), .Y(n_1108) );
BUFx2_ASAP7_75t_L g1109 ( .A(n_907), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_948), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1007), .Y(n_1111) );
OAI21xp33_ASAP7_75t_SL g1112 ( .A1(n_974), .A2(n_92), .B(n_93), .Y(n_1112) );
CKINVDCx20_ASAP7_75t_R g1113 ( .A(n_958), .Y(n_1113) );
INVx2_ASAP7_75t_L g1114 ( .A(n_909), .Y(n_1114) );
OAI21xp5_ASAP7_75t_L g1115 ( .A1(n_952), .A2(n_93), .B(n_94), .Y(n_1115) );
AOI21xp5_ASAP7_75t_L g1116 ( .A1(n_955), .A2(n_319), .B(n_398), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1007), .Y(n_1117) );
A2O1A1Ixp33_ASAP7_75t_L g1118 ( .A1(n_930), .A2(n_94), .B(n_95), .C(n_96), .Y(n_1118) );
AO31x2_ASAP7_75t_L g1119 ( .A1(n_998), .A2(n_95), .A3(n_96), .B(n_97), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1007), .Y(n_1120) );
AND2x4_ASAP7_75t_L g1121 ( .A(n_975), .B(n_97), .Y(n_1121) );
OA21x2_ASAP7_75t_L g1122 ( .A1(n_1021), .A2(n_321), .B(n_397), .Y(n_1122) );
OAI21x1_ASAP7_75t_SL g1123 ( .A1(n_1013), .A2(n_98), .B(n_99), .Y(n_1123) );
BUFx2_ASAP7_75t_L g1124 ( .A(n_945), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1023), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1003), .Y(n_1126) );
AOI21xp33_ASAP7_75t_SL g1127 ( .A1(n_1041), .A2(n_98), .B(n_100), .Y(n_1127) );
OAI21x1_ASAP7_75t_L g1128 ( .A1(n_1034), .A2(n_324), .B(n_396), .Y(n_1128) );
AND2x4_ASAP7_75t_L g1129 ( .A(n_988), .B(n_101), .Y(n_1129) );
AOI22xp5_ASAP7_75t_L g1130 ( .A1(n_904), .A2(n_102), .B1(n_104), .B2(n_105), .Y(n_1130) );
NOR2xp33_ASAP7_75t_L g1131 ( .A(n_915), .B(n_972), .Y(n_1131) );
INVx4_ASAP7_75t_L g1132 ( .A(n_994), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_916), .B(n_102), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1003), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_973), .B(n_104), .Y(n_1135) );
AO21x2_ASAP7_75t_L g1136 ( .A1(n_927), .A2(n_325), .B(n_395), .Y(n_1136) );
AO21x2_ASAP7_75t_L g1137 ( .A1(n_911), .A2(n_323), .B(n_394), .Y(n_1137) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_963), .A2(n_320), .B(n_393), .Y(n_1138) );
AND2x4_ASAP7_75t_L g1139 ( .A(n_988), .B(n_105), .Y(n_1139) );
AND2x2_ASAP7_75t_SL g1140 ( .A(n_933), .B(n_1000), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_962), .B(n_106), .Y(n_1141) );
AOI22xp5_ASAP7_75t_L g1142 ( .A1(n_1028), .A2(n_106), .B1(n_107), .B2(n_109), .Y(n_1142) );
OA21x2_ASAP7_75t_L g1143 ( .A1(n_983), .A2(n_302), .B(n_391), .Y(n_1143) );
AOI21xp5_ASAP7_75t_L g1144 ( .A1(n_923), .A2(n_301), .B(n_390), .Y(n_1144) );
OA21x2_ASAP7_75t_L g1145 ( .A1(n_1015), .A2(n_299), .B(n_389), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g1146 ( .A(n_1011), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_936), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_936), .Y(n_1148) );
NAND2x1p5_ASAP7_75t_L g1149 ( .A(n_906), .B(n_107), .Y(n_1149) );
AOI21xp5_ASAP7_75t_L g1150 ( .A1(n_923), .A2(n_333), .B(n_387), .Y(n_1150) );
AO21x2_ASAP7_75t_L g1151 ( .A1(n_997), .A2(n_293), .B(n_386), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1004), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_976), .A2(n_109), .B1(n_110), .B2(n_111), .Y(n_1153) );
INVx3_ASAP7_75t_L g1154 ( .A(n_906), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_917), .B(n_111), .Y(n_1155) );
AND2x6_ASAP7_75t_L g1156 ( .A(n_971), .B(n_113), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1019), .B(n_113), .Y(n_1157) );
AO221x2_ASAP7_75t_L g1158 ( .A1(n_1026), .A2(n_114), .B1(n_116), .B2(n_117), .C(n_118), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_947), .B(n_116), .Y(n_1159) );
OAI21x1_ASAP7_75t_SL g1160 ( .A1(n_1030), .A2(n_117), .B(n_119), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1005), .Y(n_1161) );
NAND2x1_ASAP7_75t_L g1162 ( .A(n_994), .B(n_337), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_909), .Y(n_1163) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_986), .A2(n_119), .B1(n_120), .B2(n_122), .Y(n_1164) );
OA21x2_ASAP7_75t_L g1165 ( .A1(n_1032), .A2(n_338), .B(n_384), .Y(n_1165) );
AO21x2_ASAP7_75t_L g1166 ( .A1(n_997), .A2(n_336), .B(n_380), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_940), .B(n_122), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1010), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_937), .B(n_123), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_1014), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_909), .Y(n_1171) );
AO21x2_ASAP7_75t_L g1172 ( .A1(n_1035), .A2(n_340), .B(n_369), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1017), .Y(n_1173) );
OA21x2_ASAP7_75t_L g1174 ( .A1(n_1002), .A2(n_339), .B(n_368), .Y(n_1174) );
OA21x2_ASAP7_75t_L g1175 ( .A1(n_969), .A2(n_335), .B(n_366), .Y(n_1175) );
AOI21x1_ASAP7_75t_L g1176 ( .A1(n_1030), .A2(n_334), .B(n_365), .Y(n_1176) );
OAI21x1_ASAP7_75t_L g1177 ( .A1(n_1024), .A2(n_292), .B(n_357), .Y(n_1177) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_982), .A2(n_124), .B1(n_126), .B2(n_127), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1019), .B(n_126), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1022), .Y(n_1180) );
HB1xp67_ASAP7_75t_L g1181 ( .A(n_1008), .Y(n_1181) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1018), .Y(n_1182) );
CKINVDCx5p33_ASAP7_75t_R g1183 ( .A(n_1018), .Y(n_1183) );
OAI221xp5_ASAP7_75t_SL g1184 ( .A1(n_964), .A2(n_127), .B1(n_128), .B2(n_129), .C(n_130), .Y(n_1184) );
BUFx12f_ASAP7_75t_L g1185 ( .A(n_1018), .Y(n_1185) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_1012), .Y(n_1186) );
AOI21xp5_ASAP7_75t_L g1187 ( .A1(n_918), .A2(n_290), .B(n_354), .Y(n_1187) );
AOI21xp5_ASAP7_75t_L g1188 ( .A1(n_914), .A2(n_286), .B(n_353), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_932), .B(n_128), .Y(n_1189) );
BUFx4_ASAP7_75t_SL g1190 ( .A(n_953), .Y(n_1190) );
OA21x2_ASAP7_75t_L g1191 ( .A1(n_979), .A2(n_341), .B(n_351), .Y(n_1191) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_971), .A2(n_129), .B1(n_130), .B2(n_131), .Y(n_1192) );
INVx2_ASAP7_75t_L g1193 ( .A(n_944), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_919), .B(n_131), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_920), .B(n_133), .Y(n_1195) );
AND2x4_ASAP7_75t_L g1196 ( .A(n_971), .B(n_135), .Y(n_1196) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1161), .Y(n_1197) );
INVx2_ASAP7_75t_L g1198 ( .A(n_1161), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1044), .Y(n_1199) );
CKINVDCx11_ASAP7_75t_R g1200 ( .A(n_1083), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1051), .Y(n_1201) );
INVxp67_ASAP7_75t_L g1202 ( .A(n_1064), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1048), .B(n_931), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1114), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_1042), .Y(n_1205) );
INVx2_ASAP7_75t_L g1206 ( .A(n_1051), .Y(n_1206) );
INVx1_ASAP7_75t_SL g1207 ( .A(n_1183), .Y(n_1207) );
AND2x4_ASAP7_75t_L g1208 ( .A(n_1152), .B(n_944), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1081), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1095), .B(n_931), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1061), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1104), .B(n_944), .Y(n_1212) );
INVx3_ASAP7_75t_L g1213 ( .A(n_1185), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1111), .Y(n_1214) );
OR2x6_ASAP7_75t_L g1215 ( .A(n_1080), .B(n_1020), .Y(n_1215) );
INVx1_ASAP7_75t_SL g1216 ( .A(n_1124), .Y(n_1216) );
INVx2_ASAP7_75t_SL g1217 ( .A(n_1052), .Y(n_1217) );
INVxp67_ASAP7_75t_L g1218 ( .A(n_1049), .Y(n_1218) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1193), .Y(n_1219) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1163), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1061), .Y(n_1221) );
INVx3_ASAP7_75t_L g1222 ( .A(n_1052), .Y(n_1222) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1171), .Y(n_1223) );
AOI21x1_ASAP7_75t_L g1224 ( .A1(n_1176), .A2(n_1016), .B(n_996), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1121), .Y(n_1225) );
BUFx2_ASAP7_75t_L g1226 ( .A(n_1156), .Y(n_1226) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1071), .Y(n_1227) );
BUFx2_ASAP7_75t_L g1228 ( .A(n_1156), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1121), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1104), .B(n_135), .Y(n_1230) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1071), .Y(n_1231) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1071), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1129), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1086), .B(n_924), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1235 ( .A(n_1087), .Y(n_1235) );
BUFx2_ASAP7_75t_L g1236 ( .A(n_1156), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1129), .Y(n_1237) );
HB1xp67_ASAP7_75t_L g1238 ( .A(n_1085), .Y(n_1238) );
HB1xp67_ASAP7_75t_L g1239 ( .A(n_1088), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1110), .B(n_136), .Y(n_1240) );
INVx2_ASAP7_75t_L g1241 ( .A(n_1160), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1139), .Y(n_1242) );
AO21x2_ASAP7_75t_L g1243 ( .A1(n_1134), .A2(n_136), .B(n_137), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1110), .B(n_283), .Y(n_1244) );
INVx2_ASAP7_75t_L g1245 ( .A(n_1050), .Y(n_1245) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1122), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1089), .B(n_284), .Y(n_1247) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1122), .Y(n_1248) );
HB1xp67_ASAP7_75t_L g1249 ( .A(n_1088), .Y(n_1249) );
AOI221x1_ASAP7_75t_L g1250 ( .A1(n_1144), .A2(n_342), .B1(n_343), .B2(n_344), .C(n_348), .Y(n_1250) );
INVx1_ASAP7_75t_SL g1251 ( .A(n_1047), .Y(n_1251) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1046), .Y(n_1252) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1046), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1117), .Y(n_1254) );
OR2x6_ASAP7_75t_L g1255 ( .A(n_1080), .B(n_415), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1120), .Y(n_1256) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_1158), .A2(n_1093), .B1(n_1173), .B2(n_1141), .Y(n_1257) );
NAND3xp33_ASAP7_75t_L g1258 ( .A(n_1127), .B(n_1055), .C(n_1112), .Y(n_1258) );
AO21x2_ASAP7_75t_L g1259 ( .A1(n_1070), .A2(n_1123), .B(n_1045), .Y(n_1259) );
NAND2x1p5_ASAP7_75t_L g1260 ( .A(n_1154), .B(n_1066), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1139), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1147), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1168), .B(n_1140), .Y(n_1263) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_1186), .Y(n_1264) );
HB1xp67_ASAP7_75t_L g1265 ( .A(n_1181), .Y(n_1265) );
INVxp67_ASAP7_75t_SL g1266 ( .A(n_1146), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1148), .B(n_1180), .Y(n_1267) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1159), .Y(n_1268) );
BUFx2_ASAP7_75t_L g1269 ( .A(n_1156), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1115), .B(n_1158), .Y(n_1270) );
AO21x2_ASAP7_75t_L g1271 ( .A1(n_1150), .A2(n_1166), .B(n_1151), .Y(n_1271) );
AO21x2_ASAP7_75t_L g1272 ( .A1(n_1151), .A2(n_1166), .B(n_1053), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1058), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1063), .Y(n_1274) );
INVx3_ASAP7_75t_L g1275 ( .A(n_1066), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_1092), .A2(n_1065), .B1(n_1077), .B2(n_1073), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g1277 ( .A1(n_1043), .A2(n_1169), .B1(n_1153), .B2(n_1170), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1196), .B(n_1074), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1056), .Y(n_1279) );
HB1xp67_ASAP7_75t_L g1280 ( .A(n_1109), .Y(n_1280) );
OAI21x1_ASAP7_75t_SL g1281 ( .A1(n_1103), .A2(n_1090), .B(n_1188), .Y(n_1281) );
BUFx2_ASAP7_75t_SL g1282 ( .A(n_1100), .Y(n_1282) );
INVx4_ASAP7_75t_SL g1283 ( .A(n_1196), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1072), .B(n_1108), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1079), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1099), .Y(n_1286) );
AO21x2_ASAP7_75t_L g1287 ( .A1(n_1101), .A2(n_1172), .B(n_1137), .Y(n_1287) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1082), .B(n_1182), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1091), .B(n_1097), .Y(n_1289) );
BUFx6f_ASAP7_75t_L g1290 ( .A(n_1154), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1119), .Y(n_1291) );
OA21x2_ASAP7_75t_L g1292 ( .A1(n_1068), .A2(n_1076), .B(n_1059), .Y(n_1292) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1106), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1082), .B(n_1119), .Y(n_1294) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1106), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1119), .B(n_1054), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1094), .B(n_1167), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1149), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1100), .B(n_1102), .Y(n_1299) );
CKINVDCx16_ASAP7_75t_R g1300 ( .A(n_1067), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1125), .Y(n_1301) );
INVx3_ASAP7_75t_L g1302 ( .A(n_1096), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1195), .Y(n_1303) );
AO21x2_ASAP7_75t_L g1304 ( .A1(n_1101), .A2(n_1172), .B(n_1137), .Y(n_1304) );
AND2x4_ASAP7_75t_L g1305 ( .A(n_1102), .B(n_1132), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1142), .B(n_1118), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1057), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1157), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1179), .B(n_1098), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1069), .Y(n_1310) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1165), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1155), .Y(n_1312) );
INVx2_ASAP7_75t_L g1313 ( .A(n_1174), .Y(n_1313) );
INVx4_ASAP7_75t_L g1314 ( .A(n_1132), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1131), .B(n_1133), .Y(n_1315) );
AOI21x1_ASAP7_75t_L g1316 ( .A1(n_1062), .A2(n_1143), .B(n_1145), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1078), .B(n_1130), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1194), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1189), .B(n_1135), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1192), .Y(n_1320) );
AND2x4_ASAP7_75t_L g1321 ( .A(n_1136), .B(n_1116), .Y(n_1321) );
HB1xp67_ASAP7_75t_L g1322 ( .A(n_1164), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1178), .Y(n_1323) );
INVx2_ASAP7_75t_L g1324 ( .A(n_1136), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1184), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1084), .Y(n_1326) );
OAI21x1_ASAP7_75t_L g1327 ( .A1(n_1177), .A2(n_1128), .B(n_1107), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1175), .B(n_1191), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1175), .B(n_1191), .Y(n_1329) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1162), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1060), .B(n_1187), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1075), .B(n_1138), .Y(n_1332) );
INVx2_ASAP7_75t_L g1333 ( .A(n_1190), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1105), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1113), .B(n_1048), .Y(n_1335) );
INVx2_ASAP7_75t_SL g1336 ( .A(n_1185), .Y(n_1336) );
INVx2_ASAP7_75t_SL g1337 ( .A(n_1185), .Y(n_1337) );
AO21x2_ASAP7_75t_L g1338 ( .A1(n_1160), .A2(n_1161), .B(n_1126), .Y(n_1338) );
INVx2_ASAP7_75t_SL g1339 ( .A(n_1185), .Y(n_1339) );
BUFx2_ASAP7_75t_L g1340 ( .A(n_1156), .Y(n_1340) );
OA21x2_ASAP7_75t_L g1341 ( .A1(n_1161), .A2(n_1171), .B(n_1163), .Y(n_1341) );
INVx2_ASAP7_75t_L g1342 ( .A(n_1161), .Y(n_1342) );
INVx3_ASAP7_75t_L g1343 ( .A(n_1185), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1303), .B(n_1199), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1230), .B(n_1240), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1201), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1209), .Y(n_1347) );
AND2x4_ASAP7_75t_L g1348 ( .A(n_1214), .B(n_1254), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1206), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1319), .B(n_1335), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1206), .Y(n_1351) );
HB1xp67_ASAP7_75t_L g1352 ( .A(n_1220), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1264), .Y(n_1353) );
AND2x4_ASAP7_75t_L g1354 ( .A(n_1214), .B(n_1254), .Y(n_1354) );
INVxp67_ASAP7_75t_SL g1355 ( .A(n_1204), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1273), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1319), .B(n_1335), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1286), .B(n_1263), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1263), .B(n_1238), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1274), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1267), .B(n_1212), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1230), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1240), .Y(n_1363) );
INVx3_ASAP7_75t_L g1364 ( .A(n_1314), .Y(n_1364) );
HB1xp67_ASAP7_75t_L g1365 ( .A(n_1223), .Y(n_1365) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1262), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1308), .B(n_1265), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1301), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1256), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1256), .Y(n_1370) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1266), .B(n_1235), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1299), .B(n_1216), .Y(n_1372) );
INVx4_ASAP7_75t_L g1373 ( .A(n_1255), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1225), .Y(n_1374) );
HB1xp67_ASAP7_75t_L g1375 ( .A(n_1223), .Y(n_1375) );
AND2x4_ASAP7_75t_L g1376 ( .A(n_1267), .B(n_1212), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1270), .B(n_1257), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1270), .B(n_1279), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1229), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1299), .B(n_1207), .Y(n_1380) );
HB1xp67_ASAP7_75t_L g1381 ( .A(n_1204), .Y(n_1381) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1197), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1211), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1336), .B(n_1337), .Y(n_1384) );
OR2x2_ASAP7_75t_L g1385 ( .A(n_1202), .B(n_1218), .Y(n_1385) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1205), .B(n_1280), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1221), .Y(n_1387) );
OR2x2_ASAP7_75t_L g1388 ( .A(n_1251), .B(n_1217), .Y(n_1388) );
OR2x6_ASAP7_75t_L g1389 ( .A(n_1226), .B(n_1228), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1243), .Y(n_1390) );
HB1xp67_ASAP7_75t_L g1391 ( .A(n_1219), .Y(n_1391) );
INVx2_ASAP7_75t_L g1392 ( .A(n_1198), .Y(n_1392) );
BUFx2_ASAP7_75t_L g1393 ( .A(n_1305), .Y(n_1393) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1243), .Y(n_1394) );
BUFx2_ASAP7_75t_L g1395 ( .A(n_1305), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1243), .Y(n_1396) );
INVx2_ASAP7_75t_L g1397 ( .A(n_1198), .Y(n_1397) );
HB1xp67_ASAP7_75t_L g1398 ( .A(n_1219), .Y(n_1398) );
INVx3_ASAP7_75t_L g1399 ( .A(n_1314), .Y(n_1399) );
INVx2_ASAP7_75t_L g1400 ( .A(n_1342), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1342), .Y(n_1401) );
HB1xp67_ASAP7_75t_L g1402 ( .A(n_1341), .Y(n_1402) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1341), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1336), .B(n_1337), .Y(n_1404) );
NOR2x1_ASAP7_75t_SL g1405 ( .A(n_1255), .B(n_1282), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1233), .Y(n_1406) );
NAND2x1p5_ASAP7_75t_SL g1407 ( .A(n_1333), .B(n_1306), .Y(n_1407) );
AND2x4_ASAP7_75t_L g1408 ( .A(n_1226), .B(n_1228), .Y(n_1408) );
INVx2_ASAP7_75t_L g1409 ( .A(n_1341), .Y(n_1409) );
BUFx6f_ASAP7_75t_L g1410 ( .A(n_1290), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1294), .B(n_1291), .Y(n_1411) );
NAND2x1_ASAP7_75t_L g1412 ( .A(n_1236), .B(n_1269), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1339), .B(n_1305), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1339), .B(n_1289), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1237), .Y(n_1415) );
HB1xp67_ASAP7_75t_L g1416 ( .A(n_1338), .Y(n_1416) );
BUFx2_ASAP7_75t_L g1417 ( .A(n_1255), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1217), .B(n_1282), .Y(n_1418) );
BUFx2_ASAP7_75t_L g1419 ( .A(n_1255), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1242), .Y(n_1420) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1261), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1318), .B(n_1325), .Y(n_1422) );
HB1xp67_ASAP7_75t_L g1423 ( .A(n_1338), .Y(n_1423) );
INVx3_ASAP7_75t_L g1424 ( .A(n_1314), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1268), .Y(n_1425) );
NOR2x1_ASAP7_75t_SL g1426 ( .A(n_1333), .B(n_1298), .Y(n_1426) );
NAND2x1p5_ASAP7_75t_SL g1427 ( .A(n_1306), .B(n_1317), .Y(n_1427) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1244), .Y(n_1428) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1244), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1430 ( .A(n_1323), .B(n_1276), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1317), .B(n_1285), .Y(n_1431) );
INVx2_ASAP7_75t_L g1432 ( .A(n_1338), .Y(n_1432) );
OR2x2_ASAP7_75t_L g1433 ( .A(n_1239), .B(n_1249), .Y(n_1433) );
INVx2_ASAP7_75t_L g1434 ( .A(n_1203), .Y(n_1434) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1222), .B(n_1288), .Y(n_1435) );
HB1xp67_ASAP7_75t_L g1436 ( .A(n_1208), .Y(n_1436) );
OR2x2_ASAP7_75t_L g1437 ( .A(n_1222), .B(n_1288), .Y(n_1437) );
AND2x4_ASAP7_75t_L g1438 ( .A(n_1236), .B(n_1269), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1315), .B(n_1222), .Y(n_1439) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1302), .Y(n_1440) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1302), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1213), .B(n_1343), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1302), .Y(n_1443) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1210), .Y(n_1444) );
INVx2_ASAP7_75t_SL g1445 ( .A(n_1275), .Y(n_1445) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1284), .B(n_1275), .Y(n_1446) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1343), .B(n_1213), .Y(n_1447) );
AO21x2_ASAP7_75t_L g1448 ( .A1(n_1310), .A2(n_1316), .B(n_1224), .Y(n_1448) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1210), .Y(n_1449) );
INVxp67_ASAP7_75t_L g1450 ( .A(n_1340), .Y(n_1450) );
AND2x4_ASAP7_75t_L g1451 ( .A(n_1340), .B(n_1208), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1452 ( .A(n_1284), .B(n_1297), .Y(n_1452) );
INVx2_ASAP7_75t_L g1453 ( .A(n_1208), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1343), .B(n_1213), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1275), .Y(n_1455) );
NAND2xp5_ASAP7_75t_SL g1456 ( .A(n_1278), .B(n_1283), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1309), .B(n_1247), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1309), .B(n_1247), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1278), .B(n_1297), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1234), .B(n_1326), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1322), .B(n_1312), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1312), .B(n_1260), .Y(n_1462) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1260), .B(n_1300), .Y(n_1463) );
INVx5_ASAP7_75t_L g1464 ( .A(n_1290), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1277), .B(n_1320), .Y(n_1465) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1294), .B(n_1296), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1298), .Y(n_1467) );
OR2x2_ASAP7_75t_L g1468 ( .A(n_1260), .B(n_1232), .Y(n_1468) );
OAI21xp33_ASAP7_75t_L g1469 ( .A1(n_1258), .A2(n_1296), .B(n_1307), .Y(n_1469) );
AOI22xp33_ASAP7_75t_L g1470 ( .A1(n_1259), .A2(n_1331), .B1(n_1332), .B2(n_1241), .Y(n_1470) );
NOR2xp67_ASAP7_75t_L g1471 ( .A(n_1252), .B(n_1253), .Y(n_1471) );
AND2x4_ASAP7_75t_L g1472 ( .A(n_1283), .B(n_1241), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1283), .B(n_1200), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1369), .Y(n_1474) );
AND2x4_ASAP7_75t_L g1475 ( .A(n_1453), .B(n_1283), .Y(n_1475) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1368), .Y(n_1476) );
INVx3_ASAP7_75t_L g1477 ( .A(n_1373), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1461), .B(n_1259), .Y(n_1478) );
HB1xp67_ASAP7_75t_L g1479 ( .A(n_1371), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1361), .B(n_1215), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1361), .B(n_1466), .Y(n_1481) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1347), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1466), .B(n_1215), .Y(n_1483) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1376), .B(n_1215), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1376), .B(n_1215), .Y(n_1485) );
NAND2xp5_ASAP7_75t_L g1486 ( .A(n_1431), .B(n_1259), .Y(n_1486) );
INVx2_ASAP7_75t_L g1487 ( .A(n_1403), .Y(n_1487) );
INVx2_ASAP7_75t_L g1488 ( .A(n_1403), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_1376), .B(n_1310), .Y(n_1489) );
NOR2xp67_ASAP7_75t_SL g1490 ( .A(n_1373), .B(n_1330), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1411), .B(n_1324), .Y(n_1491) );
INVx1_ASAP7_75t_SL g1492 ( .A(n_1384), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1411), .B(n_1324), .Y(n_1493) );
INVx2_ASAP7_75t_L g1494 ( .A(n_1409), .Y(n_1494) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1459), .B(n_1227), .Y(n_1495) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1444), .B(n_1328), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1352), .B(n_1232), .Y(n_1497) );
OR2x2_ASAP7_75t_L g1498 ( .A(n_1352), .B(n_1231), .Y(n_1498) );
NOR2xp67_ASAP7_75t_L g1499 ( .A(n_1373), .B(n_1321), .Y(n_1499) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1449), .B(n_1329), .Y(n_1500) );
INVx2_ASAP7_75t_L g1501 ( .A(n_1409), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1353), .Y(n_1502) );
AND2x2_ASAP7_75t_L g1503 ( .A(n_1434), .B(n_1329), .Y(n_1503) );
OR2x2_ASAP7_75t_L g1504 ( .A(n_1365), .B(n_1231), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1434), .B(n_1328), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1348), .B(n_1311), .Y(n_1506) );
HB1xp67_ASAP7_75t_L g1507 ( .A(n_1386), .Y(n_1507) );
BUFx2_ASAP7_75t_L g1508 ( .A(n_1417), .Y(n_1508) );
OR2x2_ASAP7_75t_L g1509 ( .A(n_1365), .B(n_1227), .Y(n_1509) );
HB1xp67_ASAP7_75t_L g1510 ( .A(n_1375), .Y(n_1510) );
HB1xp67_ASAP7_75t_L g1511 ( .A(n_1375), .Y(n_1511) );
BUFx2_ASAP7_75t_L g1512 ( .A(n_1419), .Y(n_1512) );
OR2x2_ASAP7_75t_L g1513 ( .A(n_1452), .B(n_1311), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1348), .B(n_1293), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1348), .B(n_1295), .Y(n_1515) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_1350), .B(n_1290), .Y(n_1516) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1425), .Y(n_1517) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1370), .Y(n_1518) );
HB1xp67_ASAP7_75t_L g1519 ( .A(n_1388), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1354), .B(n_1295), .Y(n_1520) );
INVxp67_ASAP7_75t_SL g1521 ( .A(n_1381), .Y(n_1521) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1401), .Y(n_1522) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1354), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1354), .B(n_1313), .Y(n_1524) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1346), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1391), .B(n_1398), .Y(n_1526) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1356), .Y(n_1527) );
HB1xp67_ASAP7_75t_L g1528 ( .A(n_1398), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g1529 ( .A(n_1357), .B(n_1290), .Y(n_1529) );
HB1xp67_ASAP7_75t_L g1530 ( .A(n_1446), .Y(n_1530) );
NAND2xp5_ASAP7_75t_L g1531 ( .A(n_1358), .B(n_1290), .Y(n_1531) );
BUFx3_ASAP7_75t_L g1532 ( .A(n_1364), .Y(n_1532) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1360), .Y(n_1533) );
INVx1_ASAP7_75t_SL g1534 ( .A(n_1404), .Y(n_1534) );
OR2x2_ASAP7_75t_L g1535 ( .A(n_1378), .B(n_1248), .Y(n_1535) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1344), .Y(n_1536) );
OR2x2_ASAP7_75t_L g1537 ( .A(n_1366), .B(n_1246), .Y(n_1537) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1367), .Y(n_1538) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1467), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_1362), .B(n_1200), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_1363), .B(n_1272), .Y(n_1541) );
OR2x2_ASAP7_75t_L g1542 ( .A(n_1465), .B(n_1304), .Y(n_1542) );
INVxp67_ASAP7_75t_L g1543 ( .A(n_1372), .Y(n_1543) );
INVxp67_ASAP7_75t_L g1544 ( .A(n_1414), .Y(n_1544) );
INVx3_ASAP7_75t_L g1545 ( .A(n_1472), .Y(n_1545) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1349), .Y(n_1546) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1351), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1383), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1382), .B(n_1304), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1550 ( .A(n_1382), .B(n_1304), .Y(n_1550) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1387), .Y(n_1551) );
HB1xp67_ASAP7_75t_L g1552 ( .A(n_1364), .Y(n_1552) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1406), .Y(n_1553) );
HB1xp67_ASAP7_75t_L g1554 ( .A(n_1399), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1392), .B(n_1287), .Y(n_1555) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1392), .B(n_1287), .Y(n_1556) );
AND2x4_ASAP7_75t_SL g1557 ( .A(n_1399), .B(n_1330), .Y(n_1557) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1415), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1397), .B(n_1287), .Y(n_1559) );
OR2x2_ASAP7_75t_SL g1560 ( .A(n_1436), .B(n_1292), .Y(n_1560) );
INVx3_ASAP7_75t_L g1561 ( .A(n_1472), .Y(n_1561) );
BUFx2_ASAP7_75t_L g1562 ( .A(n_1389), .Y(n_1562) );
AND2x4_ASAP7_75t_L g1563 ( .A(n_1451), .B(n_1321), .Y(n_1563) );
OR2x2_ASAP7_75t_L g1564 ( .A(n_1427), .B(n_1272), .Y(n_1564) );
NAND2xp5_ASAP7_75t_SL g1565 ( .A(n_1424), .B(n_1281), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1400), .B(n_1272), .Y(n_1566) );
INVxp67_ASAP7_75t_L g1567 ( .A(n_1426), .Y(n_1567) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1400), .Y(n_1568) );
NAND2xp5_ASAP7_75t_SL g1569 ( .A(n_1567), .B(n_1424), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1496), .B(n_1390), .Y(n_1570) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1496), .B(n_1394), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1572 ( .A(n_1481), .B(n_1359), .Y(n_1572) );
INVx2_ASAP7_75t_L g1573 ( .A(n_1526), .Y(n_1573) );
INVx2_ASAP7_75t_L g1574 ( .A(n_1526), .Y(n_1574) );
INVx2_ASAP7_75t_L g1575 ( .A(n_1528), .Y(n_1575) );
INVx4_ASAP7_75t_L g1576 ( .A(n_1532), .Y(n_1576) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1476), .Y(n_1577) );
INVx3_ASAP7_75t_L g1578 ( .A(n_1532), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1481), .B(n_1380), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1543), .B(n_1519), .Y(n_1580) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1482), .Y(n_1581) );
NAND2xp5_ASAP7_75t_L g1582 ( .A(n_1500), .B(n_1486), .Y(n_1582) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1527), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1500), .B(n_1396), .Y(n_1584) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1533), .Y(n_1585) );
NAND2xp5_ASAP7_75t_SL g1586 ( .A(n_1552), .B(n_1418), .Y(n_1586) );
AND2x4_ASAP7_75t_L g1587 ( .A(n_1562), .B(n_1451), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1588 ( .A(n_1536), .B(n_1422), .Y(n_1588) );
OR2x2_ASAP7_75t_L g1589 ( .A(n_1479), .B(n_1436), .Y(n_1589) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1480), .B(n_1460), .Y(n_1590) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1517), .Y(n_1591) );
AOI32xp33_ASAP7_75t_L g1592 ( .A1(n_1492), .A2(n_1473), .A3(n_1463), .B1(n_1377), .B2(n_1457), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g1593 ( .A(n_1522), .B(n_1469), .Y(n_1593) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1525), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1480), .B(n_1451), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1530), .B(n_1439), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1597 ( .A(n_1522), .B(n_1402), .Y(n_1597) );
INVx2_ASAP7_75t_L g1598 ( .A(n_1510), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1534), .B(n_1433), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1474), .B(n_1402), .Y(n_1600) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1474), .B(n_1470), .Y(n_1601) );
INVxp67_ASAP7_75t_SL g1602 ( .A(n_1521), .Y(n_1602) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1539), .Y(n_1603) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1502), .Y(n_1604) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1518), .Y(n_1605) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1518), .Y(n_1606) );
NAND2xp5_ASAP7_75t_SL g1607 ( .A(n_1554), .B(n_1393), .Y(n_1607) );
NAND2x1p5_ASAP7_75t_L g1608 ( .A(n_1490), .B(n_1412), .Y(n_1608) );
BUFx2_ASAP7_75t_L g1609 ( .A(n_1511), .Y(n_1609) );
INVx2_ASAP7_75t_SL g1610 ( .A(n_1507), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1483), .B(n_1395), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1483), .B(n_1408), .Y(n_1612) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1548), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_1546), .B(n_1470), .Y(n_1614) );
NAND2xp5_ASAP7_75t_L g1615 ( .A(n_1547), .B(n_1430), .Y(n_1615) );
OR2x2_ASAP7_75t_L g1616 ( .A(n_1538), .B(n_1385), .Y(n_1616) );
INVx2_ASAP7_75t_L g1617 ( .A(n_1497), .Y(n_1617) );
INVx2_ASAP7_75t_L g1618 ( .A(n_1497), .Y(n_1618) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1551), .Y(n_1619) );
INVxp67_ASAP7_75t_L g1620 ( .A(n_1478), .Y(n_1620) );
NOR2x1p5_ASAP7_75t_L g1621 ( .A(n_1477), .B(n_1438), .Y(n_1621) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1553), .Y(n_1622) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1558), .Y(n_1623) );
HB1xp67_ASAP7_75t_L g1624 ( .A(n_1498), .Y(n_1624) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1535), .Y(n_1625) );
OR2x2_ASAP7_75t_L g1626 ( .A(n_1535), .B(n_1355), .Y(n_1626) );
INVx1_ASAP7_75t_L g1627 ( .A(n_1537), .Y(n_1627) );
NAND2xp5_ASAP7_75t_L g1628 ( .A(n_1541), .B(n_1374), .Y(n_1628) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1537), .Y(n_1629) );
OR2x2_ASAP7_75t_L g1630 ( .A(n_1495), .B(n_1355), .Y(n_1630) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1513), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1489), .B(n_1438), .Y(n_1632) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1513), .Y(n_1633) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1523), .Y(n_1634) );
OR2x2_ASAP7_75t_L g1635 ( .A(n_1544), .B(n_1437), .Y(n_1635) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1542), .B(n_1379), .Y(n_1636) );
OR2x2_ASAP7_75t_L g1637 ( .A(n_1516), .B(n_1435), .Y(n_1637) );
NOR2x1p5_ASAP7_75t_L g1638 ( .A(n_1477), .B(n_1438), .Y(n_1638) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1489), .B(n_1408), .Y(n_1639) );
NOR2xp33_ASAP7_75t_L g1640 ( .A(n_1540), .B(n_1413), .Y(n_1640) );
AND2x2_ASAP7_75t_L g1641 ( .A(n_1484), .B(n_1408), .Y(n_1641) );
AND2x4_ASAP7_75t_L g1642 ( .A(n_1562), .B(n_1405), .Y(n_1642) );
NAND2xp5_ASAP7_75t_L g1643 ( .A(n_1542), .B(n_1427), .Y(n_1643) );
INVx2_ASAP7_75t_SL g1644 ( .A(n_1576), .Y(n_1644) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1577), .Y(n_1645) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1581), .Y(n_1646) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1583), .Y(n_1647) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1620), .B(n_1523), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1649 ( .A(n_1596), .B(n_1484), .Y(n_1649) );
HB1xp67_ASAP7_75t_L g1650 ( .A(n_1624), .Y(n_1650) );
INVx2_ASAP7_75t_L g1651 ( .A(n_1634), .Y(n_1651) );
INVx2_ASAP7_75t_SL g1652 ( .A(n_1576), .Y(n_1652) );
NOR2xp33_ASAP7_75t_L g1653 ( .A(n_1588), .B(n_1508), .Y(n_1653) );
AND2x2_ASAP7_75t_SL g1654 ( .A(n_1642), .B(n_1508), .Y(n_1654) );
NAND2xp5_ASAP7_75t_L g1655 ( .A(n_1620), .B(n_1503), .Y(n_1655) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1585), .Y(n_1656) );
OR2x2_ASAP7_75t_L g1657 ( .A(n_1582), .B(n_1498), .Y(n_1657) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1591), .Y(n_1658) );
INVx1_ASAP7_75t_SL g1659 ( .A(n_1599), .Y(n_1659) );
OR2x2_ASAP7_75t_L g1660 ( .A(n_1582), .B(n_1504), .Y(n_1660) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_1632), .B(n_1485), .Y(n_1661) );
INVx2_ASAP7_75t_L g1662 ( .A(n_1609), .Y(n_1662) );
OR2x6_ASAP7_75t_L g1663 ( .A(n_1608), .B(n_1389), .Y(n_1663) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_1588), .B(n_1503), .Y(n_1664) );
OR2x2_ASAP7_75t_L g1665 ( .A(n_1624), .B(n_1504), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1666 ( .A(n_1631), .B(n_1505), .Y(n_1666) );
INVxp67_ASAP7_75t_L g1667 ( .A(n_1602), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_1639), .B(n_1485), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1633), .B(n_1505), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1670 ( .A(n_1572), .B(n_1563), .Y(n_1670) );
NAND2xp33_ASAP7_75t_L g1671 ( .A(n_1621), .B(n_1477), .Y(n_1671) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_1625), .B(n_1491), .Y(n_1672) );
INVx2_ASAP7_75t_L g1673 ( .A(n_1605), .Y(n_1673) );
NOR2xp33_ASAP7_75t_L g1674 ( .A(n_1610), .B(n_1512), .Y(n_1674) );
INVxp67_ASAP7_75t_L g1675 ( .A(n_1602), .Y(n_1675) );
INVx2_ASAP7_75t_L g1676 ( .A(n_1626), .Y(n_1676) );
NAND2xp5_ASAP7_75t_L g1677 ( .A(n_1636), .B(n_1491), .Y(n_1677) );
INVxp67_ASAP7_75t_L g1678 ( .A(n_1575), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_1636), .B(n_1493), .Y(n_1679) );
OAI21xp33_ASAP7_75t_L g1680 ( .A1(n_1592), .A2(n_1564), .B(n_1563), .Y(n_1680) );
NAND2xp5_ASAP7_75t_L g1681 ( .A(n_1615), .B(n_1493), .Y(n_1681) );
AND2x2_ASAP7_75t_L g1682 ( .A(n_1590), .B(n_1563), .Y(n_1682) );
NAND2x1p5_ASAP7_75t_L g1683 ( .A(n_1578), .B(n_1490), .Y(n_1683) );
INVxp67_ASAP7_75t_L g1684 ( .A(n_1598), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1641), .B(n_1512), .Y(n_1685) );
NAND2xp5_ASAP7_75t_L g1686 ( .A(n_1615), .B(n_1529), .Y(n_1686) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1570), .B(n_1549), .Y(n_1687) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1594), .Y(n_1688) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1613), .Y(n_1689) );
OAI22xp33_ASAP7_75t_SL g1690 ( .A1(n_1586), .A2(n_1456), .B1(n_1565), .B2(n_1389), .Y(n_1690) );
AOI221xp5_ASAP7_75t_L g1691 ( .A1(n_1680), .A2(n_1643), .B1(n_1580), .B2(n_1604), .C(n_1619), .Y(n_1691) );
OAI322xp33_ASAP7_75t_L g1692 ( .A1(n_1667), .A2(n_1589), .A3(n_1643), .B1(n_1635), .B2(n_1616), .C1(n_1584), .C2(n_1570), .Y(n_1692) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1648), .Y(n_1693) );
NAND2xp5_ASAP7_75t_L g1694 ( .A(n_1650), .B(n_1601), .Y(n_1694) );
INVxp67_ASAP7_75t_SL g1695 ( .A(n_1667), .Y(n_1695) );
NOR2xp33_ASAP7_75t_L g1696 ( .A(n_1659), .B(n_1579), .Y(n_1696) );
OR2x2_ASAP7_75t_L g1697 ( .A(n_1687), .B(n_1573), .Y(n_1697) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1650), .B(n_1601), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_1670), .B(n_1595), .Y(n_1699) );
AOI22xp5_ASAP7_75t_L g1700 ( .A1(n_1653), .A2(n_1640), .B1(n_1587), .B2(n_1611), .Y(n_1700) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1653), .B(n_1627), .Y(n_1701) );
O2A1O1Ixp33_ASAP7_75t_L g1702 ( .A1(n_1690), .A2(n_1569), .B(n_1454), .C(n_1447), .Y(n_1702) );
INVx1_ASAP7_75t_SL g1703 ( .A(n_1644), .Y(n_1703) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1657), .Y(n_1704) );
O2A1O1Ixp5_ASAP7_75t_L g1705 ( .A1(n_1674), .A2(n_1607), .B(n_1578), .C(n_1642), .Y(n_1705) );
OR2x2_ASAP7_75t_L g1706 ( .A(n_1660), .B(n_1574), .Y(n_1706) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1673), .Y(n_1707) );
NOR2xp33_ASAP7_75t_L g1708 ( .A(n_1662), .B(n_1640), .Y(n_1708) );
INVx1_ASAP7_75t_SL g1709 ( .A(n_1652), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1710 ( .A(n_1675), .B(n_1629), .Y(n_1710) );
NAND2xp5_ASAP7_75t_L g1711 ( .A(n_1675), .B(n_1614), .Y(n_1711) );
AOI22xp5_ASAP7_75t_L g1712 ( .A1(n_1674), .A2(n_1587), .B1(n_1571), .B2(n_1584), .Y(n_1712) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1673), .Y(n_1713) );
O2A1O1Ixp33_ASAP7_75t_SL g1714 ( .A1(n_1678), .A2(n_1456), .B(n_1450), .C(n_1593), .Y(n_1714) );
OA21x2_ASAP7_75t_L g1715 ( .A1(n_1678), .A2(n_1600), .B(n_1597), .Y(n_1715) );
INVx1_ASAP7_75t_SL g1716 ( .A(n_1654), .Y(n_1716) );
OAI32xp33_ASAP7_75t_L g1717 ( .A1(n_1683), .A2(n_1608), .A3(n_1564), .B1(n_1561), .B2(n_1545), .Y(n_1717) );
INVx1_ASAP7_75t_SL g1718 ( .A(n_1654), .Y(n_1718) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1645), .Y(n_1719) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1646), .Y(n_1720) );
INVx2_ASAP7_75t_L g1721 ( .A(n_1665), .Y(n_1721) );
NOR3xp33_ASAP7_75t_L g1722 ( .A(n_1705), .B(n_1442), .C(n_1684), .Y(n_1722) );
AOI322xp5_ASAP7_75t_L g1723 ( .A1(n_1691), .A2(n_1664), .A3(n_1655), .B1(n_1671), .B2(n_1649), .C1(n_1685), .C2(n_1681), .Y(n_1723) );
NOR3xp33_ASAP7_75t_L g1724 ( .A(n_1705), .B(n_1684), .C(n_1671), .Y(n_1724) );
INVx2_ASAP7_75t_SL g1725 ( .A(n_1703), .Y(n_1725) );
INVx2_ASAP7_75t_L g1726 ( .A(n_1715), .Y(n_1726) );
INVxp67_ASAP7_75t_L g1727 ( .A(n_1709), .Y(n_1727) );
AOI221x1_ASAP7_75t_L g1728 ( .A1(n_1711), .A2(n_1689), .B1(n_1688), .B2(n_1647), .C(n_1656), .Y(n_1728) );
AOI211xp5_ASAP7_75t_L g1729 ( .A1(n_1702), .A2(n_1499), .B(n_1614), .C(n_1686), .Y(n_1729) );
NAND2xp5_ASAP7_75t_L g1730 ( .A(n_1695), .B(n_1658), .Y(n_1730) );
AOI21xp5_ASAP7_75t_L g1731 ( .A1(n_1702), .A2(n_1714), .B(n_1692), .Y(n_1731) );
OAI22xp33_ASAP7_75t_L g1732 ( .A1(n_1716), .A2(n_1663), .B1(n_1683), .B2(n_1679), .Y(n_1732) );
AOI221x1_ASAP7_75t_L g1733 ( .A1(n_1694), .A2(n_1407), .B1(n_1622), .B2(n_1623), .C(n_1603), .Y(n_1733) );
NOR3xp33_ASAP7_75t_L g1734 ( .A(n_1691), .B(n_1593), .C(n_1628), .Y(n_1734) );
AOI211xp5_ASAP7_75t_L g1735 ( .A1(n_1717), .A2(n_1571), .B(n_1612), .C(n_1628), .Y(n_1735) );
OAI221xp5_ASAP7_75t_SL g1736 ( .A1(n_1718), .A2(n_1663), .B1(n_1677), .B2(n_1672), .C(n_1666), .Y(n_1736) );
AOI22xp33_ASAP7_75t_L g1737 ( .A1(n_1704), .A2(n_1663), .B1(n_1638), .B2(n_1676), .Y(n_1737) );
NAND2xp5_ASAP7_75t_L g1738 ( .A(n_1698), .B(n_1651), .Y(n_1738) );
NOR3xp33_ASAP7_75t_L g1739 ( .A(n_1695), .B(n_1600), .C(n_1597), .Y(n_1739) );
AOI22xp5_ASAP7_75t_L g1740 ( .A1(n_1712), .A2(n_1669), .B1(n_1682), .B2(n_1668), .Y(n_1740) );
AOI21xp5_ASAP7_75t_L g1741 ( .A1(n_1715), .A2(n_1557), .B(n_1651), .Y(n_1741) );
AOI21xp5_ASAP7_75t_L g1742 ( .A1(n_1710), .A2(n_1557), .B(n_1630), .Y(n_1742) );
AOI221xp5_ASAP7_75t_L g1743 ( .A1(n_1693), .A2(n_1407), .B1(n_1606), .B2(n_1618), .C(n_1617), .Y(n_1743) );
NAND2xp33_ASAP7_75t_SL g1744 ( .A(n_1701), .B(n_1661), .Y(n_1744) );
AOI211xp5_ASAP7_75t_L g1745 ( .A1(n_1696), .A2(n_1458), .B(n_1450), .C(n_1545), .Y(n_1745) );
OAI21xp5_ASAP7_75t_SL g1746 ( .A1(n_1700), .A2(n_1561), .B(n_1545), .Y(n_1746) );
NAND3xp33_ASAP7_75t_L g1747 ( .A(n_1719), .B(n_1416), .C(n_1423), .Y(n_1747) );
AOI22xp5_ASAP7_75t_L g1748 ( .A1(n_1708), .A2(n_1637), .B1(n_1561), .B2(n_1531), .Y(n_1748) );
INVx2_ASAP7_75t_L g1749 ( .A(n_1707), .Y(n_1749) );
AOI221xp5_ASAP7_75t_L g1750 ( .A1(n_1720), .A2(n_1421), .B1(n_1420), .B2(n_1462), .C(n_1345), .Y(n_1750) );
NOR4xp75_ASAP7_75t_L g1751 ( .A(n_1699), .B(n_1281), .C(n_1445), .D(n_1555), .Y(n_1751) );
AOI22xp5_ASAP7_75t_L g1752 ( .A1(n_1721), .A2(n_1524), .B1(n_1506), .B2(n_1514), .Y(n_1752) );
O2A1O1Ixp5_ASAP7_75t_SL g1753 ( .A1(n_1713), .A2(n_1455), .B(n_1416), .C(n_1423), .Y(n_1753) );
NOR3xp33_ASAP7_75t_L g1754 ( .A(n_1697), .B(n_1445), .C(n_1440), .Y(n_1754) );
AOI22xp5_ASAP7_75t_L g1755 ( .A1(n_1706), .A2(n_1524), .B1(n_1506), .B2(n_1520), .Y(n_1755) );
OAI222xp33_ASAP7_75t_L g1756 ( .A1(n_1716), .A2(n_1475), .B1(n_1515), .B2(n_1514), .C1(n_1520), .C2(n_1428), .Y(n_1756) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1710), .Y(n_1757) );
AOI322xp5_ASAP7_75t_L g1758 ( .A1(n_1691), .A2(n_1429), .A3(n_1515), .B1(n_1559), .B2(n_1556), .C1(n_1555), .C2(n_1550), .Y(n_1758) );
OAI21xp5_ASAP7_75t_L g1759 ( .A1(n_1705), .A2(n_1472), .B(n_1475), .Y(n_1759) );
NOR2x1_ASAP7_75t_L g1760 ( .A(n_1731), .B(n_1732), .Y(n_1760) );
NAND3xp33_ASAP7_75t_SL g1761 ( .A(n_1724), .B(n_1735), .C(n_1729), .Y(n_1761) );
OAI321xp33_ASAP7_75t_L g1762 ( .A1(n_1736), .A2(n_1727), .A3(n_1759), .B1(n_1725), .B2(n_1737), .C(n_1743), .Y(n_1762) );
NAND3xp33_ASAP7_75t_SL g1763 ( .A(n_1722), .B(n_1723), .C(n_1751), .Y(n_1763) );
AOI221xp5_ASAP7_75t_L g1764 ( .A1(n_1734), .A2(n_1739), .B1(n_1757), .B2(n_1744), .C(n_1726), .Y(n_1764) );
NOR4xp25_ASAP7_75t_L g1765 ( .A(n_1730), .B(n_1746), .C(n_1756), .D(n_1747), .Y(n_1765) );
NOR2xp33_ASAP7_75t_L g1766 ( .A(n_1730), .B(n_1740), .Y(n_1766) );
NAND3xp33_ASAP7_75t_SL g1767 ( .A(n_1758), .B(n_1741), .C(n_1745), .Y(n_1767) );
NAND3xp33_ASAP7_75t_SL g1768 ( .A(n_1742), .B(n_1753), .C(n_1754), .Y(n_1768) );
O2A1O1Ixp33_ASAP7_75t_L g1769 ( .A1(n_1738), .A2(n_1749), .B(n_1750), .C(n_1728), .Y(n_1769) );
NAND2xp5_ASAP7_75t_SL g1770 ( .A(n_1748), .B(n_1755), .Y(n_1770) );
OR2x2_ASAP7_75t_L g1771 ( .A(n_1765), .B(n_1752), .Y(n_1771) );
AND3x2_ASAP7_75t_L g1772 ( .A(n_1764), .B(n_1733), .C(n_1475), .Y(n_1772) );
NAND5xp2_ASAP7_75t_L g1773 ( .A(n_1762), .B(n_1331), .C(n_1332), .D(n_1316), .E(n_1441), .Y(n_1773) );
INVx1_ASAP7_75t_L g1774 ( .A(n_1770), .Y(n_1774) );
NOR3x1_ASAP7_75t_L g1775 ( .A(n_1761), .B(n_1468), .C(n_1443), .Y(n_1775) );
NOR2x1_ASAP7_75t_L g1776 ( .A(n_1760), .B(n_1271), .Y(n_1776) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1769), .Y(n_1777) );
OR2x2_ASAP7_75t_L g1778 ( .A(n_1763), .B(n_1560), .Y(n_1778) );
NOR2x1p5_ASAP7_75t_L g1779 ( .A(n_1774), .B(n_1768), .Y(n_1779) );
BUFx2_ASAP7_75t_L g1780 ( .A(n_1778), .Y(n_1780) );
OR2x2_ASAP7_75t_L g1781 ( .A(n_1777), .B(n_1767), .Y(n_1781) );
HB1xp67_ASAP7_75t_L g1782 ( .A(n_1776), .Y(n_1782) );
INVx2_ASAP7_75t_L g1783 ( .A(n_1775), .Y(n_1783) );
AND2x2_ASAP7_75t_SL g1784 ( .A(n_1771), .B(n_1766), .Y(n_1784) );
INVx2_ASAP7_75t_L g1785 ( .A(n_1780), .Y(n_1785) );
INVx2_ASAP7_75t_L g1786 ( .A(n_1783), .Y(n_1786) );
INVx2_ASAP7_75t_L g1787 ( .A(n_1781), .Y(n_1787) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1784), .Y(n_1788) );
NOR2x1_ASAP7_75t_L g1789 ( .A(n_1779), .B(n_1773), .Y(n_1789) );
XNOR2x1_ASAP7_75t_L g1790 ( .A(n_1789), .B(n_1779), .Y(n_1790) );
NAND2xp5_ASAP7_75t_L g1791 ( .A(n_1786), .B(n_1772), .Y(n_1791) );
OAI22xp5_ASAP7_75t_L g1792 ( .A1(n_1785), .A2(n_1782), .B1(n_1560), .B2(n_1509), .Y(n_1792) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1787), .Y(n_1793) );
AOI222xp33_ASAP7_75t_L g1794 ( .A1(n_1793), .A2(n_1788), .B1(n_1321), .B2(n_1334), .C1(n_1432), .C2(n_1556), .Y(n_1794) );
OAI22xp5_ASAP7_75t_L g1795 ( .A1(n_1791), .A2(n_1432), .B1(n_1509), .B2(n_1464), .Y(n_1795) );
OA21x2_ASAP7_75t_L g1796 ( .A1(n_1790), .A2(n_1250), .B(n_1327), .Y(n_1796) );
AO221x2_ASAP7_75t_L g1797 ( .A1(n_1792), .A2(n_1494), .B1(n_1501), .B2(n_1488), .C(n_1487), .Y(n_1797) );
INVx1_ASAP7_75t_L g1798 ( .A(n_1795), .Y(n_1798) );
NAND3xp33_ASAP7_75t_SL g1799 ( .A(n_1794), .B(n_1250), .C(n_1559), .Y(n_1799) );
OAI21xp33_ASAP7_75t_L g1800 ( .A1(n_1797), .A2(n_1550), .B(n_1549), .Y(n_1800) );
OAI22xp33_ASAP7_75t_L g1801 ( .A1(n_1796), .A2(n_1464), .B1(n_1410), .B2(n_1494), .Y(n_1801) );
A2O1A1Ixp33_ASAP7_75t_L g1802 ( .A1(n_1798), .A2(n_1327), .B(n_1464), .C(n_1471), .Y(n_1802) );
OR2x2_ASAP7_75t_L g1803 ( .A(n_1799), .B(n_1568), .Y(n_1803) );
OAI21xp5_ASAP7_75t_L g1804 ( .A1(n_1801), .A2(n_1464), .B(n_1224), .Y(n_1804) );
OAI21xp5_ASAP7_75t_SL g1805 ( .A1(n_1800), .A2(n_1566), .B(n_1410), .Y(n_1805) );
OAI21xp33_ASAP7_75t_L g1806 ( .A1(n_1805), .A2(n_1566), .B(n_1568), .Y(n_1806) );
OAI22xp5_ASAP7_75t_L g1807 ( .A1(n_1803), .A2(n_1501), .B1(n_1487), .B2(n_1488), .Y(n_1807) );
OA21x2_ASAP7_75t_L g1808 ( .A1(n_1802), .A2(n_1804), .B(n_1245), .Y(n_1808) );
AOI22xp5_ASAP7_75t_L g1809 ( .A1(n_1806), .A2(n_1807), .B1(n_1808), .B2(n_1448), .Y(n_1809) );
endmodule