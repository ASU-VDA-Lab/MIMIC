module fake_jpeg_26573_n_49 (n_3, n_2, n_1, n_0, n_4, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_2),
.Y(n_6)
);

AND2x2_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_5),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_2),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_5),
.B(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_4),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_15),
.B(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_3),
.Y(n_18)
);

NAND3xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_21),
.C(n_22),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_14),
.B1(n_9),
.B2(n_13),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_10),
.B(n_7),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_27),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_12),
.C(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_23),
.B1(n_17),
.B2(n_7),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_29),
.B(n_24),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_26),
.B(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_17),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_42),
.C(n_30),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_12),
.B(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

OAI21x1_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_20),
.B(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_22),
.Y(n_46)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_20),
.CI(n_16),
.CON(n_48),
.SN(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_47),
.C(n_45),
.Y(n_49)
);


endmodule