module real_jpeg_29283_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_244;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_0),
.B(n_51),
.Y(n_83)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_0),
.B(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_0),
.B(n_213),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_29),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_45),
.B1(n_48),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_56),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_2),
.B(n_20),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_SL g179 ( 
.A1(n_2),
.A2(n_10),
.B(n_45),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_2),
.A2(n_50),
.B(n_52),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_2),
.B(n_62),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_4),
.A2(n_31),
.B1(n_45),
.B2(n_48),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_4),
.A2(n_31),
.B1(n_50),
.B2(n_51),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_6),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_115),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_6),
.A2(n_45),
.B1(n_48),
.B2(n_115),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_115),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_8),
.A2(n_45),
.B1(n_48),
.B2(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_131)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_10),
.Y(n_178)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_11),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_123),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_121),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_91),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_15),
.B(n_91),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_15),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_70),
.CI(n_78),
.CON(n_15),
.SN(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_38),
.B2(n_39),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_32),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_19),
.B(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_20),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_22),
.B(n_29),
.C(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_21),
.A2(n_34),
.B(n_36),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_21),
.B(n_114),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_23),
.B(n_26),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_24),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_24),
.B(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_24),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_24),
.A2(n_56),
.B(n_178),
.C(n_179),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_28),
.B(n_34),
.Y(n_257)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_33),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_35),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_36),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_37),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_40),
.B(n_136),
.C(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_40),
.A2(n_41),
.B1(n_138),
.B2(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_53),
.B(n_54),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_42),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_43),
.B(n_55),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_43),
.B(n_186),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_48),
.B1(n_60),
.B2(n_63),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_45),
.A2(n_47),
.B(n_56),
.C(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_49),
.B(n_186),
.Y(n_185)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_51),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_76),
.B(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_53),
.B(n_56),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_56),
.B(n_85),
.Y(n_228)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B(n_67),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_59),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_59),
.B(n_141),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_59),
.Y(n_260)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_62),
.B(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_68),
.B(n_151),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_71),
.B(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_72),
.B(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_72),
.A2(n_149),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_73),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_75),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_76),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B(n_90),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_80),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_82),
.B1(n_90),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_81),
.A2(n_82),
.B1(n_177),
.B2(n_180),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_82),
.B(n_177),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_86),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_83),
.B(n_86),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_83),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_84),
.Y(n_158)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_87),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_89),
.B(n_195),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_116),
.C(n_117),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_92),
.A2(n_93),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_107),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_94),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_102),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_95),
.B(n_102),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_96),
.B(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_97),
.A2(n_131),
.B(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_98),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_103),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_116),
.B(n_117),
.Y(n_281)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_277),
.B(n_282),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_264),
.B(n_276),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_171),
.B(n_246),
.C(n_263),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_159),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_127),
.B(n_159),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_142),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_129),
.B(n_135),
.C(n_142),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_130),
.B(n_133),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_132),
.B(n_212),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_134),
.B(n_185),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_137),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_144),
.B(n_147),
.C(n_152),
.Y(n_261)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_157),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_160),
.A2(n_161),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.C(n_169),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_245),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_238),
.B(n_244),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_197),
.B(n_237),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_187),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_175),
.B(n_187),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.C(n_183),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_176),
.B(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_177),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_235)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_194),
.C(n_196),
.Y(n_239)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_232),
.B(n_236),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_214),
.B(n_231),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_200),
.B(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_221),
.B(n_230),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_219),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_225),
.B(n_229),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_224),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_233),
.B(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_240),
.Y(n_244)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_247),
.B(n_248),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_261),
.B2(n_262),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_252),
.C(n_262),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_256),
.C(n_258),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_261),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_266),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_275),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_273),
.C(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);


endmodule