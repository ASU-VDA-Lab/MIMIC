module fake_jpeg_18725_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_14),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_16),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_19),
.B1(n_21),
.B2(n_18),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_35),
.B(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_21),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_24),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_21),
.B1(n_22),
.B2(n_14),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_27),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_17),
.C(n_27),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_32),
.B(n_35),
.C(n_31),
.Y(n_43)
);

AOI221xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_17),
.B1(n_11),
.B2(n_15),
.C(n_9),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_29),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_16),
.B1(n_8),
.B2(n_9),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_40),
.C(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_42),
.B(n_43),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_11),
.B(n_15),
.C(n_4),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_46),
.C(n_17),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B(n_5),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_6),
.B1(n_1),
.B2(n_3),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_3),
.Y(n_55)
);


endmodule