module real_jpeg_3242_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_321, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;
input n_321;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_0),
.A2(n_28),
.B1(n_31),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_0),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_0),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_0),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_136)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_3),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_3),
.A2(n_28),
.B1(n_31),
.B2(n_143),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_3),
.A2(n_38),
.B1(n_40),
.B2(n_143),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_143),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_4),
.A2(n_38),
.B1(n_40),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_4),
.A2(n_59),
.B1(n_65),
.B2(n_66),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_28),
.B1(n_31),
.B2(n_59),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_5),
.A2(n_28),
.B1(n_31),
.B2(n_68),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_5),
.A2(n_38),
.B1(n_40),
.B2(n_68),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_68),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_6),
.A2(n_30),
.B1(n_38),
.B2(n_40),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_30),
.B1(n_65),
.B2(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_6),
.A2(n_30),
.B1(n_50),
.B2(n_51),
.Y(n_161)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_11),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_11),
.A2(n_28),
.B1(n_31),
.B2(n_155),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_11),
.A2(n_38),
.B1(n_40),
.B2(n_155),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_155),
.Y(n_264)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_12),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_12),
.B(n_102),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_12),
.B(n_31),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_12),
.A2(n_65),
.B(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_12),
.B(n_49),
.C(n_51),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_12),
.A2(n_38),
.B1(n_40),
.B2(n_175),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_12),
.B(n_44),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_12),
.B(n_90),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_12),
.B(n_47),
.Y(n_265)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_12),
.A2(n_31),
.B(n_214),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_182),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_13),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_13),
.A2(n_28),
.B1(n_31),
.B2(n_182),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_13),
.A2(n_38),
.B1(n_40),
.B2(n_182),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_182),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_118),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_117),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_103),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.C(n_85),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_21),
.B(n_75),
.CI(n_85),
.CON(n_145),
.SN(n_145)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_60),
.B2(n_74),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_24),
.B(n_46),
.C(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_41),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_44),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_28),
.A2(n_31),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_28),
.A2(n_63),
.B(n_174),
.C(n_176),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_28),
.B(n_36),
.C(n_40),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_31),
.B(n_62),
.C(n_66),
.Y(n_176)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_32),
.A2(n_41),
.B(n_115),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_32),
.A2(n_113),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_32),
.A2(n_37),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_32),
.A2(n_37),
.B1(n_201),
.B2(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_34),
.A2(n_38),
.B(n_213),
.C(n_215),
.Y(n_212)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_37),
.A2(n_78),
.B(n_116),
.Y(n_140)
);

CKINVDCx6p67_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_40),
.B1(n_49),
.B2(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_38),
.B(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_42),
.B(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_44),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_44),
.A2(n_79),
.B1(n_179),
.B2(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_45),
.A2(n_46),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21x1_ASAP7_75t_R g46 ( 
.A1(n_47),
.A2(n_55),
.B(n_57),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_47),
.B(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_47),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_47),
.A2(n_55),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_47),
.A2(n_55),
.B1(n_247),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_58),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_48)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_51),
.B(n_259),
.Y(n_258)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_55),
.A2(n_81),
.B(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_58),
.A2(n_94),
.B(n_96),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_74),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_69),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_64),
.B1(n_72),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_61),
.A2(n_72),
.B1(n_142),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_61),
.A2(n_72),
.B1(n_154),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_61),
.A2(n_72),
.B1(n_181),
.B2(n_221),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_66),
.B(n_175),
.Y(n_174)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_99),
.B(n_101),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_72),
.A2(n_142),
.B(n_144),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_75),
.A2(n_76),
.B(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_83),
.A2(n_138),
.B(n_139),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_92),
.B(n_97),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_97),
.B1(n_98),
.B2(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_86),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_86),
.A2(n_93),
.B1(n_125),
.B2(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B(n_91),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_87),
.A2(n_160),
.B(n_162),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_87),
.A2(n_91),
.B(n_162),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_87),
.A2(n_89),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_88),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_88),
.A2(n_90),
.B1(n_161),
.B2(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_88),
.A2(n_133),
.B(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_88),
.A2(n_90),
.B1(n_175),
.B2(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_88),
.A2(n_90),
.B1(n_261),
.B2(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_91),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_89),
.A2(n_135),
.B(n_172),
.Y(n_207)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_90),
.B(n_136),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_93),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_95),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_94),
.A2(n_139),
.B1(n_210),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_102),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_146),
.B(n_317),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_145),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_121),
.B(n_145),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_127),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_126),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_127),
.A2(n_128),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_140),
.C(n_141),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_129),
.A2(n_130),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_132),
.B1(n_137),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_140),
.B(n_141),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_145),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_310),
.B(n_316),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_195),
.B(n_309),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_183),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_149),
.B(n_183),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_164),
.C(n_166),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_150),
.B(n_164),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_157),
.B2(n_158),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_156),
.C(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_159),
.B(n_163),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_166),
.B(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_177),
.C(n_180),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_167),
.A2(n_168),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_173),
.Y(n_235)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_177),
.B(n_180),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_194),
.Y(n_183)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_187),
.B(n_191),
.C(n_194),
.Y(n_315)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI321xp33_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_290),
.A3(n_301),
.B1(n_307),
.B2(n_308),
.C(n_321),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_236),
.B(n_289),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_217),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_198),
.B(n_217),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_208),
.C(n_211),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_199),
.B(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_204),
.C(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_208),
.B(n_211),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_212),
.B(n_216),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_229),
.B2(n_230),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_218),
.B(n_231),
.C(n_234),
.Y(n_302)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_220),
.B(n_224),
.C(n_228),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_284),
.B(n_288),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_274),
.B(n_283),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_255),
.B(n_273),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_248),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_252),
.C(n_254),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_250),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_267),
.B(n_272),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_262),
.B(n_266),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_265),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_279),
.C(n_281),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_287),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_293),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.C(n_300),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_295),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_303),
.Y(n_307)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_315),
.Y(n_316)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);


endmodule