module fake_jpeg_23371_n_324 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_15),
.B1(n_16),
.B2(n_22),
.Y(n_41)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_16),
.B1(n_34),
.B2(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_31),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_31),
.B1(n_38),
.B2(n_29),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_27),
.B1(n_24),
.B2(n_16),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_38),
.B1(n_30),
.B2(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_64),
.B1(n_70),
.B2(n_78),
.Y(n_80)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_65),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_39),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_30),
.Y(n_82)
);

AO22x2_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_29),
.B1(n_22),
.B2(n_13),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

CKINVDCx6p67_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_59),
.B1(n_58),
.B2(n_70),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_38),
.B(n_28),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_21),
.B(n_33),
.C(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_66),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_36),
.B1(n_30),
.B2(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_85),
.Y(n_106)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_59),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_50),
.B1(n_48),
.B2(n_42),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_96),
.B1(n_40),
.B2(n_74),
.Y(n_124)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_92),
.B1(n_40),
.B2(n_51),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_91),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_97),
.B1(n_101),
.B2(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_94),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_42),
.B1(n_36),
.B2(n_30),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_78),
.B(n_77),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_35),
.C(n_22),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_95),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_64),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_70),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_110),
.B(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_116),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_75),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_97),
.B1(n_79),
.B2(n_91),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_126),
.B(n_140),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_80),
.B1(n_83),
.B2(n_99),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_138),
.B1(n_112),
.B2(n_71),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_115),
.C(n_108),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_136),
.B1(n_137),
.B2(n_118),
.Y(n_168)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_114),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_104),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_135),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_88),
.B1(n_101),
.B2(n_63),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_63),
.B1(n_86),
.B2(n_89),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_95),
.B1(n_82),
.B2(n_36),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_146),
.B(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_13),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_163),
.C(n_32),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_114),
.B(n_103),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_152),
.A2(n_164),
.B(n_23),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_160),
.Y(n_183)
);

OAI22x1_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_109),
.B1(n_124),
.B2(n_22),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_158),
.B1(n_168),
.B2(n_170),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_155),
.B(n_161),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_145),
.B1(n_139),
.B2(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_159),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_125),
.B1(n_139),
.B2(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_131),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_13),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_176),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_119),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_111),
.B(n_13),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_146),
.B(n_130),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_169),
.A2(n_17),
.B(n_19),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_117),
.B1(n_62),
.B2(n_56),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_149),
.A2(n_86),
.B1(n_14),
.B2(n_13),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_173),
.B1(n_174),
.B2(n_68),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_62),
.B1(n_53),
.B2(n_100),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_53),
.B1(n_100),
.B2(n_86),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_76),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_32),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_159),
.B(n_81),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_180),
.B(n_198),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_33),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_185),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_33),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_33),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_28),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_192),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_17),
.C(n_19),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_102),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_89),
.Y(n_195)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_196),
.A2(n_175),
.B(n_170),
.Y(n_223)
);

OAI31xp33_ASAP7_75t_SL g197 ( 
.A1(n_154),
.A2(n_25),
.A3(n_21),
.B(n_26),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_202),
.B(n_164),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_55),
.C(n_54),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_32),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_156),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_25),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_200),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_167),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_204),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_184),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_207),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_215),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

AO22x1_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_158),
.B1(n_169),
.B2(n_172),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_18),
.B(n_1),
.Y(n_247)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_183),
.B(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_186),
.A2(n_165),
.B1(n_171),
.B2(n_14),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_224),
.A2(n_26),
.B1(n_55),
.B2(n_54),
.Y(n_231)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_190),
.B1(n_199),
.B2(n_179),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_230),
.B1(n_234),
.B2(n_242),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_202),
.CI(n_187),
.CON(n_228),
.SN(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_235),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_191),
.B1(n_189),
.B2(n_185),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_238),
.B1(n_222),
.B2(n_18),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_233),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_182),
.B1(n_183),
.B2(n_46),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_46),
.B1(n_43),
.B2(n_26),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_46),
.C(n_43),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_219),
.C(n_218),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_225),
.A2(n_211),
.B1(n_221),
.B2(n_206),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_43),
.B1(n_14),
.B2(n_21),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_32),
.B1(n_28),
.B2(n_26),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_243),
.C(n_244),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_208),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_254),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_208),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_257),
.Y(n_267)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_236),
.B(n_220),
.CI(n_209),
.CON(n_257),
.SN(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_212),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_265),
.Y(n_280)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_228),
.B(n_231),
.Y(n_277)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

XOR2x2_ASAP7_75t_SL g265 ( 
.A(n_228),
.B(n_0),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_232),
.B1(n_253),
.B2(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_275),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_239),
.B(n_247),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_265),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_251),
.A2(n_240),
.B1(n_229),
.B2(n_241),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_243),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_278),
.Y(n_286)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_245),
.C(n_2),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_1),
.C(n_2),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_289),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_273),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_285),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_267),
.B(n_257),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_293),
.C(n_281),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_250),
.B1(n_3),
.B2(n_4),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_18),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_286),
.B1(n_288),
.B2(n_290),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_2),
.C(n_3),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_18),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_18),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_296),
.B(n_11),
.Y(n_308)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_303),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_280),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_302),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_275),
.Y(n_302)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_6),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_3),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_4),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_310),
.B(n_7),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_311),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_7),
.B(n_8),
.Y(n_312)
);

A2O1A1O1Ixp25_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_295),
.B(n_302),
.C(n_300),
.D(n_10),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_316),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_300),
.B(n_301),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_307),
.B(n_308),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_315),
.C(n_9),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_8),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_317),
.B(n_9),
.Y(n_321)
);

AOI21x1_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_8),
.B(n_9),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_10),
.C(n_11),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_10),
.Y(n_324)
);


endmodule