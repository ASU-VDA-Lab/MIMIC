module fake_jpeg_30433_n_413 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_413);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_413;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_10),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_10),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_61),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_80),
.Y(n_108)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_83),
.Y(n_113)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_29),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_29),
.B1(n_43),
.B2(n_30),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_86),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_29),
.B1(n_43),
.B2(n_41),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_88),
.A2(n_112),
.B1(n_126),
.B2(n_83),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_84),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_95),
.B(n_39),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_42),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_115),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_133),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_29),
.B1(n_43),
.B2(n_32),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_39),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_73),
.A2(n_43),
.B1(n_41),
.B2(n_18),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_25),
.B1(n_37),
.B2(n_36),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_80),
.A2(n_57),
.B1(n_50),
.B2(n_53),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_48),
.A2(n_25),
.B1(n_37),
.B2(n_36),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_19),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_93),
.A2(n_58),
.B1(n_56),
.B2(n_68),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_155),
.B1(n_126),
.B2(n_86),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_145),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_19),
.B1(n_23),
.B2(n_18),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_153),
.Y(n_168)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_151),
.Y(n_188)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_149),
.Y(n_170)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_28),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_156),
.Y(n_182)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_32),
.B1(n_23),
.B2(n_28),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_158),
.Y(n_186)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_167),
.B(n_106),
.Y(n_171)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

OR2x2_ASAP7_75t_SL g179 ( 
.A(n_161),
.B(n_162),
.Y(n_179)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_111),
.A2(n_59),
.B1(n_82),
.B2(n_81),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_102),
.B1(n_98),
.B2(n_119),
.Y(n_172)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_107),
.B1(n_98),
.B2(n_109),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_146),
.B1(n_88),
.B2(n_112),
.Y(n_189)
);

AO22x1_ASAP7_75t_SL g187 ( 
.A1(n_153),
.A2(n_146),
.B1(n_87),
.B2(n_165),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_100),
.B1(n_110),
.B2(n_118),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_136),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_139),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_196),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_155),
.B(n_143),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_179),
.B(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_107),
.B1(n_87),
.B2(n_119),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_200),
.B1(n_202),
.B2(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_160),
.B(n_161),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_201),
.A2(n_113),
.B(n_177),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_109),
.B1(n_100),
.B2(n_110),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_188),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_208),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_227),
.B(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_179),
.C(n_183),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_217),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_224),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_173),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_194),
.B(n_92),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_220),
.Y(n_239)
);

AO21x2_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_187),
.B(n_173),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_218),
.B1(n_211),
.B2(n_215),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_207),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_211),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_231),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_238),
.B1(n_243),
.B2(n_247),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_214),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_196),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_210),
.C(n_212),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_203),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_245),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_200),
.B1(n_202),
.B2(n_206),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_223),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_246),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_189),
.B1(n_205),
.B2(n_206),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_192),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_244),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_195),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_200),
.B1(n_202),
.B2(n_206),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_233),
.A2(n_212),
.B(n_195),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_236),
.C(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_220),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_254),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_238),
.A2(n_205),
.B1(n_222),
.B2(n_213),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_265),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_222),
.B1(n_221),
.B2(n_206),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_266),
.B1(n_267),
.B2(n_226),
.Y(n_282)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_230),
.A2(n_221),
.B(n_206),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_222),
.B1(n_221),
.B2(n_198),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_221),
.B1(n_198),
.B2(n_226),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_235),
.B1(n_237),
.B2(n_231),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_268),
.A2(n_284),
.B1(n_288),
.B2(n_207),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_256),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_270),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_258),
.B(n_208),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_221),
.B1(n_240),
.B2(n_172),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_265),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_229),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_275),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g274 ( 
.A1(n_265),
.A2(n_227),
.B(n_241),
.C(n_229),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_170),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_242),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_289),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_227),
.B(n_223),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_260),
.B1(n_266),
.B2(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_225),
.Y(n_283)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_283),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_253),
.A2(n_234),
.B1(n_225),
.B2(n_228),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_170),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_178),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_204),
.Y(n_287)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_253),
.A2(n_224),
.B1(n_199),
.B2(n_197),
.Y(n_288)
);

BUFx12_ASAP7_75t_L g289 ( 
.A(n_257),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_248),
.B(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_255),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_295),
.B(n_305),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_297),
.A2(n_301),
.B1(n_284),
.B2(n_285),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_255),
.C(n_184),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_303),
.C(n_310),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_286),
.B1(n_278),
.B2(n_280),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_224),
.B1(n_207),
.B2(n_176),
.Y(n_302)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_184),
.C(n_183),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_289),
.B(n_224),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_288),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_307),
.B(n_289),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_178),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_313),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_180),
.C(n_174),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_178),
.Y(n_313)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_320),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_321),
.A2(n_322),
.B1(n_164),
.B2(n_134),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_293),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_323),
.B(n_325),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_296),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_331),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_293),
.B(n_274),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_272),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_334),
.Y(n_342)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_328),
.Y(n_345)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_309),
.Y(n_330)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_330),
.Y(n_354)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_332),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_274),
.B1(n_276),
.B2(n_176),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_335),
.Y(n_337)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_294),
.A2(n_274),
.B(n_162),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_180),
.C(n_174),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_14),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_316),
.A2(n_310),
.B1(n_300),
.B2(n_307),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_341),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_317),
.A2(n_300),
.B1(n_313),
.B2(n_292),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_351),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_325),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_349),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_319),
.A2(n_147),
.B1(n_166),
.B2(n_150),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_335),
.C(n_345),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_321),
.A2(n_137),
.B1(n_101),
.B2(n_159),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_163),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_352),
.Y(n_364)
);

XOR2x1_ASAP7_75t_L g353 ( 
.A(n_314),
.B(n_154),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_351),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_359),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_340),
.A2(n_314),
.B(n_318),
.Y(n_358)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_344),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_323),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_363),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_326),
.C(n_315),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_118),
.C(n_97),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_315),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_338),
.B(n_348),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_368),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_366),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_331),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_362),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_142),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_366),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_374),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_337),
.B(n_353),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_372),
.A2(n_124),
.B(n_43),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_355),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_346),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_359),
.B(n_354),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_375),
.B(n_379),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_364),
.B(n_129),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_380),
.B(n_367),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_382),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_355),
.C(n_81),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_386),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_9),
.C(n_17),
.Y(n_393)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_385),
.A2(n_378),
.B1(n_380),
.B2(n_377),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_370),
.B(n_11),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_12),
.Y(n_387)
);

AO21x1_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_389),
.B(n_391),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_376),
.A2(n_9),
.B(n_17),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_0),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_393),
.B(n_398),
.Y(n_400)
);

OAI321xp33_ASAP7_75t_L g396 ( 
.A1(n_388),
.A2(n_8),
.A3(n_17),
.B1(n_16),
.B2(n_15),
.C(n_13),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_396),
.A2(n_399),
.B(n_0),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_16),
.C(n_12),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_383),
.A2(n_16),
.B(n_12),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_395),
.B(n_390),
.C(n_8),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_402),
.C(n_403),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_33),
.C(n_1),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_404),
.B(n_396),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_0),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_400),
.A2(n_397),
.B(n_1),
.Y(n_407)
);

AOI322xp5_ASAP7_75t_L g409 ( 
.A1(n_407),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_33),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_408),
.B(n_409),
.Y(n_410)
);

OAI321xp33_ASAP7_75t_L g411 ( 
.A1(n_410),
.A2(n_405),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_1),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_411),
.B(n_4),
.Y(n_412)
);

AO21x1_ASAP7_75t_L g413 ( 
.A1(n_412),
.A2(n_4),
.B(n_33),
.Y(n_413)
);


endmodule