module fake_jpeg_27032_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_18),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_22),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_24),
.B1(n_26),
.B2(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_53),
.B1(n_54),
.B2(n_25),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_24),
.B1(n_26),
.B2(n_21),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_24),
.B1(n_26),
.B2(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_33),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_20),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_18),
.B(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_31),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_44),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_70),
.B(n_74),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_82),
.B1(n_88),
.B2(n_27),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_71),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_52),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_76),
.Y(n_102)
);

AO22x1_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_37),
.B1(n_38),
.B2(n_44),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_64),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_85),
.B(n_38),
.C(n_40),
.Y(n_110)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_86),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_45),
.B1(n_43),
.B2(n_20),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_25),
.B1(n_49),
.B2(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_45),
.B1(n_37),
.B2(n_30),
.Y(n_82)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_89),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_44),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_57),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_32),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_49),
.B1(n_55),
.B2(n_62),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_92),
.B1(n_97),
.B2(n_19),
.Y(n_134)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_47),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_103),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_32),
.B1(n_27),
.B2(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_67),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_108),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_77),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_68),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_22),
.B(n_19),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_112),
.B(n_113),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2x1p5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_85),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_112),
.B(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_129),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_132),
.Y(n_138)
);

AO22x1_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_82),
.B1(n_84),
.B2(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_86),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_101),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_87),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_134),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_87),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_80),
.B1(n_76),
.B2(n_38),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_98),
.B1(n_105),
.B2(n_109),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_150),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_143),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_99),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_152),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_100),
.B1(n_122),
.B2(n_108),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_127),
.B1(n_135),
.B2(n_98),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_119),
.B1(n_115),
.B2(n_96),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_101),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_123),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_11),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C1(n_5),
.C2(n_6),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_155),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_131),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_159),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_114),
.Y(n_161)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_135),
.C(n_118),
.Y(n_163)
);

AOI321xp33_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_164),
.A3(n_52),
.B1(n_19),
.B2(n_66),
.C(n_50),
.Y(n_186)
);

XOR2x2_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_128),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_167),
.A2(n_141),
.B1(n_151),
.B2(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_14),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_172),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_152),
.B1(n_141),
.B2(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_127),
.B1(n_142),
.B2(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_136),
.B1(n_144),
.B2(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_139),
.B(n_147),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_182),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_1),
.B(n_2),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_169),
.B(n_162),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_158),
.B(n_2),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_159),
.C(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_189),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_173),
.C(n_166),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_173),
.C(n_166),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_194),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_66),
.C(n_50),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_175),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_180),
.B1(n_187),
.B2(n_184),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_201),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_197),
.A2(n_176),
.B(n_183),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_205),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_174),
.B(n_186),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_206),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_50),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_200),
.C(n_205),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_188),
.C(n_190),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_191),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_212),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_192),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_1),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_218),
.B(n_4),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_211),
.A2(n_210),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_217),
.A2(n_3),
.B(n_4),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_2),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_216),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_6),
.C(n_8),
.Y(n_223)
);

AOI21x1_ASAP7_75t_SL g222 ( 
.A1(n_220),
.A2(n_221),
.B(n_5),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

AOI221xp5_ASAP7_75t_SL g225 ( 
.A1(n_224),
.A2(n_223),
.B1(n_9),
.B2(n_10),
.C(n_6),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_9),
.Y(n_226)
);


endmodule