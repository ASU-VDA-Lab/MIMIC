module fake_jpeg_2834_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_11),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_60),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx12_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_64),
.Y(n_81)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_43),
.B1(n_39),
.B2(n_49),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_38),
.B1(n_39),
.B2(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_58),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_56),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_77),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_53),
.Y(n_77)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_47),
.B(n_53),
.C(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_42),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_41),
.C(n_40),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_89),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_44),
.C(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_62),
.B1(n_69),
.B2(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_111),
.Y(n_119)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_16),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_25),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_83),
.B1(n_52),
.B2(n_2),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_52),
.B(n_1),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_116),
.B(n_118),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_0),
.C(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_114),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_3),
.Y(n_114)
);

OR2x2_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_4),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_88),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_126),
.B1(n_14),
.B2(n_18),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_89),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_131),
.C(n_21),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_8),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_10),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_12),
.C(n_13),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_23),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_116),
.B1(n_106),
.B2(n_26),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_137),
.B(n_27),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_141),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_128),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_142),
.A2(n_131),
.B(n_132),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_SL g147 ( 
.A(n_144),
.B(n_146),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_133),
.B1(n_138),
.B2(n_124),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_147),
.A2(n_145),
.B(n_143),
.Y(n_148)
);

OAI221xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_139),
.B1(n_124),
.B2(n_129),
.C(n_125),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_134),
.C(n_139),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_29),
.C(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_34),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_35),
.B(n_36),
.Y(n_153)
);


endmodule