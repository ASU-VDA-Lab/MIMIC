module fake_jpeg_31693_n_185 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_19),
.B(n_36),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_25),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_81),
.Y(n_91)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_85),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_54),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_72),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_75),
.B1(n_73),
.B2(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_100),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_86),
.A2(n_71),
.B1(n_75),
.B2(n_68),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_73),
.B1(n_60),
.B2(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_77),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_101),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_71),
.B1(n_68),
.B2(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_59),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_68),
.CON(n_102),
.SN(n_102)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_62),
.B(n_74),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_92),
.B1(n_88),
.B2(n_94),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_132)
);

INVx5_ASAP7_75t_SL g104 ( 
.A(n_91),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_2),
.Y(n_128)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_62),
.C(n_60),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_64),
.C(n_61),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_111),
.Y(n_133)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_78),
.B1(n_67),
.B2(n_66),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_116),
.B1(n_53),
.B2(n_49),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_58),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_122),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_55),
.B1(n_18),
.B2(n_21),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_117),
.Y(n_142)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_95),
.B(n_17),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_8),
.Y(n_140)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_1),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_24),
.A3(n_52),
.B1(n_51),
.B2(n_50),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_128),
.B(n_141),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_4),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_136),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_104),
.B1(n_117),
.B2(n_16),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_48),
.A3(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_7),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_13),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_8),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_9),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_9),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_14),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_148),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_150),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_152),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_154),
.B1(n_163),
.B2(n_125),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_30),
.B(n_32),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_155),
.A2(n_159),
.B(n_158),
.Y(n_167)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_15),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_15),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_128),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_142),
.B1(n_144),
.B2(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_170),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_148),
.A2(n_133),
.B(n_127),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_172),
.C(n_147),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_175),
.B(n_149),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_147),
.C(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

AOI321xp33_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_178),
.A3(n_149),
.B1(n_162),
.B2(n_156),
.C(n_170),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_173),
.C(n_165),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_166),
.C(n_171),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_33),
.B(n_38),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_39),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_146),
.Y(n_185)
);


endmodule