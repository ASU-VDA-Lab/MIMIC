module fake_netlist_1_2752_n_49 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_49);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_49;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_48;
wire n_46;
wire n_30;
wire n_25;
wire n_26;
wire n_33;
wire n_16;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_8), .B(n_6), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_0), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_3), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_4), .Y(n_22) );
INVx3_ASAP7_75t_L g23 ( .A(n_5), .Y(n_23) );
NOR2xp33_ASAP7_75t_SL g24 ( .A(n_14), .B(n_15), .Y(n_24) );
INVx1_ASAP7_75t_SL g25 ( .A(n_18), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
BUFx3_ASAP7_75t_L g28 ( .A(n_17), .Y(n_28) );
BUFx3_ASAP7_75t_L g29 ( .A(n_17), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_26), .B(n_20), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_28), .B(n_20), .Y(n_32) );
NOR2xp33_ASAP7_75t_SL g33 ( .A(n_30), .B(n_25), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
NAND2xp5_ASAP7_75t_SL g35 ( .A(n_33), .B(n_32), .Y(n_35) );
OR2x2_ASAP7_75t_L g36 ( .A(n_34), .B(n_18), .Y(n_36) );
NAND4xp25_ASAP7_75t_L g37 ( .A(n_36), .B(n_22), .C(n_23), .D(n_16), .Y(n_37) );
OAI21xp33_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_29), .B(n_28), .Y(n_38) );
OAI21xp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_29), .B(n_28), .Y(n_39) );
AOI22xp33_ASAP7_75t_L g40 ( .A1(n_37), .A2(n_29), .B1(n_17), .B2(n_27), .Y(n_40) );
NOR2xp33_ASAP7_75t_SL g41 ( .A(n_39), .B(n_24), .Y(n_41) );
INVx1_ASAP7_75t_SL g42 ( .A(n_38), .Y(n_42) );
OAI22xp5_ASAP7_75t_L g43 ( .A1(n_40), .A2(n_16), .B1(n_21), .B2(n_19), .Y(n_43) );
OR5x1_ASAP7_75t_L g44 ( .A(n_41), .B(n_0), .C(n_1), .D(n_2), .E(n_3), .Y(n_44) );
XOR2x1_ASAP7_75t_L g45 ( .A(n_41), .B(n_1), .Y(n_45) );
AO22x2_ASAP7_75t_L g46 ( .A1(n_44), .A2(n_42), .B1(n_4), .B2(n_5), .Y(n_46) );
INVx1_ASAP7_75t_SL g47 ( .A(n_45), .Y(n_47) );
OAI22xp5_ASAP7_75t_SL g48 ( .A1(n_47), .A2(n_43), .B1(n_2), .B2(n_10), .Y(n_48) );
AOI22xp5_ASAP7_75t_L g49 ( .A1(n_48), .A2(n_46), .B1(n_9), .B2(n_11), .Y(n_49) );
endmodule