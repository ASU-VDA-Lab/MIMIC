module fake_aes_10040_n_581 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_581);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_581;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_70;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g70 ( .A(n_27), .Y(n_70) );
CKINVDCx5p33_ASAP7_75t_R g71 ( .A(n_9), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_62), .Y(n_72) );
CKINVDCx5p33_ASAP7_75t_R g73 ( .A(n_57), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_47), .Y(n_74) );
CKINVDCx20_ASAP7_75t_R g75 ( .A(n_59), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_43), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_56), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_1), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_0), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_15), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_8), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_48), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_4), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_17), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_64), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_26), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_54), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_31), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_24), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_12), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_45), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_1), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_23), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_46), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_63), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_20), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_12), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_30), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_66), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_7), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_11), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_61), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_37), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_0), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_51), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_41), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_52), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_7), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_21), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_29), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_3), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_80), .Y(n_113) );
OR2x6_ASAP7_75t_L g114 ( .A(n_80), .B(n_32), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_75), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_89), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_83), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_106), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_83), .B(n_2), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_83), .B(n_2), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_107), .Y(n_122) );
NAND2xp33_ASAP7_75t_SL g123 ( .A(n_71), .B(n_3), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_90), .Y(n_124) );
XOR2xp5_ASAP7_75t_L g125 ( .A(n_112), .B(n_4), .Y(n_125) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_70), .A2(n_34), .B(n_68), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_70), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_72), .Y(n_129) );
NOR2xp33_ASAP7_75t_R g130 ( .A(n_73), .B(n_33), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_74), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_74), .A2(n_28), .B(n_67), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_104), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_105), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_77), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_77), .Y(n_139) );
INVxp33_ASAP7_75t_L g140 ( .A(n_79), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_99), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_86), .Y(n_144) );
NOR2xp67_ASAP7_75t_L g145 ( .A(n_92), .B(n_5), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_99), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_91), .B(n_5), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_109), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_127), .A2(n_95), .B(n_87), .C(n_88), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_118), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_118), .B(n_97), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_126), .Y(n_153) );
BUFx4f_ASAP7_75t_L g154 ( .A(n_114), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_120), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_132), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_140), .B(n_95), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_132), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_126), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
OR2x2_ASAP7_75t_SL g163 ( .A(n_116), .B(n_97), .Y(n_163) );
NAND2x1p5_ASAP7_75t_L g164 ( .A(n_120), .B(n_94), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_118), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_140), .B(n_94), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_134), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_115), .B(n_98), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_148), .B(n_98), .Y(n_170) );
OAI221xp5_ASAP7_75t_L g171 ( .A1(n_142), .A2(n_84), .B1(n_110), .B2(n_81), .C(n_101), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_116), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_124), .A2(n_84), .B1(n_110), .B2(n_81), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_136), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_136), .Y(n_175) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_137), .Y(n_176) );
AND2x6_ASAP7_75t_L g177 ( .A(n_148), .B(n_100), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_120), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_120), .Y(n_180) );
BUFx4f_ASAP7_75t_L g181 ( .A(n_114), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_120), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_131), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_121), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_115), .B(n_111), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_121), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
OAI221xp5_ASAP7_75t_L g188 ( .A1(n_142), .A2(n_102), .B1(n_101), .B2(n_93), .C(n_78), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_121), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_148), .B(n_102), .Y(n_190) );
AO22x2_ASAP7_75t_L g191 ( .A1(n_148), .A2(n_87), .B1(n_88), .B2(n_100), .Y(n_191) );
AO22x2_ASAP7_75t_L g192 ( .A1(n_148), .A2(n_121), .B1(n_125), .B2(n_146), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_121), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_114), .A2(n_103), .B1(n_96), .B2(n_85), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_157), .B(n_128), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_166), .B(n_128), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_151), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_151), .Y(n_201) );
INVx8_ASAP7_75t_L g202 ( .A(n_177), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_151), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_154), .B(n_130), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_187), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_154), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_158), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_165), .B(n_129), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_152), .B(n_114), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_165), .B(n_152), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_155), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_187), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_176), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_154), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_152), .B(n_114), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_178), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_177), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_183), .Y(n_221) );
NOR2xp33_ASAP7_75t_R g222 ( .A(n_172), .B(n_117), .Y(n_222) );
INVx2_ASAP7_75t_SL g223 ( .A(n_154), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_152), .B(n_129), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_185), .B(n_139), .Y(n_225) );
NOR3xp33_ASAP7_75t_SL g226 ( .A(n_188), .B(n_119), .C(n_122), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_178), .Y(n_227) );
NAND2xp33_ASAP7_75t_SL g228 ( .A(n_194), .B(n_130), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_168), .B(n_114), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_178), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_168), .B(n_139), .Y(n_231) );
BUFx12f_ASAP7_75t_L g232 ( .A(n_163), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_170), .B(n_145), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_170), .B(n_143), .Y(n_234) );
NOR2xp33_ASAP7_75t_R g235 ( .A(n_181), .B(n_123), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_181), .A2(n_143), .B1(n_127), .B2(n_138), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_170), .B(n_144), .Y(n_237) );
NOR2xp33_ASAP7_75t_R g238 ( .A(n_181), .B(n_178), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_186), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_192), .Y(n_240) );
BUFx10_ASAP7_75t_L g241 ( .A(n_177), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_186), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_170), .B(n_145), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_186), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_183), .Y(n_245) );
NAND3xp33_ASAP7_75t_L g246 ( .A(n_173), .B(n_123), .C(n_144), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_202), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_211), .B(n_190), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_231), .B(n_177), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_239), .Y(n_250) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_211), .B(n_181), .Y(n_251) );
OR2x6_ASAP7_75t_L g252 ( .A(n_202), .B(n_192), .Y(n_252) );
NOR2xp33_ASAP7_75t_SL g253 ( .A(n_214), .B(n_177), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_204), .A2(n_150), .B(n_138), .C(n_133), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_239), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_211), .A2(n_191), .B1(n_177), .B2(n_192), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_239), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_224), .B(n_177), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_234), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_202), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_205), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_225), .A2(n_180), .B(n_182), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_202), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_237), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_229), .B(n_177), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_197), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_229), .B(n_212), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_220), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_198), .A2(n_193), .B(n_186), .C(n_189), .Y(n_270) );
OR2x2_ASAP7_75t_L g271 ( .A(n_214), .B(n_125), .Y(n_271) );
OAI21xp33_ASAP7_75t_L g272 ( .A1(n_199), .A2(n_192), .B(n_191), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_215), .B(n_191), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_209), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_195), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_211), .A2(n_191), .B1(n_164), .B2(n_190), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_209), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_218), .B(n_190), .Y(n_278) );
INVxp67_ASAP7_75t_SL g279 ( .A(n_218), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_218), .A2(n_190), .B1(n_193), .B2(n_189), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_213), .A2(n_180), .B(n_184), .Y(n_281) );
NOR2xp33_ASAP7_75t_SL g282 ( .A(n_217), .B(n_164), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_218), .B(n_163), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_195), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_246), .B(n_171), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_220), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_241), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_210), .B(n_164), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_200), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_259), .B(n_264), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_272), .A2(n_240), .B1(n_228), .B2(n_203), .Y(n_291) );
OA21x2_ASAP7_75t_L g292 ( .A1(n_270), .A2(n_256), .B(n_281), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_256), .A2(n_217), .B1(n_203), .B2(n_200), .Y(n_293) );
NAND3xp33_ASAP7_75t_SL g294 ( .A(n_276), .B(n_235), .C(n_201), .Y(n_294) );
NOR2xp33_ASAP7_75t_R g295 ( .A(n_261), .B(n_232), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_247), .Y(n_296) );
OAI22xp33_ASAP7_75t_L g297 ( .A1(n_252), .A2(n_217), .B1(n_201), .B2(n_232), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_266), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_248), .B(n_213), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_252), .A2(n_233), .B1(n_243), .B2(n_193), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_252), .A2(n_233), .B1(n_243), .B2(n_193), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_251), .A2(n_182), .B1(n_184), .B2(n_236), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_248), .B(n_206), .Y(n_303) );
NOR2x1p5_ASAP7_75t_L g304 ( .A(n_261), .B(n_207), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_248), .A2(n_233), .B1(n_243), .B2(n_206), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_278), .B(n_223), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_275), .Y(n_307) );
BUFx3_ASAP7_75t_L g308 ( .A(n_247), .Y(n_308) );
O2A1O1Ixp5_ASAP7_75t_L g309 ( .A1(n_270), .A2(n_141), .B(n_147), .C(n_233), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_267), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_285), .A2(n_227), .B1(n_244), .B2(n_242), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_247), .Y(n_312) );
NAND2x1_ASAP7_75t_L g313 ( .A(n_275), .B(n_216), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g314 ( .A1(n_282), .A2(n_207), .B1(n_223), .B2(n_133), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_262), .A2(n_135), .B(n_126), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_278), .A2(n_207), .B1(n_244), .B2(n_242), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_278), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_290), .B(n_289), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_290), .B(n_279), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_293), .A2(n_288), .B1(n_251), .B2(n_280), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_309), .A2(n_249), .B(n_258), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_307), .B(n_273), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_294), .A2(n_283), .B1(n_222), .B2(n_268), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_298), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_297), .A2(n_226), .B1(n_283), .B2(n_254), .C(n_271), .Y(n_325) );
AOI21xp33_ASAP7_75t_L g326 ( .A1(n_297), .A2(n_253), .B(n_265), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_294), .A2(n_280), .B1(n_207), .B2(n_274), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_307), .B(n_284), .Y(n_328) );
NAND2x1_ASAP7_75t_L g329 ( .A(n_307), .B(n_312), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_293), .A2(n_207), .B1(n_284), .B2(n_156), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_291), .A2(n_277), .B1(n_260), .B2(n_247), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_300), .A2(n_238), .B1(n_255), .B2(n_250), .Y(n_332) );
AOI22xp33_ASAP7_75t_SL g333 ( .A1(n_295), .A2(n_131), .B1(n_146), .B2(n_126), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_302), .A2(n_254), .B1(n_219), .B2(n_227), .C(n_230), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_300), .A2(n_257), .B1(n_230), .B2(n_216), .Y(n_335) );
OAI221xp5_ASAP7_75t_L g336 ( .A1(n_301), .A2(n_219), .B1(n_169), .B2(n_167), .C(n_156), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_309), .B(n_147), .C(n_141), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_301), .A2(n_260), .B1(n_263), .B2(n_269), .Y(n_338) );
INVx4_ASAP7_75t_L g339 ( .A(n_312), .Y(n_339) );
AO21x2_ASAP7_75t_L g340 ( .A1(n_315), .A2(n_147), .B(n_141), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_298), .B(n_208), .Y(n_341) );
OAI31xp33_ASAP7_75t_L g342 ( .A1(n_320), .A2(n_304), .A3(n_302), .B(n_314), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_318), .Y(n_343) );
OAI21x1_ASAP7_75t_L g344 ( .A1(n_329), .A2(n_315), .B(n_313), .Y(n_344) );
NAND4xp25_ASAP7_75t_SL g345 ( .A(n_325), .B(n_291), .C(n_305), .D(n_304), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_319), .B(n_292), .Y(n_346) );
OAI211xp5_ASAP7_75t_SL g347 ( .A1(n_323), .A2(n_103), .B(n_310), .C(n_311), .Y(n_347) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_337), .A2(n_315), .B(n_311), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_324), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_330), .A2(n_314), .B1(n_292), .B2(n_310), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_330), .A2(n_317), .B1(n_292), .B2(n_303), .Y(n_351) );
NOR3xp33_ASAP7_75t_SL g352 ( .A(n_324), .B(n_76), .C(n_82), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_328), .Y(n_353) );
NAND2xp33_ASAP7_75t_SL g354 ( .A(n_318), .B(n_312), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_328), .Y(n_355) );
NAND3xp33_ASAP7_75t_L g356 ( .A(n_333), .B(n_292), .C(n_313), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_322), .B(n_292), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_340), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_327), .A2(n_317), .B1(n_299), .B2(n_303), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_322), .B(n_299), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g361 ( .A1(n_326), .A2(n_306), .B1(n_308), .B2(n_296), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_340), .Y(n_363) );
OAI31xp33_ASAP7_75t_L g364 ( .A1(n_331), .A2(n_306), .A3(n_159), .B(n_179), .Y(n_364) );
OAI33xp33_ASAP7_75t_L g365 ( .A1(n_341), .A2(n_113), .A3(n_167), .B1(n_159), .B2(n_175), .B3(n_162), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_339), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_334), .B(n_306), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_339), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_339), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_358), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_346), .B(n_339), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_349), .B(n_335), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_358), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_346), .B(n_126), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_369), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_349), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_343), .B(n_332), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_357), .B(n_135), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_347), .A2(n_321), .B1(n_337), .B2(n_338), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_358), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_357), .B(n_135), .Y(n_382) );
OAI31xp33_ASAP7_75t_L g383 ( .A1(n_345), .A2(n_336), .A3(n_131), .B(n_146), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_362), .B(n_135), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_343), .A2(n_359), .B1(n_350), .B2(n_356), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_353), .B(n_321), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_362), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_363), .B(n_135), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_363), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_363), .B(n_131), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_369), .B(n_146), .Y(n_392) );
INVx4_ASAP7_75t_L g393 ( .A(n_369), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_367), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_367), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_364), .A2(n_316), .B1(n_146), .B2(n_179), .C(n_169), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_353), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_370), .Y(n_399) );
OAI211xp5_ASAP7_75t_L g400 ( .A1(n_342), .A2(n_162), .B(n_175), .C(n_113), .Y(n_400) );
AND2x4_ASAP7_75t_SL g401 ( .A(n_370), .B(n_312), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_370), .B(n_153), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_355), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_366), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_354), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_351), .B(n_153), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_348), .B(n_153), .Y(n_409) );
NAND4xp25_ASAP7_75t_L g410 ( .A(n_342), .B(n_160), .C(n_174), .D(n_9), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_344), .Y(n_411) );
AOI211xp5_ASAP7_75t_L g412 ( .A1(n_359), .A2(n_108), .B(n_174), .C(n_160), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g413 ( .A1(n_350), .A2(n_308), .B1(n_296), .B2(n_312), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_344), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_377), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_410), .A2(n_365), .B1(n_352), .B2(n_368), .C(n_361), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_410), .A2(n_360), .B1(n_356), .B2(n_348), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_372), .B(n_348), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_398), .B(n_360), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_398), .B(n_348), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_378), .B(n_6), .Y(n_421) );
OAI33xp33_ASAP7_75t_L g422 ( .A1(n_402), .A2(n_6), .A3(n_8), .B1(n_10), .B2(n_11), .B3(n_13), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_371), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_394), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_402), .B(n_13), .Y(n_425) );
NAND2xp33_ASAP7_75t_R g426 ( .A(n_372), .B(n_14), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_394), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_372), .B(n_14), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_404), .B(n_15), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_399), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_404), .B(n_16), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_378), .B(n_16), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_395), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_393), .B(n_308), .Y(n_434) );
NAND2xp33_ASAP7_75t_SL g435 ( .A(n_393), .B(n_312), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_395), .B(n_17), .Y(n_436) );
NOR2xp33_ASAP7_75t_SL g437 ( .A(n_393), .B(n_296), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_376), .B(n_18), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_399), .Y(n_439) );
NAND5xp2_ASAP7_75t_L g440 ( .A(n_412), .B(n_19), .C(n_20), .D(n_21), .E(n_22), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_373), .B(n_19), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_373), .B(n_161), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_376), .B(n_312), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_371), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_399), .B(n_208), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_387), .B(n_161), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_393), .B(n_263), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_407), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_412), .B(n_196), .C(n_35), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_393), .B(n_399), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_387), .B(n_161), .Y(n_452) );
INVxp67_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
NOR2x1p5_ASAP7_75t_L g454 ( .A(n_405), .B(n_161), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_405), .B(n_161), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_375), .B(n_161), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_381), .B(n_384), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_405), .B(n_153), .Y(n_458) );
NAND4xp25_ASAP7_75t_L g459 ( .A(n_386), .B(n_183), .C(n_196), .D(n_221), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_371), .Y(n_460) );
AND3x1_ASAP7_75t_L g461 ( .A(n_383), .B(n_25), .C(n_36), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_375), .B(n_153), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_392), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_415), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_432), .B(n_397), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_457), .B(n_381), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_417), .A2(n_386), .B1(n_413), .B2(n_397), .Y(n_467) );
AOI32xp33_ASAP7_75t_L g468 ( .A1(n_461), .A2(n_406), .A3(n_413), .B1(n_392), .B2(n_414), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_454), .A2(n_380), .B1(n_384), .B2(n_388), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_421), .A2(n_383), .B1(n_400), .B2(n_405), .C(n_375), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_428), .B(n_401), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_424), .B(n_388), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_427), .B(n_371), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_428), .B(n_401), .Y(n_474) );
OAI211xp5_ASAP7_75t_L g475 ( .A1(n_421), .A2(n_416), .B(n_459), .C(n_436), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_419), .B(n_374), .Y(n_476) );
AOI222xp33_ASAP7_75t_L g477 ( .A1(n_422), .A2(n_408), .B1(n_400), .B2(n_379), .C1(n_382), .C2(n_391), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_463), .B(n_374), .Y(n_478) );
NAND3x2_ASAP7_75t_L g479 ( .A(n_431), .B(n_408), .C(n_391), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_418), .B(n_374), .Y(n_480) );
NAND3xp33_ASAP7_75t_SL g481 ( .A(n_436), .B(n_380), .C(n_391), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_440), .B(n_414), .C(n_379), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_433), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_447), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_453), .B(n_408), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_441), .B(n_401), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_426), .A2(n_414), .B1(n_396), .B2(n_401), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_425), .A2(n_396), .B(n_379), .C(n_382), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_426), .A2(n_396), .B1(n_390), .B2(n_411), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_451), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_418), .B(n_390), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_449), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_420), .B(n_390), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_451), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_423), .B(n_382), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_438), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_423), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_429), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_444), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_439), .B(n_409), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_439), .A2(n_403), .B1(n_411), .B2(n_409), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_444), .Y(n_502) );
NAND4xp25_ASAP7_75t_SL g503 ( .A(n_430), .B(n_411), .C(n_403), .D(n_389), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_460), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_460), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_434), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_455), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_434), .B(n_38), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_464), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_468), .B(n_435), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_498), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_489), .B(n_435), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_496), .B(n_442), .Y(n_513) );
NOR2xp33_ASAP7_75t_R g514 ( .A(n_503), .B(n_450), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_483), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_484), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_475), .A2(n_437), .B1(n_448), .B2(n_456), .C(n_462), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_492), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_467), .A2(n_445), .B(n_452), .C(n_446), .Y(n_519) );
OAI211xp5_ASAP7_75t_L g520 ( .A1(n_479), .A2(n_443), .B(n_403), .C(n_458), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_490), .B(n_434), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_467), .B(n_458), .C(n_455), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_466), .Y(n_523) );
NOR3xp33_ASAP7_75t_SL g524 ( .A(n_481), .B(n_39), .C(n_40), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_494), .B(n_389), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_476), .Y(n_526) );
NAND3xp33_ASAP7_75t_SL g527 ( .A(n_487), .B(n_385), .C(n_44), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_480), .B(n_491), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_488), .B(n_385), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_470), .A2(n_385), .B(n_153), .C(n_269), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_495), .B(n_42), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_482), .A2(n_286), .B1(n_269), .B2(n_287), .Y(n_532) );
NOR3xp33_ASAP7_75t_SL g533 ( .A(n_465), .B(n_49), .C(n_50), .Y(n_533) );
NOR3xp33_ASAP7_75t_L g534 ( .A(n_469), .B(n_245), .C(n_221), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_472), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_472), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_473), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_473), .Y(n_538) );
OAI211xp5_ASAP7_75t_L g539 ( .A1(n_510), .A2(n_477), .B(n_486), .C(n_506), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_537), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_511), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_528), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_538), .Y(n_543) );
XNOR2xp5_ASAP7_75t_L g544 ( .A(n_522), .B(n_510), .Y(n_544) );
OAI31xp33_ASAP7_75t_L g545 ( .A1(n_520), .A2(n_469), .A3(n_501), .B(n_471), .Y(n_545) );
OAI211xp5_ASAP7_75t_L g546 ( .A1(n_519), .A2(n_508), .B(n_474), .C(n_485), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_509), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_514), .A2(n_501), .B1(n_507), .B2(n_500), .Y(n_548) );
OAI211xp5_ASAP7_75t_SL g549 ( .A1(n_512), .A2(n_495), .B(n_493), .C(n_478), .Y(n_549) );
OAI311xp33_ASAP7_75t_L g550 ( .A1(n_530), .A2(n_504), .A3(n_499), .B1(n_502), .C1(n_505), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_535), .B(n_497), .Y(n_551) );
XNOR2x1_ASAP7_75t_L g552 ( .A(n_523), .B(n_53), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_512), .A2(n_286), .B(n_269), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_521), .B(n_55), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_526), .B(n_58), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_536), .B(n_60), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_515), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_543), .B(n_529), .Y(n_558) );
NAND4xp75_ASAP7_75t_L g559 ( .A(n_545), .B(n_524), .C(n_533), .D(n_513), .Y(n_559) );
OAI211xp5_ASAP7_75t_SL g560 ( .A1(n_539), .A2(n_530), .B(n_517), .C(n_532), .Y(n_560) );
AOI322xp5_ASAP7_75t_L g561 ( .A1(n_548), .A2(n_525), .A3(n_518), .B1(n_516), .B2(n_527), .C1(n_534), .C2(n_514), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_547), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_544), .B(n_531), .Y(n_563) );
OAI211xp5_ASAP7_75t_L g564 ( .A1(n_546), .A2(n_525), .B(n_286), .C(n_287), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_540), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_544), .A2(n_286), .B1(n_245), .B2(n_69), .C(n_65), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_552), .A2(n_541), .B1(n_542), .B2(n_555), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_557), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_549), .A2(n_241), .B1(n_287), .B2(n_552), .Y(n_569) );
AOI221xp5_ASAP7_75t_L g570 ( .A1(n_550), .A2(n_551), .B1(n_553), .B2(n_554), .C(n_556), .Y(n_570) );
OAI211xp5_ASAP7_75t_L g571 ( .A1(n_555), .A2(n_545), .B(n_539), .C(n_548), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_571), .B(n_558), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_561), .B(n_560), .C(n_564), .Y(n_573) );
NOR3xp33_ASAP7_75t_SL g574 ( .A(n_566), .B(n_567), .C(n_559), .Y(n_574) );
NAND4xp75_ASAP7_75t_L g575 ( .A(n_574), .B(n_563), .C(n_570), .D(n_569), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_573), .A2(n_563), .B1(n_565), .B2(n_568), .C(n_562), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_576), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_575), .Y(n_578) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_578), .Y(n_579) );
BUFx2_ASAP7_75t_L g580 ( .A(n_579), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_580), .A2(n_577), .B(n_572), .Y(n_581) );
endmodule