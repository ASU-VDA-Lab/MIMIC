module fake_jpeg_4600_n_180 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g15 ( 
.A(n_14),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_34),
.B(n_16),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_28),
.Y(n_44)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_56),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_40),
.B1(n_20),
.B2(n_16),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_19),
.B1(n_18),
.B2(n_30),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_75),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_40),
.B1(n_19),
.B2(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_71),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_30),
.B(n_26),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_95),
.B(n_29),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_32),
.B(n_27),
.C(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_25),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_35),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_69),
.Y(n_100)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_27),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_38),
.B1(n_33),
.B2(n_48),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_35),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_61),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_66),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_104),
.B(n_80),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_74),
.B(n_62),
.Y(n_104)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_81),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_58),
.C(n_33),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

AOI221xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.C(n_79),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_111),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_123),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_94),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_119),
.C(n_127),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_102),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_77),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_104),
.Y(n_132)
);

HAxp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_78),
.CON(n_126),
.SN(n_126)
);

OAI31xp33_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_111),
.A3(n_110),
.B(n_38),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_129),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_86),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_105),
.C(n_107),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_136),
.C(n_22),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_125),
.B(n_122),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_114),
.B1(n_103),
.B2(n_24),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_82),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_17),
.B1(n_24),
.B2(n_91),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_125),
.B1(n_103),
.B2(n_22),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_126),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_142),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_144),
.B1(n_135),
.B2(n_137),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_131),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_122),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_149),
.C(n_150),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_48),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_21),
.B(n_22),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_0),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_21),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_160),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_152),
.A2(n_142),
.B(n_136),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_159),
.B(n_154),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_23),
.B1(n_21),
.B2(n_3),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_148),
.C(n_152),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_9),
.C(n_12),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_158),
.B(n_146),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_165),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_23),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_155),
.B1(n_166),
.B2(n_4),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_170),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_155),
.B(n_11),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_4),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_7),
.B(n_13),
.C(n_1),
.D(n_2),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_175),
.C(n_171),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_177),
.B(n_173),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_169),
.C(n_1),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_1),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g180 ( 
.A(n_179),
.Y(n_180)
);


endmodule