module fake_jpeg_31810_n_112 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_56),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_39),
.B1(n_36),
.B2(n_37),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_61),
.B1(n_31),
.B2(n_3),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_35),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_1),
.Y(n_72)
);

AO22x2_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_40),
.B1(n_32),
.B2(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_71),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_55),
.B1(n_51),
.B2(n_57),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_73),
.B(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_2),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_2),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_4),
.Y(n_81)
);

HAxp5_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_3),
.CON(n_79),
.SN(n_79)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_88),
.B(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_13),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_64),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_86),
.C(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_87),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g85 ( 
.A(n_63),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_24),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_5),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_5),
.B(n_6),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_7),
.B(n_8),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_9),
.B(n_12),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_94),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_97),
.C(n_99),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_27),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

AOI21x1_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_90),
.B(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_106),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_86),
.B(n_97),
.C(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_92),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_99),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_103),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_101),
.Y(n_112)
);


endmodule