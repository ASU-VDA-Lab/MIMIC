module fake_netlist_1_8551_n_867 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_867);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_867;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_141;
wire n_119;
wire n_560;
wire n_517;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g107 ( .A(n_98), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_79), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_99), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_27), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_64), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_58), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_97), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_31), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_89), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_65), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_53), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_23), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_81), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_13), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_34), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_106), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_28), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_40), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_80), .Y(n_125) );
INVx2_ASAP7_75t_SL g126 ( .A(n_105), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_20), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_0), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_96), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_22), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_1), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_17), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_25), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_35), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
BUFx2_ASAP7_75t_SL g137 ( .A(n_74), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_72), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_41), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_1), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_18), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_61), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_93), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_36), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_25), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_34), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_73), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_71), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_20), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_110), .B(n_0), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_111), .B(n_126), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_109), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_110), .B(n_132), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_116), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_111), .B(n_2), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_132), .B(n_2), .Y(n_156) );
NOR2xp33_ASAP7_75t_SL g157 ( .A(n_107), .B(n_48), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_112), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_116), .Y(n_159) );
BUFx12f_ASAP7_75t_L g160 ( .A(n_111), .Y(n_160) );
NOR2xp33_ASAP7_75t_SL g161 ( .A(n_107), .B(n_49), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_116), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_126), .B(n_3), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_135), .B(n_3), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_112), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_135), .B(n_4), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_120), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_120), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_120), .Y(n_169) );
INVx5_ASAP7_75t_L g170 ( .A(n_126), .Y(n_170) );
BUFx8_ASAP7_75t_L g171 ( .A(n_115), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_115), .Y(n_172) );
OR2x6_ASAP7_75t_L g173 ( .A(n_153), .B(n_137), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_150), .A2(n_146), .B1(n_139), .B2(n_145), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_163), .A2(n_155), .B1(n_171), .B2(n_151), .Y(n_175) );
OAI22xp33_ASAP7_75t_R g176 ( .A1(n_155), .A2(n_145), .B1(n_128), .B2(n_140), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_163), .B(n_139), .Y(n_177) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_152), .A2(n_146), .B1(n_122), .B2(n_109), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_163), .A2(n_151), .B1(n_153), .B2(n_150), .Y(n_181) );
AO22x2_ASAP7_75t_L g182 ( .A1(n_163), .A2(n_133), .B1(n_140), .B2(n_128), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_160), .B(n_117), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_163), .B(n_128), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_153), .B(n_133), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g186 ( .A1(n_150), .A2(n_122), .B1(n_114), .B2(n_118), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_160), .B(n_117), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_155), .A2(n_149), .B1(n_121), .B2(n_123), .Y(n_188) );
OAI22xp33_ASAP7_75t_R g189 ( .A1(n_158), .A2(n_140), .B1(n_133), .B2(n_130), .Y(n_189) );
NOR2x1p5_ASAP7_75t_L g190 ( .A(n_152), .B(n_124), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_171), .A2(n_134), .B1(n_131), .B2(n_144), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_158), .B(n_129), .Y(n_192) );
OAI22xp33_ASAP7_75t_R g193 ( .A1(n_158), .A2(n_130), .B1(n_136), .B2(n_147), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_156), .A2(n_127), .B1(n_141), .B2(n_129), .Y(n_194) );
INVx5_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
NAND3x1_ASAP7_75t_L g196 ( .A(n_156), .B(n_136), .C(n_147), .Y(n_196) );
AO22x2_ASAP7_75t_L g197 ( .A1(n_151), .A2(n_137), .B1(n_5), .B2(n_6), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_171), .A2(n_120), .B1(n_148), .B2(n_142), .Y(n_198) );
OR2x6_ASAP7_75t_L g199 ( .A(n_156), .B(n_120), .Y(n_199) );
OAI22xp33_ASAP7_75t_L g200 ( .A1(n_164), .A2(n_120), .B1(n_138), .B2(n_125), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_171), .A2(n_120), .B1(n_143), .B2(n_119), .Y(n_201) );
OAI22xp33_ASAP7_75t_R g202 ( .A1(n_158), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_171), .A2(n_113), .B1(n_108), .B2(n_9), .Y(n_203) );
AO22x2_ASAP7_75t_L g204 ( .A1(n_151), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_154), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_151), .Y(n_206) );
OAI22xp33_ASAP7_75t_SL g207 ( .A1(n_164), .A2(n_7), .B1(n_8), .B2(n_10), .Y(n_207) );
OAI22xp33_ASAP7_75t_SL g208 ( .A1(n_164), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_160), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_151), .B(n_11), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g211 ( .A1(n_166), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_171), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_171), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_171), .A2(n_18), .B1(n_19), .B2(n_21), .Y(n_214) );
AO22x2_ASAP7_75t_L g215 ( .A1(n_166), .A2(n_19), .B1(n_21), .B2(n_22), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_154), .Y(n_216) );
OAI22xp33_ASAP7_75t_SL g217 ( .A1(n_166), .A2(n_23), .B1(n_24), .B2(n_26), .Y(n_217) );
OA22x2_ASAP7_75t_L g218 ( .A1(n_165), .A2(n_24), .B1(n_26), .B2(n_27), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_180), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_206), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_173), .Y(n_221) );
XNOR2x2_ASAP7_75t_L g222 ( .A(n_197), .B(n_165), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_177), .B(n_160), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_183), .A2(n_170), .B(n_165), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_181), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_182), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_192), .B(n_160), .Y(n_228) );
AND2x2_ASAP7_75t_SL g229 ( .A(n_210), .B(n_157), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_188), .B(n_165), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_179), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_182), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_179), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_195), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_205), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_179), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_216), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g238 ( .A(n_209), .B(n_157), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_205), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
XNOR2x2_ASAP7_75t_L g241 ( .A(n_197), .B(n_167), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_195), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_210), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_184), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_185), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_191), .B(n_170), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_199), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_187), .B(n_172), .Y(n_248) );
XOR2xp5_ASAP7_75t_L g249 ( .A(n_178), .B(n_28), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_199), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_215), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_173), .B(n_172), .Y(n_253) );
AND2x6_ASAP7_75t_L g254 ( .A(n_175), .B(n_172), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_203), .B(n_172), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_194), .B(n_172), .Y(n_256) );
NOR2xp67_ASAP7_75t_L g257 ( .A(n_212), .B(n_170), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_215), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_204), .Y(n_260) );
NOR2xp67_ASAP7_75t_L g261 ( .A(n_213), .B(n_170), .Y(n_261) );
XNOR2xp5_ASAP7_75t_L g262 ( .A(n_186), .B(n_190), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_214), .B(n_170), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_196), .B(n_170), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_189), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_189), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_211), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_198), .Y(n_268) );
INVxp33_ASAP7_75t_L g269 ( .A(n_174), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_207), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_200), .B(n_170), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_201), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_208), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_176), .B(n_154), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_217), .B(n_170), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_176), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_193), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_193), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_202), .Y(n_279) );
BUFx4f_ASAP7_75t_SL g280 ( .A(n_254), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_235), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_225), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_274), .B(n_170), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_267), .B(n_170), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_235), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_239), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_267), .B(n_170), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_239), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_225), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_219), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_219), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_274), .B(n_170), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_253), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_220), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_226), .B(n_170), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_226), .B(n_154), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_227), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_230), .B(n_157), .Y(n_298) );
OAI21xp5_ASAP7_75t_L g299 ( .A1(n_275), .A2(n_224), .B(n_268), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_243), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_243), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_254), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_245), .B(n_154), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_227), .Y(n_304) );
NOR2xp33_ASAP7_75t_R g305 ( .A(n_229), .B(n_161), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_254), .Y(n_306) );
INVx2_ASAP7_75t_SL g307 ( .A(n_229), .Y(n_307) );
NOR2xp33_ASAP7_75t_SL g308 ( .A(n_229), .B(n_161), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_223), .B(n_154), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_221), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_237), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g312 ( .A1(n_268), .A2(n_154), .B(n_167), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_247), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_220), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_245), .B(n_270), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_254), .B(n_154), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_270), .B(n_202), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_234), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_237), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_234), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_232), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_234), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_254), .B(n_162), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_277), .B(n_29), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_237), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_264), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_232), .Y(n_327) );
NOR2xp33_ASAP7_75t_R g328 ( .A(n_254), .B(n_161), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_273), .B(n_159), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_285), .B(n_265), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_285), .Y(n_334) );
OR2x6_ASAP7_75t_L g335 ( .A(n_302), .B(n_259), .Y(n_335) );
BUFx8_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
BUFx12f_ASAP7_75t_L g337 ( .A(n_310), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_282), .B(n_253), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_315), .B(n_276), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_282), .B(n_260), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_286), .B(n_265), .Y(n_341) );
BUFx4f_ASAP7_75t_L g342 ( .A(n_286), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_293), .B(n_269), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_315), .B(n_276), .Y(n_344) );
BUFx4f_ASAP7_75t_L g345 ( .A(n_286), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_286), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_315), .B(n_277), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_286), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_281), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_293), .B(n_266), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_283), .B(n_266), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_282), .B(n_260), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_281), .Y(n_354) );
NOR2xp33_ASAP7_75t_SL g355 ( .A(n_280), .B(n_254), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_281), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_283), .B(n_244), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_311), .Y(n_358) );
BUFx4f_ASAP7_75t_L g359 ( .A(n_307), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_283), .B(n_244), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_315), .B(n_278), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_342), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_342), .Y(n_363) );
BUFx24_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_331), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_342), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_342), .Y(n_367) );
INVx4_ASAP7_75t_L g368 ( .A(n_342), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_342), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_331), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_345), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_331), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_334), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_330), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_330), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_345), .B(n_302), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_348), .A2(n_324), .B1(n_252), .B2(n_258), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_348), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_334), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_334), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_337), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_334), .Y(n_382) );
BUFx2_ASAP7_75t_SL g383 ( .A(n_334), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_352), .A2(n_317), .B1(n_279), .B2(n_222), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_345), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_346), .Y(n_387) );
BUFx12f_ASAP7_75t_L g388 ( .A(n_336), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_345), .Y(n_389) );
CKINVDCx6p67_ASAP7_75t_R g390 ( .A(n_335), .Y(n_390) );
INVx4_ASAP7_75t_L g391 ( .A(n_388), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_388), .A2(n_279), .B1(n_317), .B2(n_278), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_381), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_365), .A2(n_345), .B1(n_324), .B2(n_280), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_388), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_378), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_388), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_388), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_365), .A2(n_345), .B1(n_324), .B2(n_280), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_381), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_378), .Y(n_402) );
BUFx2_ASAP7_75t_SL g403 ( .A(n_365), .Y(n_403) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_390), .A2(n_324), .B1(n_355), .B2(n_337), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_373), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_385), .B(n_317), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_385), .A2(n_343), .B1(n_351), .B2(n_352), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_378), .B(n_373), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_378), .B(n_346), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_388), .A2(n_306), .B1(n_302), .B2(n_343), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g413 ( .A1(n_383), .A2(n_222), .B1(n_241), .B2(n_337), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_383), .A2(n_241), .B1(n_337), .B2(n_308), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_385), .A2(n_306), .B1(n_298), .B2(n_352), .Y(n_415) );
CKINVDCx6p67_ASAP7_75t_R g416 ( .A(n_364), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_375), .A2(n_351), .B1(n_352), .B2(n_298), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_373), .B(n_348), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_370), .Y(n_419) );
CKINVDCx6p67_ASAP7_75t_R g420 ( .A(n_364), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_390), .A2(n_306), .B1(n_298), .B2(n_254), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_375), .A2(n_361), .B1(n_347), .B2(n_355), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_390), .A2(n_355), .B1(n_337), .B2(n_308), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_390), .A2(n_306), .B1(n_335), .B2(n_358), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_373), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_373), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_387), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_390), .A2(n_249), .B1(n_273), .B2(n_307), .Y(n_428) );
BUFx2_ASAP7_75t_SL g429 ( .A(n_370), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_372), .B(n_347), .Y(n_431) );
BUFx8_ASAP7_75t_L g432 ( .A(n_384), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_416), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_416), .Y(n_434) );
OAI22xp5_ASAP7_75t_SL g435 ( .A1(n_391), .A2(n_249), .B1(n_381), .B2(n_383), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_420), .A2(n_383), .B1(n_370), .B2(n_374), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_391), .A2(n_368), .B1(n_307), .B2(n_336), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g438 ( .A1(n_406), .A2(n_428), .B1(n_262), .B2(n_361), .C1(n_347), .C2(n_392), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_391), .A2(n_368), .B1(n_307), .B2(n_336), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
NOR2x1_ASAP7_75t_R g441 ( .A(n_399), .B(n_395), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_399), .A2(n_368), .B1(n_307), .B2(n_336), .Y(n_442) );
INVx6_ASAP7_75t_L g443 ( .A(n_432), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_397), .Y(n_444) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_404), .A2(n_384), .B(n_262), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_399), .A2(n_368), .B1(n_336), .B2(n_384), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_420), .A2(n_383), .B1(n_374), .B2(n_368), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_418), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_432), .A2(n_368), .B1(n_336), .B2(n_384), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_411), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_403), .A2(n_374), .B1(n_368), .B2(n_384), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_402), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g455 ( .A1(n_395), .A2(n_368), .B1(n_366), .B2(n_363), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_432), .A2(n_368), .B1(n_336), .B2(n_360), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_408), .B(n_387), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_432), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_418), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_403), .A2(n_368), .B1(n_379), .B2(n_372), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_412), .Y(n_461) );
OAI21xp5_ASAP7_75t_SL g462 ( .A1(n_413), .A2(n_377), .B(n_364), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_408), .B(n_372), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_398), .A2(n_308), .B1(n_335), .B2(n_367), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_398), .A2(n_361), .B1(n_377), .B2(n_344), .C1(n_339), .C2(n_251), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_417), .A2(n_379), .B1(n_372), .B2(n_367), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_425), .B(n_387), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_407), .A2(n_377), .B1(n_360), .B2(n_357), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_409), .B(n_387), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_425), .B(n_387), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_426), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_426), .Y(n_473) );
BUFx12f_ASAP7_75t_L g474 ( .A(n_418), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_427), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_427), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_418), .B(n_387), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_393), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_424), .A2(n_366), .B1(n_371), .B2(n_369), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_394), .A2(n_366), .B1(n_371), .B2(n_369), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_430), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_396), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_430), .B(n_379), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g484 ( .A1(n_417), .A2(n_335), .B1(n_367), .B2(n_369), .Y(n_484) );
OAI21xp5_ASAP7_75t_SL g485 ( .A1(n_414), .A2(n_377), .B(n_376), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_400), .A2(n_366), .B1(n_371), .B2(n_369), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_407), .A2(n_335), .B1(n_367), .B2(n_363), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_405), .B(n_380), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_415), .A2(n_357), .B1(n_360), .B2(n_338), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_419), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_419), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_422), .A2(n_367), .B1(n_335), .B2(n_363), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_422), .A2(n_335), .B1(n_363), .B2(n_366), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_421), .A2(n_360), .B1(n_357), .B2(n_338), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_423), .A2(n_357), .B1(n_338), .B2(n_258), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_410), .A2(n_338), .B1(n_252), .B2(n_257), .Y(n_496) );
BUFx12f_ASAP7_75t_L g497 ( .A(n_409), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_429), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_429), .B(n_380), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_431), .A2(n_338), .B1(n_257), .B2(n_261), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_401), .A2(n_338), .B1(n_261), .B2(n_305), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_411), .Y(n_502) );
OAI221xp5_ASAP7_75t_L g503 ( .A1(n_445), .A2(n_251), .B1(n_344), .B2(n_339), .C(n_310), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_451), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_438), .A2(n_305), .B1(n_328), .B2(n_338), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_435), .A2(n_305), .B1(n_328), .B2(n_369), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_468), .B(n_380), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_435), .A2(n_328), .B1(n_363), .B2(n_366), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_457), .B(n_380), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_497), .A2(n_371), .B1(n_363), .B2(n_369), .Y(n_510) );
AO22x1_ASAP7_75t_L g511 ( .A1(n_433), .A2(n_369), .B1(n_371), .B2(n_389), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_497), .A2(n_371), .B1(n_340), .B2(n_353), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_497), .A2(n_371), .B1(n_340), .B2(n_353), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_471), .B(n_380), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_487), .A2(n_353), .B1(n_340), .B2(n_263), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_484), .A2(n_353), .B1(n_340), .B2(n_263), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_458), .B(n_380), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_469), .A2(n_353), .B1(n_340), .B2(n_263), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_462), .A2(n_389), .B1(n_386), .B2(n_362), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_469), .A2(n_339), .B1(n_344), .B2(n_341), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_466), .A2(n_474), .B1(n_493), .B2(n_492), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_445), .A2(n_332), .B1(n_341), .B2(n_340), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_466), .A2(n_340), .B1(n_353), .B2(n_263), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_474), .A2(n_353), .B1(n_332), .B2(n_341), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_462), .A2(n_380), .B1(n_382), .B2(n_346), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_495), .A2(n_341), .B1(n_332), .B2(n_326), .Y(n_526) );
OAI221xp5_ASAP7_75t_SL g527 ( .A1(n_485), .A2(n_316), .B1(n_293), .B2(n_256), .C(n_323), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_456), .A2(n_332), .B1(n_326), .B2(n_386), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_482), .B(n_159), .C(n_162), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_443), .A2(n_389), .B1(n_386), .B2(n_362), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_443), .A2(n_389), .B1(n_386), .B2(n_362), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_450), .A2(n_380), .B1(n_382), .B2(n_346), .Y(n_532) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_485), .A2(n_312), .B(n_323), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_443), .A2(n_389), .B1(n_386), .B2(n_362), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_443), .A2(n_326), .B1(n_386), .B2(n_389), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_471), .B(n_380), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_489), .A2(n_346), .B1(n_333), .B2(n_350), .Y(n_537) );
OAI222xp33_ASAP7_75t_L g538 ( .A1(n_458), .A2(n_362), .B1(n_376), .B2(n_356), .C1(n_354), .C2(n_350), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_479), .A2(n_326), .B1(n_362), .B2(n_282), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g540 ( .A(n_441), .B(n_434), .C(n_433), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_457), .B(n_461), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_446), .A2(n_362), .B1(n_376), .B2(n_380), .Y(n_542) );
AOI21xp5_ASAP7_75t_SL g543 ( .A1(n_441), .A2(n_382), .B(n_380), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_464), .A2(n_326), .B1(n_362), .B2(n_282), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_433), .A2(n_326), .B1(n_289), .B2(n_329), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_433), .A2(n_326), .B1(n_289), .B2(n_329), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_434), .A2(n_382), .B1(n_380), .B2(n_376), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_461), .B(n_380), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_434), .A2(n_382), .B1(n_380), .B2(n_376), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_434), .A2(n_376), .B1(n_382), .B2(n_350), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_494), .A2(n_326), .B1(n_289), .B2(n_329), .Y(n_551) );
NOR3xp33_ASAP7_75t_L g552 ( .A(n_498), .B(n_329), .C(n_316), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_480), .A2(n_326), .B1(n_289), .B2(n_354), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_455), .A2(n_376), .B1(n_382), .B2(n_356), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_467), .A2(n_452), .B1(n_500), .B2(n_501), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_448), .A2(n_382), .B1(n_376), .B2(n_333), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_436), .A2(n_382), .B1(n_333), .B2(n_356), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_486), .A2(n_289), .B1(n_354), .B2(n_299), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_437), .A2(n_299), .B1(n_333), .B2(n_316), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_465), .B(n_382), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_439), .A2(n_299), .B1(n_333), .B2(n_296), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_442), .A2(n_382), .B1(n_358), .B2(n_333), .Y(n_562) );
OAI222xp33_ASAP7_75t_L g563 ( .A1(n_460), .A2(n_333), .B1(n_358), .B2(n_349), .C1(n_323), .C2(n_314), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_477), .A2(n_382), .B1(n_358), .B2(n_349), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_496), .A2(n_296), .B1(n_382), .B2(n_314), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_459), .A2(n_296), .B1(n_382), .B2(n_314), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_478), .A2(n_382), .B1(n_314), .B2(n_349), .Y(n_567) );
NAND3xp33_ASAP7_75t_L g568 ( .A(n_465), .B(n_162), .C(n_159), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_459), .A2(n_296), .B1(n_291), .B2(n_294), .Y(n_569) );
AOI221xp5_ASAP7_75t_SL g570 ( .A1(n_440), .A2(n_159), .B1(n_162), .B2(n_313), .C(n_303), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_451), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_449), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_459), .A2(n_349), .B1(n_303), .B2(n_359), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_459), .A2(n_349), .B1(n_303), .B2(n_359), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_498), .A2(n_303), .B1(n_238), .B2(n_255), .C(n_309), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_449), .A2(n_296), .B1(n_291), .B2(n_294), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_449), .A2(n_440), .B1(n_453), .B2(n_447), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_449), .A2(n_296), .B1(n_291), .B2(n_294), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_449), .A2(n_359), .B1(n_255), .B2(n_296), .Y(n_579) );
OAI222xp33_ASAP7_75t_L g580 ( .A1(n_472), .A2(n_481), .B1(n_463), .B2(n_454), .C1(n_451), .C2(n_476), .Y(n_580) );
AOI222xp33_ASAP7_75t_L g581 ( .A1(n_444), .A2(n_296), .B1(n_327), .B2(n_290), .C1(n_301), .C2(n_300), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_454), .B(n_159), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_470), .A2(n_313), .B1(n_290), .B2(n_359), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_472), .B(n_327), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_449), .A2(n_290), .B1(n_304), .B2(n_321), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_444), .A2(n_321), .B1(n_304), .B2(n_297), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_447), .A2(n_321), .B1(n_304), .B2(n_297), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_481), .A2(n_313), .B1(n_359), .B2(n_297), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_453), .A2(n_327), .B1(n_359), .B2(n_288), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_454), .B(n_159), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_483), .A2(n_327), .B1(n_359), .B2(n_288), .Y(n_591) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_499), .A2(n_283), .B1(n_292), .B2(n_309), .Y(n_592) );
OAI222xp33_ASAP7_75t_L g593 ( .A1(n_473), .A2(n_309), .B1(n_264), .B2(n_288), .C1(n_325), .C2(n_311), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_473), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_473), .B(n_29), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_502), .A2(n_312), .B(n_325), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_475), .B(n_159), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_502), .A2(n_325), .B1(n_319), .B2(n_311), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_483), .A2(n_300), .B1(n_301), .B2(n_292), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_541), .B(n_475), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_509), .B(n_490), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_509), .B(n_490), .Y(n_602) );
NAND4xp25_ASAP7_75t_L g603 ( .A(n_521), .B(n_238), .C(n_491), .D(n_490), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_533), .B(n_491), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_571), .B(n_475), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_594), .B(n_476), .Y(n_606) );
NAND4xp25_ASAP7_75t_L g607 ( .A(n_503), .B(n_491), .C(n_499), .D(n_502), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_504), .B(n_488), .Y(n_608) );
NOR2xp33_ASAP7_75t_SL g609 ( .A(n_540), .B(n_488), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_529), .B(n_159), .C(n_162), .Y(n_610) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_522), .B(n_228), .C(n_167), .D(n_292), .Y(n_611) );
NOR3xp33_ASAP7_75t_SL g612 ( .A(n_527), .B(n_246), .C(n_284), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_533), .B(n_167), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_533), .B(n_168), .Y(n_614) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_525), .A2(n_292), .B1(n_159), .B2(n_162), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_533), .B(n_168), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_507), .B(n_159), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_522), .A2(n_325), .B1(n_311), .B2(n_319), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_572), .B(n_168), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_577), .B(n_168), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_514), .B(n_159), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_536), .B(n_162), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_520), .B(n_162), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_520), .B(n_162), .Y(n_624) );
NAND3xp33_ASAP7_75t_SL g625 ( .A(n_525), .B(n_30), .C(n_31), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_555), .B(n_162), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_523), .A2(n_325), .B1(n_319), .B2(n_320), .Y(n_627) );
OAI21xp5_ASAP7_75t_SL g628 ( .A1(n_547), .A2(n_162), .B(n_250), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_529), .B(n_162), .C(n_168), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_570), .B(n_168), .C(n_169), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_570), .B(n_543), .C(n_549), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g632 ( .A1(n_505), .A2(n_300), .B1(n_301), .B2(n_312), .C(n_284), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_555), .B(n_30), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_548), .B(n_32), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_582), .B(n_168), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_516), .B(n_287), .C(n_284), .D(n_271), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_543), .B(n_168), .C(n_169), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_560), .B(n_32), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_515), .A2(n_295), .B1(n_287), .B2(n_301), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_554), .A2(n_295), .B1(n_319), .B2(n_320), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_582), .B(n_168), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_590), .B(n_33), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_590), .B(n_33), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_597), .B(n_35), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_580), .A2(n_168), .B1(n_169), .B2(n_300), .C(n_287), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_595), .B(n_36), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_567), .B(n_37), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g648 ( .A1(n_511), .A2(n_168), .B(n_169), .C(n_247), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_556), .B(n_168), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_592), .A2(n_295), .B1(n_322), .B2(n_320), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_517), .B(n_38), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_552), .A2(n_295), .B1(n_322), .B2(n_320), .Y(n_652) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_518), .A2(n_250), .B1(n_272), .B2(n_319), .C(n_318), .Y(n_653) );
NOR2xp33_ASAP7_75t_R g654 ( .A(n_512), .B(n_38), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_568), .B(n_169), .C(n_295), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_542), .A2(n_295), .B1(n_322), .B2(n_318), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_538), .A2(n_295), .B(n_169), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_513), .A2(n_320), .B1(n_318), .B2(n_322), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_583), .B(n_39), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_534), .A2(n_295), .B(n_169), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_583), .B(n_39), .Y(n_661) );
NOR2xp33_ASAP7_75t_SL g662 ( .A(n_593), .B(n_318), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_598), .B(n_40), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_575), .A2(n_169), .B1(n_322), .B2(n_318), .C(n_248), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_557), .A2(n_169), .B(n_42), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_598), .B(n_41), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_568), .B(n_322), .C(n_268), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_599), .B(n_42), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_599), .B(n_43), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_532), .A2(n_322), .B1(n_242), .B2(n_240), .C(n_46), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_584), .B(n_43), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_564), .B(n_44), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_564), .B(n_44), .Y(n_673) );
AOI221xp5_ASAP7_75t_SL g674 ( .A1(n_519), .A2(n_45), .B1(n_47), .B2(n_272), .C(n_51), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_558), .B(n_45), .C(n_234), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_511), .B(n_50), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_544), .B(n_52), .Y(n_677) );
OAI21xp33_ASAP7_75t_L g678 ( .A1(n_573), .A2(n_54), .B(n_55), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g679 ( .A1(n_550), .A2(n_56), .B(n_57), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_510), .B(n_59), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_562), .A2(n_236), .B1(n_233), .B2(n_231), .C(n_66), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_524), .A2(n_60), .B1(n_62), .B2(n_63), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_508), .B(n_67), .Y(n_683) );
AOI221x1_ASAP7_75t_SL g684 ( .A1(n_588), .A2(n_68), .B1(n_69), .B2(n_70), .C(n_75), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_581), .B(n_76), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_574), .B(n_77), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_561), .B(n_78), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_553), .B(n_539), .C(n_535), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_530), .B(n_82), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_579), .A2(n_83), .B(n_86), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_531), .B(n_87), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_506), .A2(n_88), .B1(n_90), .B2(n_91), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_591), .B(n_92), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_596), .B(n_94), .Y(n_694) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_605), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_633), .B(n_588), .C(n_563), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_601), .B(n_528), .Y(n_697) );
NAND4xp75_ASAP7_75t_L g698 ( .A(n_674), .B(n_537), .C(n_596), .D(n_581), .Y(n_698) );
OA21x2_ASAP7_75t_L g699 ( .A1(n_604), .A2(n_566), .B(n_537), .Y(n_699) );
AO21x2_ASAP7_75t_L g700 ( .A1(n_614), .A2(n_559), .B(n_589), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_631), .B(n_578), .C(n_576), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_600), .B(n_526), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_601), .B(n_569), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_602), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_626), .B(n_565), .C(n_585), .Y(n_705) );
INVx3_ASAP7_75t_SL g706 ( .A(n_686), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_604), .B(n_546), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_637), .B(n_545), .C(n_586), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_602), .B(n_551), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_675), .B(n_587), .C(n_236), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_613), .B(n_95), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_665), .B(n_233), .C(n_231), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_608), .B(n_100), .Y(n_713) );
NAND4xp75_ASAP7_75t_L g714 ( .A(n_686), .B(n_101), .C(n_102), .D(n_103), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_613), .B(n_104), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_606), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_614), .B(n_616), .Y(n_717) );
NOR2xp33_ASAP7_75t_SL g718 ( .A(n_609), .B(n_690), .Y(n_718) );
OA211x2_ASAP7_75t_L g719 ( .A1(n_662), .A2(n_625), .B(n_691), .C(n_689), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_617), .B(n_621), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_622), .B(n_619), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_616), .B(n_619), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_635), .B(n_641), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_603), .A2(n_611), .B1(n_654), .B2(n_688), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_635), .B(n_641), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_628), .A2(n_660), .B1(n_690), .B2(n_685), .Y(n_726) );
OA21x2_ASAP7_75t_L g727 ( .A1(n_676), .A2(n_620), .B(n_649), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_649), .B(n_620), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_654), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_656), .B(n_694), .Y(n_730) );
NAND4xp75_ASAP7_75t_L g731 ( .A(n_689), .B(n_691), .C(n_612), .D(n_683), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_668), .A2(n_669), .B1(n_661), .B2(n_659), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_646), .B(n_651), .C(n_638), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_634), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_623), .B(n_624), .Y(n_735) );
AO21x2_ASAP7_75t_L g736 ( .A1(n_672), .A2(n_673), .B(n_647), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_648), .B(n_645), .C(n_615), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_642), .B(n_643), .Y(n_738) );
NOR2xp33_ASAP7_75t_SL g739 ( .A(n_678), .B(n_653), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_671), .B(n_632), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_644), .Y(n_741) );
NOR3xp33_ASAP7_75t_SL g742 ( .A(n_618), .B(n_682), .C(n_692), .Y(n_742) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_670), .B(n_663), .C(n_666), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_610), .B(n_629), .C(n_640), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_636), .A2(n_664), .B1(n_650), .B2(n_652), .Y(n_745) );
OAI211xp5_ASAP7_75t_SL g746 ( .A1(n_639), .A2(n_679), .B(n_681), .C(n_658), .Y(n_746) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_655), .B(n_667), .C(n_630), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_683), .B(n_680), .C(n_687), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_627), .B(n_680), .Y(n_749) );
NOR2x1_ASAP7_75t_L g750 ( .A(n_693), .B(n_677), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_684), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_677), .B(n_633), .C(n_626), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_603), .A2(n_503), .B1(n_438), .B2(n_521), .Y(n_753) );
NAND3xp33_ASAP7_75t_SL g754 ( .A(n_654), .B(n_657), .C(n_665), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_600), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_601), .B(n_602), .Y(n_756) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_631), .B(n_626), .C(n_633), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_601), .B(n_602), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_631), .B(n_626), .C(n_633), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_601), .B(n_602), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_633), .B(n_607), .Y(n_761) );
NOR2xp33_ASAP7_75t_SL g762 ( .A(n_609), .B(n_441), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_603), .A2(n_503), .B1(n_438), .B2(n_521), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_695), .B(n_755), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_704), .B(n_756), .Y(n_765) );
OAI22xp33_ASAP7_75t_SL g766 ( .A1(n_706), .A2(n_762), .B1(n_718), .B2(n_729), .Y(n_766) );
XOR2x2_ASAP7_75t_L g767 ( .A(n_706), .B(n_754), .Y(n_767) );
XNOR2x2_ASAP7_75t_L g768 ( .A(n_731), .B(n_698), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_716), .B(n_761), .Y(n_769) );
NOR2x1_ASAP7_75t_L g770 ( .A(n_757), .B(n_759), .Y(n_770) );
INVx6_ASAP7_75t_L g771 ( .A(n_728), .Y(n_771) );
INVx3_ASAP7_75t_L g772 ( .A(n_717), .Y(n_772) );
XOR2xp5_ASAP7_75t_L g773 ( .A(n_738), .B(n_725), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_761), .B(n_736), .Y(n_774) );
NOR4xp25_ASAP7_75t_L g775 ( .A(n_751), .B(n_734), .C(n_741), .D(n_724), .Y(n_775) );
INVxp67_ASAP7_75t_L g776 ( .A(n_702), .Y(n_776) );
NAND4xp75_ASAP7_75t_L g777 ( .A(n_719), .B(n_750), .C(n_726), .D(n_742), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_758), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_736), .B(n_697), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_736), .B(n_697), .Y(n_780) );
NAND4xp75_ASAP7_75t_L g781 ( .A(n_740), .B(n_727), .C(n_699), .D(n_709), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_717), .Y(n_782) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_760), .Y(n_783) );
XNOR2x1_ASAP7_75t_L g784 ( .A(n_748), .B(n_730), .Y(n_784) );
INVxp67_ASAP7_75t_L g785 ( .A(n_733), .Y(n_785) );
NAND4xp75_ASAP7_75t_L g786 ( .A(n_727), .B(n_699), .C(n_709), .D(n_735), .Y(n_786) );
INVxp67_ASAP7_75t_L g787 ( .A(n_739), .Y(n_787) );
AND2x4_ASAP7_75t_SL g788 ( .A(n_723), .B(n_722), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_724), .A2(n_763), .B1(n_753), .B2(n_752), .Y(n_789) );
NAND4xp75_ASAP7_75t_L g790 ( .A(n_711), .B(n_715), .C(n_730), .D(n_699), .Y(n_790) );
AND4x2_ASAP7_75t_L g791 ( .A(n_753), .B(n_763), .C(n_696), .D(n_732), .Y(n_791) );
XOR2xp5_ASAP7_75t_L g792 ( .A(n_703), .B(n_721), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_743), .A2(n_701), .B1(n_707), .B2(n_732), .Y(n_793) );
XNOR2xp5_ASAP7_75t_L g794 ( .A(n_723), .B(n_705), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_728), .B(n_700), .Y(n_795) );
NAND4xp75_ASAP7_75t_L g796 ( .A(n_712), .B(n_746), .C(n_714), .D(n_708), .Y(n_796) );
XNOR2xp5_ASAP7_75t_L g797 ( .A(n_768), .B(n_745), .Y(n_797) );
XNOR2x2_ASAP7_75t_L g798 ( .A(n_767), .B(n_744), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_764), .Y(n_799) );
XOR2x2_ASAP7_75t_L g800 ( .A(n_767), .B(n_737), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_783), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_765), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_776), .B(n_700), .Y(n_803) );
INVx1_ASAP7_75t_SL g804 ( .A(n_788), .Y(n_804) );
XNOR2xp5_ASAP7_75t_L g805 ( .A(n_768), .B(n_745), .Y(n_805) );
INVx1_ASAP7_75t_SL g806 ( .A(n_788), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_789), .B(n_749), .Y(n_807) );
XNOR2x1_ASAP7_75t_SL g808 ( .A(n_791), .B(n_710), .Y(n_808) );
INVx2_ASAP7_75t_SL g809 ( .A(n_771), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_778), .Y(n_810) );
XOR2x2_ASAP7_75t_L g811 ( .A(n_777), .B(n_747), .Y(n_811) );
INVx2_ASAP7_75t_SL g812 ( .A(n_771), .Y(n_812) );
INVx1_ASAP7_75t_SL g813 ( .A(n_771), .Y(n_813) );
XNOR2x2_ASAP7_75t_L g814 ( .A(n_781), .B(n_713), .Y(n_814) );
OA22x2_ASAP7_75t_L g815 ( .A1(n_793), .A2(n_700), .B1(n_720), .B2(n_787), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_772), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_774), .B(n_795), .Y(n_817) );
INVxp67_ASAP7_75t_L g818 ( .A(n_777), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_795), .B(n_769), .Y(n_819) );
XOR2x2_ASAP7_75t_L g820 ( .A(n_794), .B(n_784), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_802), .Y(n_821) );
OAI22x1_ASAP7_75t_L g822 ( .A1(n_797), .A2(n_770), .B1(n_794), .B2(n_785), .Y(n_822) );
XNOR2x1_ASAP7_75t_L g823 ( .A(n_797), .B(n_796), .Y(n_823) );
OA22x2_ASAP7_75t_L g824 ( .A1(n_805), .A2(n_791), .B1(n_773), .B2(n_792), .Y(n_824) );
INVx4_ASAP7_75t_L g825 ( .A(n_811), .Y(n_825) );
XOR2x2_ASAP7_75t_L g826 ( .A(n_800), .B(n_766), .Y(n_826) );
XOR2x2_ASAP7_75t_L g827 ( .A(n_800), .B(n_796), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_816), .Y(n_828) );
BUFx3_ASAP7_75t_L g829 ( .A(n_798), .Y(n_829) );
OA22x2_ASAP7_75t_L g830 ( .A1(n_818), .A2(n_780), .B1(n_779), .B2(n_775), .Y(n_830) );
BUFx2_ASAP7_75t_L g831 ( .A(n_804), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_798), .Y(n_832) );
XNOR2xp5_ASAP7_75t_L g833 ( .A(n_820), .B(n_784), .Y(n_833) );
OAI22x1_ASAP7_75t_L g834 ( .A1(n_807), .A2(n_782), .B1(n_772), .B2(n_786), .Y(n_834) );
XNOR2xp5_ASAP7_75t_L g835 ( .A(n_820), .B(n_790), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_831), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_821), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_830), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_828), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_828), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_830), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_829), .Y(n_842) );
OAI322xp33_ASAP7_75t_L g843 ( .A1(n_832), .A2(n_815), .A3(n_807), .B1(n_814), .B2(n_803), .C1(n_817), .C2(n_808), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_836), .Y(n_844) );
AO22x2_ASAP7_75t_L g845 ( .A1(n_842), .A2(n_823), .B1(n_825), .B2(n_829), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_836), .A2(n_835), .B1(n_832), .B2(n_833), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_839), .Y(n_847) );
AND4x1_ASAP7_75t_L g848 ( .A(n_838), .B(n_827), .C(n_825), .D(n_823), .Y(n_848) );
O2A1O1Ixp33_ASAP7_75t_L g849 ( .A1(n_846), .A2(n_842), .B(n_841), .C(n_843), .Y(n_849) );
O2A1O1Ixp33_ASAP7_75t_L g850 ( .A1(n_844), .A2(n_827), .B(n_825), .C(n_837), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_847), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_851), .Y(n_852) );
AO22x1_ASAP7_75t_L g853 ( .A1(n_849), .A2(n_848), .B1(n_845), .B2(n_837), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_853), .A2(n_824), .B1(n_822), .B2(n_826), .Y(n_854) );
AOI22xp33_ASAP7_75t_SL g855 ( .A1(n_852), .A2(n_824), .B1(n_845), .B2(n_848), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_854), .Y(n_856) );
AND4x1_ASAP7_75t_L g857 ( .A(n_855), .B(n_850), .C(n_808), .D(n_822), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_856), .Y(n_858) );
AO22x2_ASAP7_75t_L g859 ( .A1(n_857), .A2(n_826), .B1(n_840), .B2(n_806), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_858), .A2(n_811), .B1(n_815), .B2(n_834), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_860), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g862 ( .A1(n_861), .A2(n_859), .B1(n_834), .B2(n_799), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_862), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_863), .A2(n_840), .B1(n_819), .B2(n_813), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_864), .Y(n_865) );
AOI221xp5_ASAP7_75t_L g866 ( .A1(n_865), .A2(n_801), .B1(n_809), .B2(n_812), .C(n_816), .Y(n_866) );
AOI211xp5_ASAP7_75t_L g867 ( .A1(n_866), .A2(n_809), .B(n_812), .C(n_810), .Y(n_867) );
endmodule