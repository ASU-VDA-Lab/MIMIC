module fake_jpeg_23594_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_39),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g38 ( 
.A(n_26),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_2),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_52),
.Y(n_58)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_28),
.B1(n_31),
.B2(n_22),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_28),
.B1(n_31),
.B2(n_22),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_38),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_28),
.B1(n_22),
.B2(n_31),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_19),
.B1(n_16),
.B2(n_26),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_65),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_39),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_73),
.C(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_51),
.Y(n_67)
);

HB1xp67_ASAP7_75t_SL g93 ( 
.A(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_54),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_80),
.B1(n_86),
.B2(n_29),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_35),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_32),
.B(n_19),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_36),
.B1(n_30),
.B2(n_26),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_34),
.B1(n_32),
.B2(n_16),
.Y(n_89)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_45),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_45),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_29),
.B1(n_19),
.B2(n_16),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_37),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_17),
.C(n_20),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_99),
.B1(n_77),
.B2(n_60),
.Y(n_119)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_71),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_58),
.B(n_79),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_103),
.B1(n_114),
.B2(n_69),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_29),
.B1(n_23),
.B2(n_27),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_37),
.B1(n_20),
.B2(n_21),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_21),
.B1(n_27),
.B2(n_23),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_86),
.B1(n_88),
.B2(n_61),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_104),
.C(n_95),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_25),
.B1(n_24),
.B2(n_17),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_129),
.B1(n_91),
.B2(n_110),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_118),
.B1(n_125),
.B2(n_140),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_115),
.A2(n_74),
.B1(n_79),
.B2(n_60),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_132),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_74),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_123),
.B(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_81),
.B1(n_65),
.B2(n_87),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_98),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_127),
.B(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_82),
.B1(n_67),
.B2(n_70),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_24),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_93),
.A2(n_21),
.B(n_18),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_91),
.B1(n_96),
.B2(n_90),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_98),
.Y(n_135)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_18),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_18),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_21),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_142),
.B(n_66),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_66),
.B1(n_14),
.B2(n_13),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_14),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_100),
.C(n_110),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_103),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_149),
.A2(n_162),
.B(n_164),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_160),
.B1(n_165),
.B2(n_166),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_161),
.B1(n_129),
.B2(n_141),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_103),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_120),
.C(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_11),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_135),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_96),
.B1(n_101),
.B2(n_92),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_101),
.B1(n_92),
.B2(n_102),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_102),
.B(n_4),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_5),
.B(n_6),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_170),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_140),
.B1(n_125),
.B2(n_122),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_183),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_173),
.Y(n_195)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_121),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_181),
.C(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_182),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_142),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_176),
.Y(n_191)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_133),
.C(n_9),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_8),
.C(n_10),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_11),
.C(n_12),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_205),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_201),
.C(n_203),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_152),
.C(n_158),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_155),
.C(n_161),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_170),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_210),
.B(n_211),
.Y(n_230)
);

HAxp5_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_188),
.CON(n_208),
.SN(n_208)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_146),
.B1(n_171),
.B2(n_153),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_213),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_185),
.B(n_188),
.C(n_149),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_195),
.A2(n_164),
.B(n_185),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_144),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_189),
.C(n_148),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_216),
.C(n_196),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_201),
.C(n_203),
.Y(n_216)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_204),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_205),
.B1(n_155),
.B2(n_193),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_180),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_225),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_169),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_160),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_228),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_191),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_215),
.B(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_223),
.B(n_218),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_236),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

XOR2x1_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_184),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_228),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_242),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_230),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_231),
.Y(n_245)
);

OAI221xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_237),
.B1(n_235),
.B2(n_229),
.C(n_187),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_244),
.B(n_165),
.C(n_146),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_224),
.C(n_154),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_163),
.B(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_252),
.B(n_247),
.C(n_11),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_149),
.Y(n_252)
);

AO21x2_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_12),
.B(n_253),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_255),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_256),
.Y(n_257)
);


endmodule