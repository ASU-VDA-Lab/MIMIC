module fake_jpeg_11189_n_636 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_636);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_636;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_31),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_60),
.B(n_72),
.Y(n_151)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_37),
.Y(n_62)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_31),
.B(n_9),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_94),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_78),
.Y(n_220)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_80),
.Y(n_221)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_81),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_83),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_85),
.Y(n_197)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_92),
.Y(n_192)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_8),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_96),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_97),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_8),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_98),
.B(n_112),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_99),
.Y(n_211)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_105),
.Y(n_216)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_111),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_45),
.B(n_10),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_20),
.Y(n_115)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_26),
.Y(n_117)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_118),
.A2(n_57),
.B1(n_51),
.B2(n_44),
.Y(n_189)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_29),
.B(n_7),
.C(n_17),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_123),
.Y(n_169)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_29),
.Y(n_122)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_45),
.B(n_7),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_30),
.Y(n_125)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_34),
.Y(n_127)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_45),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_56),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_53),
.B(n_7),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_129),
.B(n_14),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_53),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_133),
.B(n_138),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_56),
.B1(n_54),
.B2(n_34),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_137),
.A2(n_167),
.B1(n_168),
.B2(n_173),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_53),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_141),
.B(n_92),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_111),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_145),
.B(n_210),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_71),
.A2(n_23),
.B1(n_51),
.B2(n_44),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_153),
.A2(n_189),
.B1(n_0),
.B2(n_1),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_161),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_107),
.B(n_40),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_165),
.B(n_193),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_73),
.A2(n_42),
.B1(n_56),
.B2(n_54),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_103),
.A2(n_54),
.B1(n_43),
.B2(n_42),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_62),
.B(n_43),
.Y(n_170)
);

NAND2x1_ASAP7_75t_L g265 ( 
.A(n_170),
.B(n_39),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_83),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_118),
.A2(n_43),
.B1(n_42),
.B2(n_40),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_178),
.A2(n_180),
.B1(n_21),
.B2(n_23),
.Y(n_248)
);

AO22x2_ASAP7_75t_L g180 ( 
.A1(n_99),
.A2(n_57),
.B1(n_51),
.B2(n_44),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_108),
.A2(n_38),
.B1(n_36),
.B2(n_40),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_185),
.A2(n_200),
.B1(n_24),
.B2(n_23),
.Y(n_226)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_109),
.B(n_36),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_110),
.A2(n_38),
.B1(n_41),
.B2(n_39),
.Y(n_200)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_95),
.Y(n_205)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_64),
.B(n_15),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_214),
.B(n_217),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_89),
.B(n_15),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_74),
.B(n_41),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_219),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_88),
.B(n_41),
.Y(n_219)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_222),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_226),
.A2(n_274),
.B(n_265),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_93),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_227),
.Y(n_345)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_228),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_230),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_161),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_231),
.B(n_248),
.Y(n_330)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_136),
.Y(n_233)
);

INVx8_ASAP7_75t_L g352 ( 
.A(n_233),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_178),
.A2(n_78),
.B1(n_77),
.B2(n_80),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_234),
.A2(n_276),
.B1(n_283),
.B2(n_220),
.Y(n_350)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_132),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_154),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_237),
.Y(n_313)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_149),
.Y(n_238)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_238),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_131),
.B(n_21),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_239),
.B(n_253),
.C(n_267),
.Y(n_320)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_149),
.Y(n_240)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_240),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_139),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_241),
.Y(n_324)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_143),
.Y(n_242)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_196),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_244),
.B(n_257),
.Y(n_318)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_246),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_247),
.B(n_250),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_249),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_146),
.Y(n_251)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_176),
.Y(n_252)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_24),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_254),
.Y(n_338)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_255),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_136),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_152),
.A2(n_97),
.B(n_57),
.C(n_39),
.Y(n_261)
);

MAJx3_ASAP7_75t_L g327 ( 
.A(n_261),
.B(n_210),
.C(n_151),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_169),
.B(n_25),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_290),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_185),
.A2(n_91),
.B1(n_87),
.B2(n_84),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_263),
.A2(n_130),
.B1(n_140),
.B2(n_183),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_265),
.Y(n_353)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_270),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_25),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_156),
.A2(n_82),
.B1(n_97),
.B2(n_7),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_268),
.A2(n_272),
.B1(n_275),
.B2(n_291),
.Y(n_333)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_160),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_271),
.B(n_282),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_181),
.A2(n_18),
.B1(n_16),
.B2(n_13),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_207),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_171),
.A2(n_18),
.B1(n_13),
.B2(n_12),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_206),
.A2(n_13),
.B1(n_12),
.B2(n_2),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_198),
.B(n_1),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_281),
.C(n_217),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_166),
.B(n_12),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_279),
.B(n_287),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_169),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_280),
.A2(n_158),
.B1(n_172),
.B2(n_211),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_188),
.B(n_3),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_166),
.B(n_12),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_153),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_155),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_192),
.Y(n_285)
);

INVx13_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_180),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_286),
.B(n_288),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_151),
.B(n_4),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_203),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g289 ( 
.A(n_155),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_289),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_152),
.B(n_4),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_208),
.A2(n_5),
.B1(n_182),
.B2(n_150),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_175),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_292),
.Y(n_344)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_164),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_293),
.A2(n_294),
.B1(n_299),
.B2(n_191),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_162),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_136),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_295),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_215),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_296),
.Y(n_337)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_142),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_297),
.Y(n_354)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_180),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_298),
.B(n_168),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_162),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_305),
.A2(n_238),
.B1(n_240),
.B2(n_233),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_307),
.B(n_335),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_286),
.A2(n_221),
.B1(n_204),
.B2(n_178),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_314),
.A2(n_315),
.B1(n_317),
.B2(n_357),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_172),
.B1(n_158),
.B2(n_134),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_277),
.A2(n_220),
.B1(n_191),
.B2(n_195),
.Y(n_317)
);

OAI22x1_ASAP7_75t_SL g325 ( 
.A1(n_276),
.A2(n_137),
.B1(n_167),
.B2(n_200),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_350),
.B1(n_227),
.B2(n_278),
.Y(n_360)
);

MAJx2_ASAP7_75t_L g388 ( 
.A(n_326),
.B(n_251),
.C(n_273),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_327),
.A2(n_331),
.B(n_340),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_260),
.B(n_174),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_332),
.B(n_336),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_262),
.B(n_177),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_247),
.B(n_148),
.Y(n_336)
);

AOI32xp33_ASAP7_75t_L g340 ( 
.A1(n_290),
.A2(n_225),
.A3(n_245),
.B1(n_223),
.B2(n_231),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_341),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_224),
.A2(n_215),
.B1(n_201),
.B2(n_144),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_342),
.A2(n_355),
.B1(n_229),
.B2(n_273),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_224),
.A2(n_199),
.B1(n_163),
.B2(n_179),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_347),
.A2(n_358),
.B(n_274),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_229),
.A2(n_5),
.B1(n_179),
.B2(n_228),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_248),
.A2(n_5),
.B1(n_179),
.B2(n_280),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_227),
.C(n_255),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_359),
.B(n_368),
.C(n_392),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_360),
.A2(n_358),
.B1(n_353),
.B2(n_320),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_361),
.Y(n_429)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_362),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_363),
.A2(n_300),
.B(n_327),
.Y(n_423)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_350),
.A2(n_235),
.B1(n_248),
.B2(n_278),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_366),
.A2(n_367),
.B1(n_375),
.B2(n_383),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_330),
.A2(n_248),
.B1(n_261),
.B2(n_281),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_256),
.C(n_232),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_281),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_373),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_253),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_308),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_374),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_331),
.A2(n_253),
.B1(n_267),
.B2(n_239),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_308),
.Y(n_379)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_318),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_380),
.B(n_402),
.Y(n_425)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_320),
.B(n_283),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_381),
.B(n_385),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_267),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_393),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_325),
.A2(n_239),
.B1(n_259),
.B2(n_258),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_346),
.Y(n_384)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_322),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_386),
.A2(n_390),
.B1(n_403),
.B2(n_354),
.Y(n_406)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_387),
.B(n_396),
.Y(n_414)
);

XNOR2x1_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_316),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_356),
.A2(n_297),
.B1(n_237),
.B2(n_293),
.Y(n_389)
);

AO21x2_ASAP7_75t_L g441 ( 
.A1(n_389),
.A2(n_311),
.B(n_319),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_314),
.A2(n_246),
.B1(n_242),
.B2(n_236),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_324),
.A2(n_243),
.B1(n_252),
.B2(n_285),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_391),
.A2(n_305),
.B1(n_333),
.B2(n_347),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_335),
.B(n_264),
.Y(n_392)
);

INVx8_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_348),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_398),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_254),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_395),
.B(n_399),
.Y(n_408)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_338),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_397),
.B(n_400),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_332),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_321),
.B(n_292),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_348),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_309),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_404),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_302),
.Y(n_402)
);

OAI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_317),
.A2(n_288),
.B1(n_269),
.B2(n_299),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_309),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_409),
.B1(n_441),
.B2(n_383),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_407),
.A2(n_419),
.B1(n_428),
.B2(n_369),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_324),
.B1(n_327),
.B2(n_353),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_378),
.C(n_359),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_417),
.C(n_440),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_399),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_413),
.B(n_437),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_316),
.C(n_326),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_418),
.A2(n_370),
.B1(n_371),
.B2(n_381),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_360),
.A2(n_307),
.B1(n_327),
.B2(n_300),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_421),
.B(n_436),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_423),
.A2(n_426),
.B(n_439),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_363),
.A2(n_351),
.B(n_343),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_366),
.A2(n_340),
.B1(n_343),
.B2(n_310),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_378),
.B(n_310),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_395),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_365),
.B(n_344),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_365),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_367),
.A2(n_337),
.B(n_323),
.Y(n_439)
);

MAJx2_ASAP7_75t_L g440 ( 
.A(n_381),
.B(n_311),
.C(n_323),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_392),
.B(n_319),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_364),
.C(n_384),
.Y(n_458)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_443),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_465),
.B1(n_466),
.B2(n_477),
.Y(n_478)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_435),
.Y(n_445)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_445),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_423),
.A2(n_373),
.B(n_381),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_446),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_447),
.A2(n_450),
.B1(n_462),
.B2(n_464),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_398),
.Y(n_448)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_448),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_449),
.Y(n_500)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_435),
.Y(n_451)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_451),
.Y(n_506)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_408),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_454),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_428),
.B(n_368),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_453),
.B(n_468),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_414),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_409),
.Y(n_456)
);

OAI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_456),
.A2(n_462),
.B1(n_464),
.B2(n_476),
.Y(n_495)
);

OAI32xp33_ASAP7_75t_L g457 ( 
.A1(n_420),
.A2(n_372),
.A3(n_382),
.B1(n_375),
.B2(n_362),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_463),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_461),
.C(n_469),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_417),
.B(n_372),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_419),
.A2(n_390),
.B1(n_377),
.B2(n_374),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_410),
.A2(n_379),
.B1(n_402),
.B2(n_400),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_434),
.A2(n_385),
.B1(n_387),
.B2(n_397),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_432),
.A2(n_396),
.B1(n_393),
.B2(n_401),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g467 ( 
.A(n_426),
.B(n_404),
.C(n_306),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_467),
.B(n_470),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_408),
.B(n_394),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_412),
.B(n_222),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_427),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_250),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_473),
.C(n_442),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_393),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_472),
.B(n_475),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_230),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_411),
.B(n_344),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_410),
.A2(n_313),
.B1(n_312),
.B2(n_349),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_476),
.A2(n_441),
.B1(n_430),
.B2(n_422),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_434),
.A2(n_313),
.B1(n_284),
.B2(n_294),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_440),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_480),
.B(n_484),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_411),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_455),
.B(n_407),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_485),
.B(n_488),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_463),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_455),
.B(n_420),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_456),
.A2(n_418),
.B1(n_429),
.B2(n_424),
.Y(n_489)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_489),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_447),
.A2(n_429),
.B1(n_441),
.B2(n_406),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_491),
.A2(n_495),
.B1(n_507),
.B2(n_477),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_460),
.B(n_450),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_492),
.B(n_501),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_445),
.A2(n_424),
.B1(n_439),
.B2(n_431),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_496),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_459),
.A2(n_427),
.B(n_430),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_494),
.A2(n_481),
.B(n_508),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_451),
.A2(n_416),
.B1(n_431),
.B2(n_405),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_422),
.C(n_416),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_508),
.C(n_470),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_460),
.B(n_415),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_498),
.B(n_503),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_473),
.B(n_415),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_454),
.B(n_405),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_448),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_446),
.B(n_458),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_459),
.B(n_301),
.C(n_312),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_512),
.B(n_521),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_479),
.B(n_466),
.Y(n_515)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_515),
.Y(n_543)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_496),
.Y(n_516)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_516),
.Y(n_551)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_490),
.Y(n_517)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_517),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_505),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_518),
.B(n_532),
.Y(n_542)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_506),
.Y(n_519)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_519),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_520),
.A2(n_483),
.B1(n_486),
.B2(n_497),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_465),
.C(n_443),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_522),
.B(n_488),
.C(n_487),
.Y(n_545)
);

XNOR2x1_ASAP7_75t_L g526 ( 
.A(n_503),
.B(n_472),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g555 ( 
.A(n_526),
.B(n_536),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_449),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_527),
.B(n_529),
.Y(n_547)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_528),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_509),
.B(n_474),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_510),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_530),
.B(n_531),
.Y(n_560)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_510),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_493),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_499),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_533),
.B(n_303),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_534),
.A2(n_478),
.B1(n_441),
.B2(n_494),
.Y(n_546)
);

OA21x2_ASAP7_75t_L g535 ( 
.A1(n_481),
.A2(n_491),
.B(n_489),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_535),
.A2(n_501),
.B(n_498),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g536 ( 
.A(n_480),
.B(n_492),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_537),
.A2(n_539),
.B(n_511),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_482),
.B(n_457),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_538),
.B(n_539),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_482),
.B(n_441),
.Y(n_539)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_540),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_534),
.A2(n_478),
.B1(n_441),
.B2(n_504),
.Y(n_544)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_544),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_557),
.C(n_558),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_546),
.A2(n_535),
.B1(n_524),
.B2(n_511),
.Y(n_567)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_549),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_525),
.B(n_485),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_550),
.B(n_552),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_525),
.B(n_376),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_528),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_523),
.B(n_301),
.C(n_303),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_523),
.B(n_303),
.C(n_352),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_524),
.A2(n_349),
.B1(n_352),
.B2(n_328),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_559),
.A2(n_551),
.B1(n_548),
.B2(n_553),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_561),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g563 ( 
.A(n_547),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_563),
.B(n_568),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_565),
.A2(n_543),
.B1(n_551),
.B2(n_554),
.Y(n_586)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_567),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_542),
.B(n_529),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_546),
.A2(n_535),
.B1(n_515),
.B2(n_527),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_569),
.B(n_575),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_562),
.B(n_521),
.C(n_513),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_570),
.B(n_573),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_562),
.B(n_513),
.C(n_512),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_522),
.C(n_538),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_576),
.B(n_579),
.C(n_580),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_547),
.B(n_537),
.Y(n_578)
);

CKINVDCx14_ASAP7_75t_R g583 ( 
.A(n_578),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_550),
.B(n_526),
.C(n_536),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_541),
.B(n_514),
.C(n_352),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_560),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_581),
.B(n_556),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g584 ( 
.A1(n_578),
.A2(n_561),
.B(n_543),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_584),
.A2(n_591),
.B(n_596),
.Y(n_608)
);

INVxp33_ASAP7_75t_SL g607 ( 
.A(n_586),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_581),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_594),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_574),
.B(n_552),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_588),
.B(n_579),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_590),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_566),
.A2(n_549),
.B(n_541),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_564),
.B(n_558),
.C(n_557),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_572),
.B(n_556),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_595),
.B(n_597),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_566),
.A2(n_559),
.B(n_553),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_577),
.A2(n_514),
.B1(n_555),
.B2(n_328),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_593),
.B(n_587),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_600),
.B(n_610),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_583),
.A2(n_571),
.B(n_576),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_601),
.B(n_602),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_587),
.A2(n_575),
.B1(n_564),
.B2(n_574),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_604),
.B(n_585),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_584),
.Y(n_605)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_605),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_594),
.B(n_570),
.C(n_573),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_606),
.B(n_609),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_582),
.A2(n_580),
.B1(n_569),
.B2(n_567),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_592),
.B(n_555),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_606),
.B(n_585),
.C(n_582),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_611),
.B(n_618),
.Y(n_626)
);

A2O1A1Ixp33_ASAP7_75t_SL g612 ( 
.A1(n_608),
.A2(n_591),
.B(n_596),
.C(n_589),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_612),
.A2(n_607),
.B(n_609),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_617),
.B(n_619),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_598),
.B(n_590),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_599),
.B(n_589),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_586),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_620),
.B(n_588),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_616),
.A2(n_604),
.B(n_603),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_621),
.A2(n_613),
.B(n_607),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_622),
.A2(n_623),
.B1(n_624),
.B2(n_614),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_616),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_625),
.B(n_615),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_627),
.A2(n_630),
.B(n_329),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_628),
.B(n_629),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_626),
.B(n_612),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_632),
.A2(n_296),
.B1(n_289),
.B2(n_339),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_633),
.B(n_631),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_634),
.B(n_339),
.C(n_289),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_635),
.B(n_339),
.Y(n_636)
);


endmodule