module real_jpeg_26063_n_16 (n_5, n_4, n_8, n_0, n_12, n_359, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_359;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_1),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_1),
.A2(n_69),
.B(n_74),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_1),
.B(n_87),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_1),
.A2(n_131),
.B1(n_155),
.B2(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_1),
.A2(n_33),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_1),
.B(n_60),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_2),
.A2(n_37),
.B1(n_73),
.B2(n_74),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_2),
.A2(n_37),
.B1(n_49),
.B2(n_300),
.Y(n_299)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_5),
.A2(n_73),
.B1(n_74),
.B2(n_119),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_119),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_5),
.A2(n_48),
.B1(n_84),
.B2(n_119),
.Y(n_245)
);

INVx8_ASAP7_75t_SL g56 ( 
.A(n_6),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_7),
.A2(n_47),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_62),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_7),
.A2(n_62),
.B1(n_73),
.B2(n_74),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_62),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_8),
.A2(n_42),
.B1(n_46),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_8),
.A2(n_42),
.B1(n_73),
.B2(n_74),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_9),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_9),
.A2(n_50),
.B1(n_73),
.B2(n_74),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_50),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_11),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_11),
.A2(n_73),
.B1(n_74),
.B2(n_128),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_128),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_11),
.A2(n_58),
.B1(n_84),
.B2(n_128),
.Y(n_257)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_13),
.A2(n_73),
.B1(n_74),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_13),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_136),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_136),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_13),
.A2(n_48),
.B1(n_84),
.B2(n_136),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_15),
.Y(n_134)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_15),
.Y(n_140)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_15),
.Y(n_148)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_15),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_103),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_101),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_90),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_19),
.B(n_90),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_78),
.B2(n_89),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.C(n_65),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_22),
.A2(n_23),
.B1(n_65),
.B2(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_25),
.A2(n_39),
.B(n_239),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_26),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_26),
.A2(n_38),
.B(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_26)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_40)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_27),
.A2(n_29),
.A3(n_33),
.B1(n_174),
.B2(n_183),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_28),
.A2(n_29),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_28),
.B(n_31),
.Y(n_183)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_29),
.A2(n_71),
.B(n_115),
.C(n_121),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_32),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_32),
.A2(n_100),
.B(n_175),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_34),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_33),
.B(n_55),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_34),
.B(n_115),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_34),
.A2(n_54),
.A3(n_63),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_39),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_39),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_39),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_39),
.A2(n_87),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_39),
.A2(n_87),
.B1(n_200),
.B2(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_39),
.A2(n_87),
.B1(n_98),
.B2(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_41),
.B(n_87),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_43),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_53),
.B(n_95),
.Y(n_94)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_49),
.B(n_115),
.Y(n_225)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_49),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_61),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_83),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_51),
.A2(n_60),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_51),
.A2(n_60),
.B1(n_245),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_52),
.A2(n_53),
.B1(n_257),
.B2(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_52),
.A2(n_274),
.B(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_52),
.A2(n_82),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_60),
.B(n_299),
.Y(n_298)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_65),
.A2(n_66),
.B1(n_97),
.B2(n_344),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_94),
.C(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_76),
.B(n_77),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_67),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_67),
.A2(n_76),
.B1(n_118),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_67),
.A2(n_76),
.B1(n_127),
.B2(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_67),
.A2(n_77),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_67),
.B(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_72),
.B(n_115),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_72),
.B(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_72),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_72),
.A2(n_116),
.B1(n_263),
.B2(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_73),
.B(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_76),
.B(n_77),
.Y(n_215)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_84),
.A2(n_115),
.B(n_225),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.C(n_96),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_342),
.Y(n_349)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_94),
.A2(n_342),
.B1(n_343),
.B2(n_345),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_94),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_96),
.B(n_349),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_97),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI321xp33_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_339),
.A3(n_350),
.B1(n_355),
.B2(n_356),
.C(n_359),
.Y(n_103)
);

AOI311xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_290),
.A3(n_329),
.B(n_333),
.C(n_334),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_247),
.C(n_285),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_219),
.B(n_246),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_193),
.B(n_218),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_167),
.B(n_192),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_141),
.B(n_166),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_122),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_111),
.B(n_122),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_120),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_113),
.B1(n_120),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_140),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_116),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_116),
.A2(n_280),
.B(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_120),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_129),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_129),
.C(n_130),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_135),
.B(n_137),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_145),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_131),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_131),
.A2(n_186),
.B(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_131),
.A2(n_156),
.B(n_185),
.Y(n_305)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_132),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_132),
.B(n_189),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_132),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_227)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_137),
.B(n_209),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_151),
.B(n_165),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_149),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_149),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_159),
.B(n_164),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_154),
.Y(n_164)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_169),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_181),
.B1(n_190),
.B2(n_191),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_170)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_180),
.C(n_190),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_184),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_194),
.B(n_195),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_210),
.B2(n_211),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_213),
.C(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_203),
.C(n_204),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_208),
.B(n_209),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_216),
.B2(n_217),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_215),
.B(n_264),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_220),
.B(n_221),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_236),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_222)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_223),
.B(n_235),
.C(n_236),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_227),
.B1(n_231),
.B2(n_232),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_231),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_227),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_243),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_240),
.C(n_243),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g335 ( 
.A1(n_248),
.A2(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_266),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_249),
.B(n_266),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_258),
.C(n_259),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_251),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_254),
.C(n_255),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_258),
.B(n_259),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_262),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_277),
.B2(n_281),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_268),
.B(n_281),
.C(n_284),
.Y(n_331)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_276),
.Y(n_269)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_275),
.C(n_276),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_277),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_279),
.Y(n_295)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_282),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_287),
.Y(n_336)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

O2A1O1Ixp33_ASAP7_75t_SL g334 ( 
.A1(n_291),
.A2(n_330),
.B(n_335),
.C(n_338),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_311),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_311),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_304),
.C(n_310),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g332 ( 
.A(n_293),
.B(n_304),
.CI(n_310),
.CON(n_332),
.SN(n_332)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_303),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_297),
.C(n_301),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_301),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_299),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_302),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_309),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_305),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_307),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_309),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_309),
.A2(n_319),
.B(n_323),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_328),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_318),
.B1(n_326),
.B2(n_327),
.Y(n_312)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_316),
.B(n_317),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_314),
.B(n_316),
.Y(n_317)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_317),
.A2(n_341),
.B1(n_346),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_326),
.C(n_328),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_321),
.B2(n_325),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_331),
.B(n_332),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g358 ( 
.A(n_332),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_348),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_340),
.B(n_348),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_346),
.C(n_347),
.Y(n_340)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_343),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_347),
.B(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_351),
.B(n_352),
.Y(n_355)
);


endmodule