module fake_jpeg_12962_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_1),
.B(n_25),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_23),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_56),
.B1(n_45),
.B2(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_3),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_47),
.Y(n_73)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_4),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_46),
.B1(n_56),
.B2(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_77),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_51),
.B(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_57),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_82),
.C(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_58),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_57),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_42),
.A3(n_43),
.B1(n_55),
.B2(n_37),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_87),
.Y(n_100)
);

A2O1A1O1Ixp25_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_54),
.B(n_76),
.C(n_75),
.D(n_70),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_91),
.B(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_95),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_98),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_40),
.C(n_21),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_8),
.C(n_9),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_6),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_9),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_13),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_16),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_109)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_36),
.B(n_33),
.Y(n_115)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_28),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_32),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_126),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_101),
.B1(n_100),
.B2(n_110),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_117),
.C(n_120),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_129),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_101),
.C(n_118),
.Y(n_129)
);

OAI21x1_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_128),
.B(n_126),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_131),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_115),
.Y(n_134)
);


endmodule