module fake_jpeg_31023_n_341 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_341);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_53),
.Y(n_83)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_56),
.Y(n_102)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_60),
.Y(n_109)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_67),
.Y(n_110)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_66),
.Y(n_100)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_74),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_76),
.A2(n_86),
.B1(n_88),
.B2(n_93),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_41),
.B1(n_38),
.B2(n_20),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_77),
.A2(n_94),
.B1(n_106),
.B2(n_14),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_78),
.B(n_85),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_26),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_82),
.B(n_17),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_38),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_28),
.B1(n_31),
.B2(n_30),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_29),
.B1(n_34),
.B2(n_39),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_8),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_31),
.B1(n_28),
.B2(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_34),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_29),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_30),
.B1(n_22),
.B2(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_30),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_101),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_59),
.A2(n_43),
.B1(n_37),
.B2(n_35),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_105),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_35),
.B1(n_32),
.B2(n_24),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_37),
.B1(n_32),
.B2(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_23),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_23),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_104),
.B(n_107),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_37),
.B1(n_2),
.B2(n_4),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_45),
.A2(n_42),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_1),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_63),
.A2(n_1),
.B1(n_4),
.B2(n_7),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_8),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_14),
.C(n_16),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_123),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_115),
.A2(n_106),
.B1(n_151),
.B2(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_79),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_11),
.B(n_12),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_71),
.Y(n_123)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_132),
.Y(n_154)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_77),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_151),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_13),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_134),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_139),
.B1(n_108),
.B2(n_80),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_148),
.B1(n_18),
.B2(n_80),
.Y(n_186)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_18),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_78),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_150),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_85),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_157),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_112),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_107),
.B(n_74),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_158),
.A2(n_177),
.B(n_119),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_161),
.B(n_183),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_110),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_137),
.B1(n_143),
.B2(n_148),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_90),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_175),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_95),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_94),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_113),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_100),
.B(n_113),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_100),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_188),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_100),
.C(n_86),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_133),
.C(n_129),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_93),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_142),
.B1(n_139),
.B2(n_131),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_91),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_114),
.B(n_118),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_189),
.A2(n_162),
.B(n_174),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_158),
.B(n_125),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_200),
.C(n_206),
.Y(n_221)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

BUFx24_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_131),
.B(n_118),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_193),
.A2(n_205),
.B1(n_210),
.B2(n_169),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_142),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_194),
.B(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_198),
.A2(n_201),
.B1(n_203),
.B2(n_197),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_199),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_131),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_128),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_89),
.B1(n_117),
.B2(n_121),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_212),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_141),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_185),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_217),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_171),
.C(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_162),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_166),
.B(n_134),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_116),
.Y(n_223)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_170),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_224),
.B(n_188),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_225),
.B(n_231),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_162),
.B1(n_168),
.B2(n_164),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_190),
.C(n_214),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_216),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_153),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_242),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_243),
.B(n_246),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_164),
.B(n_177),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_245),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_164),
.B(n_178),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_199),
.B1(n_205),
.B2(n_206),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_249),
.B(n_262),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_256),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_270),
.B1(n_248),
.B2(n_238),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_216),
.C(n_197),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_258),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_201),
.C(n_199),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_241),
.C(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_267),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_165),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_263),
.B(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_165),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_266),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_198),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_217),
.C(n_161),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_248),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_210),
.B1(n_215),
.B2(n_218),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_239),
.B(n_230),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_278),
.B(n_284),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_231),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_276),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_239),
.Y(n_277)
);

OAI21x1_ASAP7_75t_SL g295 ( 
.A1(n_277),
.A2(n_278),
.B(n_272),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_250),
.A2(n_246),
.B1(n_236),
.B2(n_227),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_281),
.B(n_282),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_189),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_250),
.A2(n_227),
.B(n_242),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_269),
.B1(n_270),
.B2(n_253),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_255),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_298),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_296),
.B1(n_300),
.B2(n_303),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_287),
.B(n_258),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_261),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_267),
.B(n_251),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_285),
.Y(n_308)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_275),
.C(n_273),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_307),
.B(n_309),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_310),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_275),
.C(n_285),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_288),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_288),
.C(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_314),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_226),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_238),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_298),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_300),
.B1(n_292),
.B2(n_290),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_316),
.A2(n_322),
.B1(n_306),
.B2(n_308),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_292),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_319),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_303),
.B(n_235),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_324),
.B(n_235),
.Y(n_326)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_226),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_326),
.Y(n_335)
);

OAI321xp33_ASAP7_75t_L g327 ( 
.A1(n_317),
.A2(n_306),
.A3(n_234),
.B1(n_312),
.B2(n_229),
.C(n_209),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_327),
.A2(n_328),
.B1(n_169),
.B2(n_173),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_234),
.B1(n_229),
.B2(n_204),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_187),
.C(n_185),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_155),
.C(n_124),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_320),
.A2(n_179),
.B(n_172),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_318),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_330),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_336),
.B(n_334),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_338),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_337),
.B(n_331),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_339),
.Y(n_341)
);


endmodule