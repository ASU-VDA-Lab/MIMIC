module fake_jpeg_26667_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_1),
.B(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_49),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_33),
.B1(n_20),
.B2(n_28),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_54),
.B1(n_56),
.B2(n_22),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_48),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_64),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_55),
.Y(n_82)
);

NAND2xp67_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_21),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_21),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_33),
.B1(n_20),
.B2(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_33),
.B1(n_22),
.B2(n_26),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_39),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_39),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_79),
.B1(n_62),
.B2(n_52),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_39),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_68),
.Y(n_117)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_69),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_76),
.Y(n_99)
);

INVxp33_ASAP7_75t_SL g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_74),
.B(n_91),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_86),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_49),
.B(n_50),
.C(n_58),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_66),
.B(n_68),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_55),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_43),
.B1(n_34),
.B2(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_88),
.B1(n_87),
.B2(n_65),
.Y(n_139)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_39),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_66),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_67),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_62),
.B1(n_60),
.B2(n_19),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_106),
.A2(n_76),
.B1(n_65),
.B2(n_58),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_81),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_120),
.C(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_59),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_59),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_92),
.B1(n_77),
.B2(n_52),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_85),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_122),
.B(n_143),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_132),
.B(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_78),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_133),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_111),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_80),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_80),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_141),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_85),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_138),
.Y(n_157)
);

AO21x2_ASAP7_75t_SL g137 ( 
.A1(n_104),
.A2(n_117),
.B(n_120),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_117),
.B(n_102),
.C(n_120),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_69),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_105),
.B1(n_112),
.B2(n_114),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_84),
.Y(n_145)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_48),
.Y(n_146)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_148),
.A2(n_112),
.B1(n_105),
.B2(n_103),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_58),
.C(n_52),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_102),
.C(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_158),
.B1(n_150),
.B2(n_144),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_176),
.B1(n_177),
.B2(n_121),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_111),
.B1(n_113),
.B2(n_104),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_170),
.C(n_179),
.Y(n_185)
);

CKINVDCx10_ASAP7_75t_R g162 ( 
.A(n_147),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_168),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_169),
.B(n_172),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_167),
.B(n_17),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_137),
.B(n_132),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_117),
.C(n_103),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_40),
.B(n_116),
.C(n_16),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_101),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_173),
.B(n_174),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_35),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_137),
.B1(n_148),
.B2(n_124),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_114),
.B1(n_98),
.B2(n_93),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_98),
.C(n_93),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_126),
.B(n_89),
.C(n_35),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_127),
.C(n_89),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_118),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_121),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_19),
.B(n_24),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_131),
.B(n_130),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_190),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_166),
.B(n_138),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_189),
.B(n_151),
.Y(n_219)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_198),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_149),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_196),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_123),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_202),
.B1(n_204),
.B2(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_206),
.B(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_169),
.A2(n_127),
.B1(n_139),
.B2(n_122),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_160),
.C(n_180),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_135),
.B1(n_19),
.B2(n_24),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_156),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_205),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_173),
.B(n_165),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_177),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_17),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_161),
.A2(n_0),
.B(n_1),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_29),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_174),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_191),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_223),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_218),
.B1(n_228),
.B2(n_188),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_164),
.B1(n_178),
.B2(n_162),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_219),
.B(n_220),
.Y(n_255)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_233),
.C(n_203),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_231),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_183),
.B1(n_179),
.B2(n_151),
.Y(n_228)
);

NOR4xp25_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_172),
.C(n_157),
.D(n_21),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_229),
.B(n_232),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_191),
.B(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_185),
.B(n_157),
.C(n_21),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_31),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_234),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_188),
.B(n_25),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_13),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_240),
.C(n_247),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_215),
.C(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_251),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_217),
.A2(n_206),
.B1(n_189),
.B2(n_195),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_194),
.C(n_196),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_212),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_250),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_212),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_210),
.C(n_192),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_236),
.C(n_222),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_195),
.B(n_186),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_221),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_232),
.A2(n_224),
.B1(n_214),
.B2(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_256),
.B(n_258),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_31),
.B1(n_25),
.B2(n_27),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_219),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_268),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_252),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_269),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_216),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_216),
.Y(n_269)
);

FAx1_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_213),
.CI(n_223),
.CON(n_270),
.SN(n_270)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_254),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_222),
.C(n_235),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_255),
.C(n_238),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_271),
.Y(n_296)
);

AOI221xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_246),
.B1(n_236),
.B2(n_242),
.C(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_255),
.CI(n_250),
.CON(n_278),
.SN(n_278)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_283),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_281),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_266),
.B1(n_274),
.B2(n_260),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_249),
.C(n_251),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_264),
.C(n_271),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_27),
.B1(n_10),
.B2(n_15),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_6),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_27),
.B1(n_12),
.B2(n_9),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_11),
.B1(n_14),
.B2(n_12),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_290),
.A2(n_292),
.B1(n_299),
.B2(n_1),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_276),
.A2(n_280),
.B1(n_278),
.B2(n_282),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_285),
.B(n_284),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_9),
.B(n_29),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_281),
.C(n_278),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_297),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_7),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_6),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_1),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_27),
.C(n_32),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_32),
.C(n_29),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_306),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_295),
.C(n_296),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_305),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_29),
.A3(n_6),
.B1(n_14),
.B2(n_9),
.C1(n_32),
.C2(n_5),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_32),
.C(n_29),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_307),
.A2(n_308),
.B(n_2),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_32),
.B(n_2),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_300),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_292),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_316),
.B(n_302),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_313),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_5),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_2),
.C(n_3),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_315),
.B1(n_310),
.B2(n_5),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_3),
.B(n_4),
.Y(n_322)
);

OAI321xp33_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_3),
.A3(n_4),
.B1(n_317),
.B2(n_320),
.C(n_302),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_3),
.Y(n_324)
);


endmodule