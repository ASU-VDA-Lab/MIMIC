module fake_jpeg_17954_n_207 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_207);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_0),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_24),
.Y(n_50)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_27),
.B1(n_31),
.B2(n_24),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_53),
.B1(n_56),
.B2(n_23),
.Y(n_74)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_15),
.B1(n_21),
.B2(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_62),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_15),
.B1(n_19),
.B2(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_25),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_30),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_34),
.B1(n_33),
.B2(n_29),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_29),
.B1(n_23),
.B2(n_20),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_74),
.B1(n_20),
.B2(n_28),
.Y(n_103)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_42),
.B1(n_41),
.B2(n_36),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_45),
.B1(n_52),
.B2(n_42),
.Y(n_85)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_83),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_103),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_71),
.Y(n_106)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_30),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_38),
.A3(n_30),
.B1(n_69),
.B2(n_40),
.C1(n_65),
.C2(n_43),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_100),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_82),
.Y(n_124)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_41),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_82),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_123),
.Y(n_142)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_87),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_116),
.B(n_95),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_90),
.C(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_98),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_18),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_122),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_75),
.B1(n_78),
.B2(n_76),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_125),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_103),
.B1(n_100),
.B2(n_88),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_113),
.B1(n_18),
.B2(n_22),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_85),
.B(n_84),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_140),
.B(n_117),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_141),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_99),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_56),
.B(n_66),
.C(n_43),
.D(n_55),
.Y(n_144)
);

OA21x2_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_127),
.B(n_129),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_72),
.C(n_44),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_114),
.C(n_115),
.Y(n_148)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_156),
.C(n_142),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_149),
.C(n_150),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_106),
.C(n_110),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_122),
.C(n_118),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_125),
.C(n_117),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_158),
.C(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_126),
.C(n_107),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_141),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_126),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_144),
.B1(n_143),
.B2(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_171),
.C(n_22),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_160),
.Y(n_178)
);

BUFx12_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_143),
.C(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_133),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_170),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_149),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_180),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_150),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_16),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_183),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_175),
.A2(n_169),
.B1(n_171),
.B2(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_185),
.B(n_192),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_184),
.A2(n_162),
.B(n_165),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_187),
.B(n_9),
.Y(n_193)
);

AOI21x1_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_170),
.B(n_3),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_8),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_9),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_5),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_181),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_193),
.A2(n_197),
.B1(n_7),
.B2(n_12),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_11),
.C(n_14),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_196),
.A2(n_190),
.B(n_189),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_189),
.B(n_4),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_0),
.B(n_4),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_204),
.B(n_0),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_201),
.Y(n_204)
);

OAI31xp33_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_202),
.A3(n_12),
.B(n_16),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_16),
.Y(n_207)
);


endmodule