module fake_jpeg_30904_n_539 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_539);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_539;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_10),
.B(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_38),
.B(n_0),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_68),
.B(n_84),
.Y(n_126)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_81),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_44),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g153 ( 
.A(n_80),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_37),
.B(n_1),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx11_ASAP7_75t_SL g83 ( 
.A(n_21),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_21),
.B(n_1),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_37),
.B(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_95),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_20),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx16f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g145 ( 
.A(n_97),
.Y(n_145)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_100),
.B(n_102),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_20),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_105),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_114),
.B(n_123),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_25),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_115),
.B(n_149),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_120),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_33),
.B1(n_42),
.B2(n_53),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_121),
.A2(n_122),
.B1(n_26),
.B2(n_46),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_58),
.A2(n_24),
.B1(n_29),
.B2(n_50),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_24),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_41),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_124),
.B(n_29),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_132),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_40),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_134),
.B(n_154),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_47),
.B(n_51),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_68),
.A2(n_34),
.B(n_45),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_82),
.B(n_41),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_54),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

INVx2_ASAP7_75t_R g162 ( 
.A(n_104),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_57),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_168),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_115),
.A2(n_47),
.B1(n_48),
.B2(n_22),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_169),
.B(n_204),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_50),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_171),
.B(n_172),
.Y(n_230)
);

INVx4_ASAP7_75t_SL g172 ( 
.A(n_162),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_167),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_180),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_121),
.A2(n_33),
.B1(n_55),
.B2(n_66),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_174),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_116),
.A2(n_33),
.B1(n_98),
.B2(n_70),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_175),
.Y(n_236)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_46),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_126),
.B(n_26),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_201),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_183),
.A2(n_186),
.B1(n_214),
.B2(n_85),
.Y(n_235)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_126),
.A2(n_92),
.B1(n_101),
.B2(n_62),
.Y(n_186)
);

CKINVDCx12_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_187),
.B(n_188),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_30),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_109),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_191),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_132),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_192),
.B(n_198),
.Y(n_252)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_150),
.Y(n_194)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_26),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_140),
.B(n_31),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_135),
.B(n_30),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_205),
.B(n_206),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_31),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_135),
.B(n_40),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_208),
.B(n_209),
.Y(n_262)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_107),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_210),
.B(n_217),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_113),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_211),
.A2(n_164),
.B1(n_165),
.B2(n_127),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_147),
.B(n_48),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_213),
.Y(n_237)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_127),
.A2(n_103),
.B1(n_65),
.B2(n_93),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_106),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_215),
.B(n_156),
.Y(n_251)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_218),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_142),
.B(n_51),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_79),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_220),
.Y(n_245)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_159),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_45),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_168),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_78),
.B1(n_72),
.B2(n_73),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_232),
.A2(n_243),
.B1(n_246),
.B2(n_263),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_235),
.A2(n_191),
.B1(n_143),
.B2(n_214),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_179),
.A2(n_142),
.B(n_130),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_250),
.B(n_254),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_179),
.A2(n_152),
.B1(n_136),
.B2(n_165),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_242),
.A2(n_253),
.B1(n_191),
.B2(n_181),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_136),
.B1(n_152),
.B2(n_129),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_219),
.A2(n_129),
.B1(n_164),
.B2(n_113),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_168),
.A2(n_130),
.B(n_69),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_251),
.B(n_257),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_172),
.A2(n_155),
.B1(n_141),
.B2(n_108),
.Y(n_253)
);

NAND2x1_ASAP7_75t_L g254 ( 
.A(n_182),
.B(n_45),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_77),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_207),
.B(n_20),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_265),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_178),
.A2(n_87),
.B1(n_91),
.B2(n_157),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_176),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_282),
.Y(n_316)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_224),
.B(n_201),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_271),
.B(n_280),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

INVx3_ASAP7_75t_SL g320 ( 
.A(n_272),
.Y(n_320)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_177),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_274),
.B(n_296),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_221),
.C(n_185),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_276),
.B(n_251),
.C(n_230),
.Y(n_329)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_224),
.B(n_212),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_281),
.A2(n_286),
.B1(n_291),
.B2(n_293),
.Y(n_305)
);

OAI32xp33_ASAP7_75t_L g282 ( 
.A1(n_234),
.A2(n_186),
.A3(n_169),
.B1(n_184),
.B2(n_218),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_244),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_283),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_243),
.A2(n_264),
.B1(n_236),
.B2(n_232),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_285),
.A2(n_299),
.B1(n_303),
.B2(n_242),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_235),
.A2(n_157),
.B1(n_216),
.B2(n_209),
.Y(n_286)
);

AO22x2_ASAP7_75t_L g287 ( 
.A1(n_236),
.A2(n_215),
.B1(n_204),
.B2(n_193),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_302),
.Y(n_334)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_SL g289 ( 
.A(n_227),
.B(n_45),
.C(n_197),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_300),
.B(n_250),
.Y(n_309)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_264),
.A2(n_199),
.B1(n_221),
.B2(n_211),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_225),
.B(n_190),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_227),
.B(n_90),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_298),
.Y(n_325)
);

BUFx4f_ASAP7_75t_SL g298 ( 
.A(n_229),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_246),
.A2(n_220),
.B1(n_170),
.B2(n_195),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_227),
.A2(n_203),
.B(n_181),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_244),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_301),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_234),
.A2(n_170),
.B1(n_200),
.B2(n_128),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_255),
.A2(n_189),
.B1(n_194),
.B2(n_128),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_260),
.Y(n_304)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_237),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_328),
.C(n_329),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_309),
.B(n_223),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_279),
.B(n_237),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_312),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_289),
.A2(n_259),
.B1(n_233),
.B2(n_260),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_311),
.A2(n_272),
.B1(n_223),
.B2(n_238),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_258),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_SL g314 ( 
.A1(n_284),
.A2(n_257),
.B(n_245),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_336),
.B1(n_337),
.B2(n_287),
.Y(n_353)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_262),
.B(n_249),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_293),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_270),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_318),
.B(n_322),
.Y(n_354)
);

XNOR2x2_ASAP7_75t_L g321 ( 
.A(n_267),
.B(n_254),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_321),
.A2(n_332),
.B1(n_286),
.B2(n_302),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_230),
.B(n_256),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_327),
.A2(n_309),
.B(n_317),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_282),
.B(n_245),
.Y(n_328)
);

OAI32xp33_ASAP7_75t_L g335 ( 
.A1(n_280),
.A2(n_263),
.A3(n_254),
.B1(n_261),
.B2(n_240),
.Y(n_335)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_335),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_275),
.A2(n_266),
.B1(n_241),
.B2(n_226),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_275),
.A2(n_285),
.B1(n_301),
.B2(n_283),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_261),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_340),
.B(n_346),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_322),
.Y(n_341)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_344),
.A2(n_353),
.B1(n_355),
.B2(n_361),
.Y(n_400)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_307),
.Y(n_345)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_345),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_271),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_334),
.A2(n_278),
.B1(n_299),
.B2(n_294),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_347),
.A2(n_370),
.B1(n_324),
.B2(n_338),
.Y(n_386)
);

AO21x1_ASAP7_75t_L g385 ( 
.A1(n_348),
.A2(n_368),
.B(n_372),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_297),
.B(n_287),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_350),
.Y(n_379)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_351),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_354),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_337),
.A2(n_328),
.B1(n_332),
.B2(n_336),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_333),
.B(n_273),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_356),
.B(n_359),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_317),
.A2(n_294),
.B1(n_287),
.B2(n_288),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_357),
.A2(n_366),
.B1(n_369),
.B2(n_326),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_292),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_329),
.C(n_312),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_325),
.B(n_287),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_362),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_305),
.A2(n_277),
.B1(n_272),
.B2(n_269),
.Y(n_361)
);

AND2x6_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_327),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_310),
.B(n_228),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_363),
.B(n_367),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_334),
.A2(n_304),
.B(n_266),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_364),
.Y(n_398)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_305),
.A2(n_266),
.B1(n_268),
.B2(n_298),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_315),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_323),
.A2(n_241),
.B1(n_238),
.B2(n_228),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_323),
.B(n_226),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_371),
.B(n_331),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_96),
.Y(n_372)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_375),
.B(n_377),
.Y(n_412)
);

OAI22x1_ASAP7_75t_L g376 ( 
.A1(n_357),
.A2(n_298),
.B1(n_326),
.B2(n_313),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_376),
.A2(n_366),
.B(n_372),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_331),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_383),
.A2(n_391),
.B1(n_376),
.B2(n_364),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_386),
.A2(n_390),
.B1(n_397),
.B2(n_403),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_338),
.C(n_313),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_343),
.C(n_358),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_342),
.A2(n_320),
.B1(n_339),
.B2(n_306),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_344),
.A2(n_320),
.B1(n_306),
.B2(n_339),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_295),
.Y(n_392)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_203),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_394),
.B(n_396),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_320),
.Y(n_395)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_395),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_359),
.B(n_196),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_348),
.A2(n_206),
.B1(n_67),
.B2(n_60),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_352),
.B(n_45),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_371),
.Y(n_413)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_345),
.Y(n_402)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_402),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_348),
.A2(n_145),
.B1(n_18),
.B2(n_53),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_349),
.Y(n_404)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_404),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_379),
.A2(n_360),
.B(n_350),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_405),
.B(n_430),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_406),
.B(n_416),
.C(n_424),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_408),
.A2(n_411),
.B1(n_431),
.B2(n_397),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_391),
.A2(n_347),
.B1(n_355),
.B2(n_362),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_423),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_353),
.C(n_367),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_365),
.Y(n_417)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_417),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_395),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_420),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_387),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_351),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_429),
.Y(n_447)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_422),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_375),
.B(n_368),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_361),
.C(n_372),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_387),
.B(n_370),
.Y(n_426)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_426),
.Y(n_443)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_374),
.Y(n_427)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_427),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_374),
.B(n_2),
.Y(n_428)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_2),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_400),
.A2(n_145),
.B1(n_3),
.B2(n_4),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_432),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_20),
.C(n_117),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_380),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_434),
.A2(n_453),
.B1(n_455),
.B2(n_425),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_411),
.A2(n_382),
.B1(n_419),
.B2(n_408),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_435),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_404),
.C(n_379),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_449),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_414),
.B(n_388),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_437),
.B(n_456),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_431),
.A2(n_386),
.B1(n_390),
.B2(n_403),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_445),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_426),
.A2(n_398),
.B1(n_401),
.B2(n_384),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_409),
.A2(n_398),
.B1(n_400),
.B2(n_385),
.Y(n_448)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_448),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_416),
.B(n_385),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_L g453 ( 
.A1(n_427),
.A2(n_385),
.B1(n_373),
.B2(n_402),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_405),
.A2(n_401),
.B(n_384),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_454),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_415),
.A2(n_380),
.B1(n_18),
.B2(n_4),
.Y(n_455)
);

NOR3xp33_ASAP7_75t_L g457 ( 
.A(n_452),
.B(n_442),
.C(n_439),
.Y(n_457)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_457),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_439),
.A2(n_407),
.B(n_432),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_458),
.B(n_467),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_443),
.A2(n_430),
.B1(n_415),
.B2(n_407),
.Y(n_459)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_459),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_423),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_460),
.B(n_438),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_425),
.Y(n_463)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_463),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_464),
.A2(n_463),
.B1(n_472),
.B2(n_471),
.Y(n_476)
);

BUFx12f_ASAP7_75t_SL g465 ( 
.A(n_436),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_465),
.A2(n_450),
.B(n_444),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_443),
.A2(n_424),
.B1(n_428),
.B2(n_410),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_474),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_440),
.A2(n_422),
.B(n_410),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_412),
.C(n_413),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_470),
.C(n_475),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_412),
.C(n_433),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_446),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_43),
.C(n_117),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_476),
.A2(n_463),
.B1(n_472),
.B2(n_459),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_467),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_483),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_478),
.B(n_484),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_454),
.C(n_440),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_480),
.B(n_482),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_461),
.C(n_460),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_447),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_448),
.C(n_434),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_487),
.A2(n_464),
.B(n_475),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_465),
.A2(n_444),
.B(n_450),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_488),
.A2(n_458),
.B(n_474),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_455),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_53),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_473),
.B(n_446),
.Y(n_491)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_491),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_492),
.Y(n_493)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_493),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_495),
.A2(n_489),
.B1(n_479),
.B2(n_478),
.Y(n_508)
);

AOI21x1_ASAP7_75t_L g513 ( 
.A1(n_496),
.A2(n_497),
.B(n_493),
.Y(n_513)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_488),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_501),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_507),
.Y(n_511)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_481),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_504),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_482),
.A2(n_120),
.B(n_3),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_503),
.A2(n_5),
.B(n_6),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_487),
.A2(n_485),
.B1(n_490),
.B2(n_480),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_8),
.Y(n_519)
);

MAJx2_ASAP7_75t_L g507 ( 
.A(n_479),
.B(n_2),
.C(n_3),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_515),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_513),
.A2(n_496),
.B(n_495),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_120),
.C(n_18),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_516),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_494),
.B(n_4),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_500),
.B(n_4),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_518),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_500),
.B(n_6),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_519),
.A2(n_507),
.B1(n_10),
.B2(n_11),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_522),
.A2(n_525),
.B(n_511),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_526),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_509),
.A2(n_9),
.B(n_11),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_12),
.C(n_13),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_520),
.A2(n_512),
.B(n_514),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_527),
.A2(n_528),
.B(n_12),
.Y(n_532)
);

OAI31xp33_ASAP7_75t_SL g528 ( 
.A1(n_523),
.A2(n_508),
.A3(n_511),
.B(n_517),
.Y(n_528)
);

AOI322xp5_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_521),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.C1(n_17),
.C2(n_12),
.Y(n_531)
);

AOI21x1_ASAP7_75t_SL g535 ( 
.A1(n_531),
.A2(n_532),
.B(n_533),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_530),
.B(n_14),
.Y(n_533)
);

OAI31xp33_ASAP7_75t_SL g534 ( 
.A1(n_532),
.A2(n_14),
.A3(n_16),
.B(n_43),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_534),
.A2(n_14),
.B(n_16),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_535),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_43),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_43),
.Y(n_539)
);


endmodule