module fake_netlist_5_2134_n_1742 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1742);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1742;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1543;
wire n_1399;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_81),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_21),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_89),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_123),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_16),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_84),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_53),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_108),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_67),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_90),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_88),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_59),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_46),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_127),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_37),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_86),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_82),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_12),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_25),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_53),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_121),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_150),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_1),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_76),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_130),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_48),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_122),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_3),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_26),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_26),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_35),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_97),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_129),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_38),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_91),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_87),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_69),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_66),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_32),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_95),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_124),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_58),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_8),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_114),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_142),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_107),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_35),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_27),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_5),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_85),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_40),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_33),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_65),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_21),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_19),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_110),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_40),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_120),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_75),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_93),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_38),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_20),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_113),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_20),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_94),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_28),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_30),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_16),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_68),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_24),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_48),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_139),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_55),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_80),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_137),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_52),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_6),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_59),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_103),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_12),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_112),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_55),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_30),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_46),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_54),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_7),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_154),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_78),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_101),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_138),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_15),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_98),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_2),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_71),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_29),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_39),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_43),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_9),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_1),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_58),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_79),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_47),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_153),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_73),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_29),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_106),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_36),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_105),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_44),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_56),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_2),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_15),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_28),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_56),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_126),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_13),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_118),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_34),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_102),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_42),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_14),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_52),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_49),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_4),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_54),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_51),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_152),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_60),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_99),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_24),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_13),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_141),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_100),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_33),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_41),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_155),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_44),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_42),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_60),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_158),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_161),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_269),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_211),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_269),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_269),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_269),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_230),
.B(n_0),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_277),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_174),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_162),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_298),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_164),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_165),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_180),
.Y(n_331)
);

BUFx2_ASAP7_75t_SL g332 ( 
.A(n_198),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_166),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_168),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_169),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_170),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_171),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_272),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_160),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g341 ( 
.A(n_198),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_174),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_207),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_207),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_272),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_272),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_198),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_272),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_248),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_163),
.B(n_0),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_182),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_160),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_175),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_179),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_230),
.B(n_3),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_248),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_183),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_311),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_311),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_184),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_248),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_163),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_163),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_231),
.B(n_4),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_172),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_163),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_192),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_192),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_186),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_194),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_185),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_189),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_194),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_191),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_228),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_193),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_228),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_199),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_202),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_276),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_203),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_231),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_317),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_368),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_339),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_339),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_325),
.B(n_280),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_344),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

OA21x2_ASAP7_75t_L g401 ( 
.A1(n_368),
.A2(n_306),
.B(n_276),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_279),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_351),
.B(n_299),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_325),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_319),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_369),
.B(n_279),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_320),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_347),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_347),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_320),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_370),
.B(n_227),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_349),
.B(n_279),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_327),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_351),
.B(n_361),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_348),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_329),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_348),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_328),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_328),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_177),
.Y(n_425)
);

AND2x2_ASAP7_75t_SL g426 ( 
.A(n_321),
.B(n_177),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_361),
.B(n_210),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_330),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_361),
.B(n_212),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_352),
.Y(n_433)
);

NOR3xp33_ASAP7_75t_L g434 ( 
.A(n_359),
.B(n_173),
.C(n_172),
.Y(n_434)
);

AND2x2_ASAP7_75t_SL g435 ( 
.A(n_353),
.B(n_157),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_352),
.Y(n_436)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_333),
.A2(n_167),
.B(n_157),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_333),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_358),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_372),
.B(n_214),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_357),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_360),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_360),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_366),
.B(n_216),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_362),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_316),
.A2(n_302),
.B1(n_297),
.B2(n_288),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_372),
.B(n_167),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_354),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_366),
.B(n_178),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_364),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_367),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_366),
.B(n_219),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_439),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_401),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_390),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_388),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

INVx8_ASAP7_75t_L g465 ( 
.A(n_453),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_SL g466 ( 
.A(n_452),
.B(n_323),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_418),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_393),
.B(n_332),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_401),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_388),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_401),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_401),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_415),
.B(n_312),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_415),
.B(n_314),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_426),
.B(n_324),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_393),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_391),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_418),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_414),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_426),
.B(n_326),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_435),
.A2(n_353),
.B1(n_306),
.B2(n_214),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_426),
.B(n_334),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_414),
.Y(n_491)
);

NOR3xp33_ASAP7_75t_L g492 ( 
.A(n_450),
.B(n_375),
.C(n_355),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_452),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_404),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_439),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_402),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_435),
.B(n_335),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_392),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_389),
.B(n_332),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_420),
.B(n_331),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_404),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_446),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_435),
.B(n_336),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_446),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_404),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_426),
.B(n_337),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_420),
.B(n_338),
.Y(n_509)
);

NOR3xp33_ASAP7_75t_L g510 ( 
.A(n_450),
.B(n_371),
.C(n_340),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_416),
.B(n_341),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_414),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_389),
.B(n_341),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_435),
.A2(n_434),
.B1(n_396),
.B2(n_236),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_414),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_402),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_427),
.B(n_356),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_390),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_396),
.B(n_377),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_392),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_407),
.B(n_378),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_427),
.B(n_382),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_430),
.B(n_384),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_407),
.B(n_385),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_430),
.B(n_445),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_417),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_390),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_407),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_417),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_445),
.B(n_365),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_408),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_416),
.B(n_380),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_417),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_390),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_440),
.B(n_373),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_405),
.B(n_387),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_390),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_SL g541 ( 
.A(n_450),
.B(n_342),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_456),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_456),
.B(n_343),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_405),
.B(n_178),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_440),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_417),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_417),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_417),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_440),
.B(n_214),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_434),
.A2(n_229),
.B1(n_263),
.B2(n_267),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_408),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_408),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_423),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_423),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_423),
.B(n_367),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_409),
.B(n_345),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_409),
.A2(n_286),
.B1(n_209),
.B2(n_213),
.Y(n_557)
);

INVx4_ASAP7_75t_SL g558 ( 
.A(n_453),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_423),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_409),
.B(n_159),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_423),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_423),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_409),
.B(n_252),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_408),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_409),
.B(n_159),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_409),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_410),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_451),
.B(n_159),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_451),
.B(n_373),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_399),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_424),
.B(n_322),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_399),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_425),
.B(n_159),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_410),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_451),
.B(n_222),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_424),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_410),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_424),
.B(n_289),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_399),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_399),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_424),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_410),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_451),
.A2(n_195),
.B1(n_246),
.B2(n_247),
.Y(n_583)
);

INVx5_ASAP7_75t_L g584 ( 
.A(n_453),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_451),
.B(n_225),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_424),
.B(n_304),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_424),
.B(n_200),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_399),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_438),
.B(n_205),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_451),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_438),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_425),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_438),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_438),
.Y(n_594)
);

BUFx4f_ASAP7_75t_L g595 ( 
.A(n_399),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_438),
.B(n_226),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_422),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_425),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_425),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_453),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_422),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_422),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_425),
.B(n_386),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_438),
.B(n_208),
.Y(n_604)
);

AND3x2_ASAP7_75t_L g605 ( 
.A(n_425),
.B(n_188),
.C(n_187),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_399),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_461),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_542),
.B(n_399),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_511),
.B(n_399),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_511),
.B(n_400),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_461),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_590),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_464),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_467),
.A2(n_429),
.B(n_422),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_528),
.B(n_400),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_499),
.B(n_400),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_519),
.B(n_400),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_496),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_469),
.B(n_400),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_485),
.A2(n_437),
.B1(n_453),
.B2(n_432),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_598),
.Y(n_621)
);

BUFx6f_ASAP7_75t_SL g622 ( 
.A(n_544),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_505),
.B(n_400),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_566),
.B(n_590),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_600),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_469),
.B(n_400),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_464),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_586),
.B(n_400),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_566),
.B(n_400),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_481),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_485),
.B(n_494),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_502),
.B(n_233),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_481),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_482),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_470),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_482),
.Y(n_636)
);

NOR3xp33_ASAP7_75t_L g637 ( 
.A(n_556),
.B(n_201),
.C(n_217),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_545),
.B(n_411),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_545),
.B(n_411),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_592),
.B(n_411),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_494),
.B(n_411),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_478),
.B(n_220),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_526),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_526),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_465),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_592),
.B(n_411),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_470),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_472),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_500),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_569),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_569),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_531),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_500),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_522),
.B(n_374),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_503),
.B(n_411),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_480),
.B(n_411),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_503),
.B(n_411),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_487),
.B(n_411),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_603),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_507),
.B(n_429),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_507),
.B(n_429),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_488),
.A2(n_437),
.B1(n_453),
.B2(n_432),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_603),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_501),
.B(n_515),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_587),
.B(n_429),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_589),
.B(n_432),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_472),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_604),
.B(n_432),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_599),
.B(n_453),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_501),
.B(n_437),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_522),
.B(n_374),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_490),
.A2(n_250),
.B1(n_244),
.B2(n_271),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_493),
.B(n_252),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_524),
.B(n_453),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_508),
.A2(n_273),
.B1(n_258),
.B2(n_257),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_525),
.B(n_453),
.Y(n_676)
);

BUFx6f_ASAP7_75t_SL g677 ( 
.A(n_544),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_473),
.Y(n_678)
);

NAND2xp33_ASAP7_75t_L g679 ( 
.A(n_473),
.B(n_453),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_533),
.B(n_453),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_457),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_L g682 ( 
.A(n_484),
.B(n_453),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_578),
.B(n_437),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_573),
.B(n_238),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_600),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_550),
.A2(n_278),
.B1(n_265),
.B2(n_261),
.C(n_253),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_501),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_549),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_484),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_543),
.B(n_241),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_486),
.B(n_394),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_571),
.B(n_243),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_486),
.B(n_491),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_549),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_530),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_491),
.B(n_394),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_497),
.B(n_394),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_501),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_497),
.B(n_395),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_538),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_512),
.B(n_395),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_474),
.B(n_224),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_501),
.A2(n_258),
.B1(n_257),
.B2(n_237),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_544),
.A2(n_187),
.B1(n_188),
.B2(n_273),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_515),
.A2(n_256),
.B1(n_259),
.B2(n_260),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_512),
.B(n_395),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_463),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_539),
.B(n_235),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_468),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_515),
.A2(n_237),
.B1(n_190),
.B2(n_305),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_509),
.B(n_239),
.Y(n_711)
);

OR2x4_ASAP7_75t_L g712 ( 
.A(n_563),
.B(n_173),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_538),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_513),
.B(n_397),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_513),
.B(n_517),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_468),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_535),
.B(n_515),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_530),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_596),
.A2(n_398),
.B(n_397),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_517),
.B(n_397),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_544),
.A2(n_305),
.B1(n_190),
.B2(n_291),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_471),
.Y(n_722)
);

NOR3xp33_ASAP7_75t_L g723 ( 
.A(n_466),
.B(n_240),
.C(n_254),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_521),
.B(n_523),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_529),
.B(n_398),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_595),
.A2(n_406),
.B(n_398),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_529),
.B(n_403),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_504),
.B(n_506),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_515),
.B(n_204),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_471),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_532),
.B(n_262),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_475),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_475),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_544),
.A2(n_204),
.B1(n_308),
.B2(n_223),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_532),
.B(n_264),
.Y(n_735)
);

INVx8_ASAP7_75t_L g736 ( 
.A(n_465),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_476),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_557),
.B(n_376),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_536),
.B(n_403),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_563),
.A2(n_232),
.B(n_176),
.C(n_181),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_536),
.B(n_275),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_527),
.B(n_242),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_510),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_530),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_546),
.B(n_403),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_476),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_546),
.B(n_287),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_547),
.B(n_206),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_465),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_547),
.B(n_406),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_548),
.B(n_301),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_595),
.A2(n_421),
.B(n_406),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_548),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_L g754 ( 
.A(n_553),
.B(n_206),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_553),
.B(n_412),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_479),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_516),
.B(n_292),
.C(n_249),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_479),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_492),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_483),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_557),
.B(n_251),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_554),
.B(n_412),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_559),
.B(n_412),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_559),
.B(n_413),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_561),
.B(n_223),
.Y(n_765)
);

OR2x6_ASAP7_75t_L g766 ( 
.A(n_465),
.B(n_291),
.Y(n_766)
);

BUFx8_ASAP7_75t_L g767 ( 
.A(n_541),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_516),
.A2(n_308),
.B1(n_421),
.B2(n_449),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_465),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_561),
.B(n_442),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_568),
.A2(n_428),
.B1(n_413),
.B2(n_449),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_562),
.B(n_442),
.Y(n_772)
);

INVx8_ASAP7_75t_L g773 ( 
.A(n_530),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_562),
.B(n_413),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_483),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_576),
.B(n_419),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_576),
.B(n_419),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_631),
.B(n_581),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_625),
.B(n_581),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_753),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_645),
.A2(n_595),
.B(n_460),
.Y(n_781)
);

AOI21x1_ASAP7_75t_L g782 ( 
.A1(n_683),
.A2(n_593),
.B(n_591),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_642),
.B(n_550),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_759),
.B(n_583),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_615),
.B(n_591),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_625),
.B(n_593),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_645),
.A2(n_460),
.B(n_459),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_607),
.B(n_611),
.Y(n_788)
);

AOI21x1_ASAP7_75t_L g789 ( 
.A1(n_683),
.A2(n_594),
.B(n_585),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_645),
.A2(n_460),
.B(n_459),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_607),
.B(n_594),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_609),
.A2(n_495),
.B(n_489),
.Y(n_792)
);

CKINVDCx8_ASAP7_75t_R g793 ( 
.A(n_618),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_625),
.B(n_537),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_611),
.B(n_583),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_614),
.A2(n_462),
.B(n_458),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_649),
.B(n_560),
.Y(n_797)
);

INVx11_ASAP7_75t_L g798 ( 
.A(n_767),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_645),
.A2(n_477),
.B(n_459),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_761),
.B(n_688),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_645),
.A2(n_477),
.B(n_459),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_773),
.A2(n_608),
.B(n_610),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_613),
.B(n_565),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_619),
.A2(n_626),
.B(n_623),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_654),
.B(n_575),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_612),
.A2(n_555),
.B1(n_540),
.B2(n_458),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_773),
.A2(n_520),
.B(n_477),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_694),
.Y(n_808)
);

AOI21xp33_ASAP7_75t_L g809 ( 
.A1(n_702),
.A2(n_268),
.B(n_255),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_613),
.B(n_458),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_SL g811 ( 
.A(n_622),
.B(n_176),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_653),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_625),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_627),
.B(n_462),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_627),
.B(n_462),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_671),
.B(n_376),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_773),
.A2(n_736),
.B(n_617),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_635),
.B(n_540),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_612),
.A2(n_540),
.B1(n_579),
.B2(n_588),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_773),
.A2(n_520),
.B(n_477),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_685),
.B(n_537),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_686),
.A2(n_282),
.B(n_278),
.C(n_309),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_736),
.A2(n_606),
.B(n_520),
.Y(n_823)
);

OAI21xp33_ASAP7_75t_L g824 ( 
.A1(n_711),
.A2(n_270),
.B(n_284),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_685),
.B(n_537),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_717),
.A2(n_579),
.B1(n_588),
.B2(n_520),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_635),
.B(n_579),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_736),
.A2(n_606),
.B(n_570),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_628),
.A2(n_606),
.B(n_570),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_647),
.B(n_588),
.Y(n_830)
);

OAI21xp33_ASAP7_75t_L g831 ( 
.A1(n_742),
.A2(n_274),
.B(n_281),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_675),
.A2(n_514),
.B(n_602),
.C(n_601),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_650),
.A2(n_514),
.B(n_602),
.C(n_601),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_647),
.B(n_489),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_665),
.A2(n_570),
.B(n_572),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_648),
.B(n_495),
.Y(n_836)
);

OR2x6_ASAP7_75t_L g837 ( 
.A(n_664),
.B(n_181),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_648),
.B(n_498),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_667),
.B(n_498),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_666),
.A2(n_572),
.B(n_537),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_700),
.B(n_713),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_667),
.B(n_678),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_668),
.A2(n_572),
.B(n_537),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_678),
.B(n_518),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_689),
.B(n_518),
.Y(n_845)
);

AND2x4_ASAP7_75t_SL g846 ( 
.A(n_698),
.B(n_580),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_685),
.Y(n_847)
);

CKINVDCx8_ASAP7_75t_R g848 ( 
.A(n_681),
.Y(n_848)
);

INVx11_ASAP7_75t_L g849 ( 
.A(n_767),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_724),
.A2(n_572),
.B1(n_597),
.B2(n_551),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_689),
.B(n_534),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_707),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_651),
.B(n_534),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_659),
.B(n_663),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_630),
.B(n_633),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_634),
.B(n_551),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_SL g857 ( 
.A(n_728),
.B(n_283),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_636),
.B(n_552),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_749),
.B(n_584),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_749),
.A2(n_580),
.B(n_597),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_616),
.A2(n_552),
.B(n_564),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_612),
.B(n_643),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_644),
.B(n_564),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_685),
.B(n_580),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_660),
.B(n_567),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_616),
.A2(n_567),
.B(n_574),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_SL g867 ( 
.A1(n_623),
.A2(n_196),
.B(n_215),
.C(n_218),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_680),
.B(n_674),
.Y(n_868)
);

BUFx4f_ASAP7_75t_L g869 ( 
.A(n_664),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_769),
.A2(n_580),
.B(n_582),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_621),
.B(n_558),
.Y(n_871)
);

AND2x4_ASAP7_75t_SL g872 ( 
.A(n_698),
.B(n_580),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_712),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_769),
.A2(n_582),
.B(n_577),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_641),
.A2(n_657),
.B(n_655),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_712),
.Y(n_876)
);

BUFx12f_ASAP7_75t_L g877 ( 
.A(n_767),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_738),
.B(n_379),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_768),
.A2(n_310),
.B(n_197),
.C(n_215),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_664),
.A2(n_574),
.B1(n_577),
.B2(n_290),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_661),
.B(n_419),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_629),
.A2(n_584),
.B(n_448),
.Y(n_882)
);

NAND3xp33_ASAP7_75t_L g883 ( 
.A(n_757),
.B(n_285),
.C(n_293),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_693),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_676),
.B(n_558),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_715),
.Y(n_886)
);

NOR2xp67_ASAP7_75t_SL g887 ( 
.A(n_695),
.B(n_584),
.Y(n_887)
);

CKINVDCx8_ASAP7_75t_R g888 ( 
.A(n_652),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_679),
.A2(n_682),
.B(n_620),
.Y(n_889)
);

OAI21xp33_ASAP7_75t_L g890 ( 
.A1(n_673),
.A2(n_294),
.B(n_295),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_629),
.A2(n_584),
.B(n_448),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_624),
.A2(n_584),
.B(n_448),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_679),
.A2(n_428),
.B(n_436),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_632),
.B(n_421),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_664),
.A2(n_296),
.B1(n_307),
.B2(n_428),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_682),
.A2(n_765),
.B(n_740),
.C(n_703),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_624),
.A2(n_447),
.B1(n_433),
.B2(n_436),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_715),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_669),
.A2(n_584),
.B(n_448),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_690),
.B(n_431),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_690),
.B(n_431),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_638),
.A2(n_444),
.B(n_436),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_638),
.B(n_431),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_698),
.B(n_558),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_656),
.B(n_558),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_743),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_640),
.A2(n_455),
.B(n_447),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_640),
.A2(n_455),
.B(n_447),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_646),
.A2(n_455),
.B(n_444),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_656),
.B(n_442),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_646),
.A2(n_455),
.B(n_444),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_708),
.B(n_379),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_658),
.B(n_442),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_658),
.A2(n_639),
.B(n_662),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_639),
.A2(n_433),
.B(n_441),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_704),
.A2(n_734),
.B(n_721),
.C(n_687),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_695),
.A2(n_449),
.B(n_433),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_705),
.B(n_442),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_707),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_692),
.B(n_441),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_709),
.B(n_442),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_709),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_692),
.B(n_441),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_716),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_622),
.B(n_5),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_716),
.B(n_722),
.Y(n_926)
);

AND2x2_ASAP7_75t_SL g927 ( 
.A(n_637),
.B(n_748),
.Y(n_927)
);

AO22x1_ASAP7_75t_L g928 ( 
.A1(n_723),
.A2(n_265),
.B1(n_197),
.B2(n_218),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_722),
.B(n_605),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_672),
.A2(n_300),
.B(n_221),
.Y(n_930)
);

AO21x1_ASAP7_75t_L g931 ( 
.A1(n_710),
.A2(n_196),
.B(n_221),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_730),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_719),
.A2(n_303),
.B(n_234),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_730),
.B(n_442),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_729),
.B(n_684),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_732),
.B(n_442),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_729),
.B(n_232),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_684),
.A2(n_303),
.B(n_245),
.C(n_253),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_732),
.Y(n_939)
);

AO21x1_ASAP7_75t_L g940 ( 
.A1(n_731),
.A2(n_735),
.B(n_741),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_733),
.B(n_454),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_733),
.B(n_454),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_729),
.Y(n_943)
);

BUFx8_ASAP7_75t_SL g944 ( 
.A(n_677),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_737),
.B(n_454),
.Y(n_945)
);

BUFx12f_ASAP7_75t_L g946 ( 
.A(n_729),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_737),
.B(n_454),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_746),
.B(n_443),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_677),
.B(n_6),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_765),
.A2(n_300),
.B(n_245),
.C(n_261),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_748),
.A2(n_234),
.B(n_266),
.C(n_282),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_718),
.A2(n_744),
.B(n_731),
.Y(n_952)
);

BUFx12f_ASAP7_75t_L g953 ( 
.A(n_766),
.Y(n_953)
);

BUFx12f_ASAP7_75t_L g954 ( 
.A(n_766),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_735),
.B(n_741),
.Y(n_955)
);

BUFx4f_ASAP7_75t_L g956 ( 
.A(n_766),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_744),
.A2(n_443),
.B(n_386),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_746),
.B(n_443),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_783),
.A2(n_670),
.B1(n_744),
.B2(n_766),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_780),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_800),
.B(n_747),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_800),
.B(n_670),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_812),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_884),
.B(n_747),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_877),
.Y(n_965)
);

CKINVDCx8_ASAP7_75t_R g966 ( 
.A(n_906),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_783),
.B(n_751),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_857),
.B(n_784),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_R g969 ( 
.A(n_848),
.B(n_754),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_813),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_809),
.A2(n_751),
.B(n_754),
.C(n_691),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_852),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_807),
.A2(n_670),
.B(n_726),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_955),
.B(n_940),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_784),
.A2(n_670),
.B1(n_771),
.B2(n_770),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_SL g976 ( 
.A1(n_889),
.A2(n_752),
.B(n_756),
.C(n_775),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_812),
.B(n_696),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_820),
.A2(n_745),
.B(n_776),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_823),
.A2(n_739),
.B(n_697),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_873),
.Y(n_980)
);

OAI21xp33_ASAP7_75t_L g981 ( 
.A1(n_831),
.A2(n_266),
.B(n_309),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_795),
.A2(n_755),
.B1(n_699),
.B2(n_774),
.Y(n_982)
);

O2A1O1Ixp5_ASAP7_75t_L g983 ( 
.A1(n_918),
.A2(n_777),
.B(n_701),
.C(n_706),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_805),
.B(n_714),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_878),
.B(n_756),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_927),
.B(n_775),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_896),
.A2(n_750),
.B(n_720),
.C(n_764),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_856),
.Y(n_988)
);

O2A1O1Ixp5_ASAP7_75t_L g989 ( 
.A1(n_918),
.A2(n_725),
.B(n_763),
.C(n_762),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_858),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_813),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_828),
.A2(n_727),
.B(n_770),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_822),
.A2(n_310),
.B(n_772),
.C(n_758),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_802),
.A2(n_760),
.B(n_758),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_803),
.A2(n_383),
.B1(n_381),
.B2(n_156),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_808),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_SL g997 ( 
.A(n_793),
.B(n_383),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_816),
.B(n_381),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_912),
.B(n_841),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_935),
.A2(n_148),
.B1(n_146),
.B2(n_145),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_808),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_817),
.A2(n_144),
.B(n_143),
.Y(n_1002)
);

INVxp67_ASAP7_75t_SL g1003 ( 
.A(n_788),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_SL g1004 ( 
.A(n_888),
.B(n_136),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_R g1005 ( 
.A(n_811),
.B(n_847),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_914),
.A2(n_132),
.B(n_131),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_863),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_922),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_875),
.A2(n_119),
.B(n_117),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_781),
.A2(n_115),
.B(n_111),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_924),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_869),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_869),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_873),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_785),
.A2(n_109),
.B(n_104),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_939),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_927),
.B(n_92),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_804),
.A2(n_74),
.B(n_72),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_853),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_840),
.A2(n_64),
.B(n_63),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_SL g1021 ( 
.A(n_797),
.B(n_7),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_854),
.B(n_8),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_843),
.A2(n_62),
.B(n_61),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_868),
.A2(n_9),
.B(n_10),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_822),
.A2(n_10),
.B(n_11),
.C(n_14),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_938),
.A2(n_11),
.B(n_17),
.C(n_18),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_824),
.A2(n_898),
.B(n_886),
.C(n_916),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_868),
.A2(n_835),
.B(n_842),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_787),
.A2(n_790),
.B(n_829),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_946),
.B(n_17),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_799),
.A2(n_57),
.B(n_22),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_876),
.B(n_18),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_SL g1033 ( 
.A1(n_925),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_876),
.B(n_23),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_801),
.A2(n_57),
.B(n_31),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_847),
.B(n_27),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_794),
.A2(n_51),
.B(n_32),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_778),
.B(n_31),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_956),
.B(n_34),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_916),
.A2(n_36),
.B(n_37),
.C(n_39),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_956),
.B(n_41),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_855),
.B(n_43),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_794),
.A2(n_45),
.B(n_47),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_826),
.A2(n_49),
.B1(n_50),
.B2(n_862),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_821),
.A2(n_50),
.B(n_825),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_890),
.B(n_943),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_943),
.B(n_883),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_937),
.B(n_925),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_821),
.A2(n_825),
.B(n_864),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_944),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_837),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_864),
.A2(n_865),
.B(n_779),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_937),
.B(n_949),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_779),
.A2(n_786),
.B(n_814),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_938),
.A2(n_879),
.B(n_930),
.C(n_950),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_871),
.Y(n_1056)
);

O2A1O1Ixp5_ASAP7_75t_L g1057 ( 
.A1(n_894),
.A2(n_880),
.B(n_933),
.C(n_905),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_900),
.A2(n_901),
.B(n_920),
.C(n_923),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_837),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_885),
.B(n_952),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_895),
.B(n_837),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_885),
.B(n_953),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_871),
.B(n_846),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_879),
.A2(n_950),
.B(n_867),
.C(n_951),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_867),
.A2(n_929),
.B(n_949),
.C(n_905),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_881),
.B(n_919),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_932),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_954),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_791),
.B(n_903),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_782),
.A2(n_796),
.B(n_902),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_850),
.A2(n_786),
.B1(n_904),
.B2(n_830),
.Y(n_1071)
);

INVxp33_ASAP7_75t_SL g1072 ( 
.A(n_798),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_926),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_810),
.B(n_827),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_931),
.A2(n_893),
.B(n_833),
.C(n_910),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_904),
.A2(n_818),
.B1(n_815),
.B2(n_872),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_846),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_928),
.B(n_836),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_849),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_872),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_859),
.Y(n_1081)
);

OAI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_897),
.A2(n_839),
.B(n_845),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_834),
.A2(n_851),
.B1(n_844),
.B2(n_838),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_789),
.B(n_892),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_859),
.A2(n_819),
.B1(n_910),
.B2(n_913),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_SL g1086 ( 
.A1(n_913),
.A2(n_921),
.B(n_941),
.C(n_948),
.Y(n_1086)
);

AOI21x1_ASAP7_75t_L g1087 ( 
.A1(n_921),
.A2(n_941),
.B(n_870),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_SL g1088 ( 
.A(n_957),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_915),
.A2(n_832),
.B(n_806),
.C(n_917),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_934),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_936),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_792),
.A2(n_861),
.B1(n_866),
.B2(n_911),
.Y(n_1092)
);

NOR2xp67_ASAP7_75t_L g1093 ( 
.A(n_899),
.B(n_882),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_942),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_907),
.A2(n_908),
.B1(n_909),
.B2(n_958),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_874),
.B(n_860),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_945),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_947),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_891),
.B(n_887),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_914),
.A2(n_889),
.B(n_505),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_807),
.A2(n_645),
.B(n_773),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_808),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_966),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_SL g1104 ( 
.A1(n_1027),
.A2(n_1017),
.B(n_1040),
.C(n_974),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_999),
.B(n_1048),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_1071),
.A2(n_1085),
.A3(n_987),
.B(n_1028),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1070),
.A2(n_1029),
.B(n_994),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_968),
.B(n_967),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_979),
.A2(n_978),
.B(n_1100),
.Y(n_1109)
);

AO22x1_ASAP7_75t_L g1110 ( 
.A1(n_1061),
.A2(n_1034),
.B1(n_1032),
.B2(n_1046),
.Y(n_1110)
);

CKINVDCx6p67_ASAP7_75t_R g1111 ( 
.A(n_965),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1057),
.A2(n_989),
.B(n_983),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_973),
.A2(n_1058),
.B(n_992),
.Y(n_1113)
);

BUFx8_ASAP7_75t_L g1114 ( 
.A(n_980),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1021),
.A2(n_984),
.B1(n_1053),
.B2(n_1041),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_977),
.B(n_963),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_974),
.A2(n_1092),
.B(n_1084),
.Y(n_1117)
);

BUFx8_ASAP7_75t_L g1118 ( 
.A(n_1079),
.Y(n_1118)
);

AOI221xp5_ASAP7_75t_SL g1119 ( 
.A1(n_1025),
.A2(n_1026),
.B1(n_981),
.B2(n_1055),
.C(n_1044),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1012),
.Y(n_1120)
);

OAI21xp33_ASAP7_75t_L g1121 ( 
.A1(n_997),
.A2(n_984),
.B(n_977),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_971),
.A2(n_1046),
.B(n_1065),
.C(n_1061),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_996),
.Y(n_1123)
);

OAI22x1_ASAP7_75t_L g1124 ( 
.A1(n_1039),
.A2(n_1041),
.B1(n_1047),
.B2(n_1062),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1096),
.A2(n_1069),
.B(n_1003),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1039),
.A2(n_962),
.B1(n_1047),
.B2(n_961),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1011),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1101),
.A2(n_1003),
.B(n_1096),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1087),
.A2(n_1054),
.B(n_1049),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_982),
.A2(n_1060),
.B(n_1089),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1060),
.A2(n_1083),
.B(n_1092),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_959),
.A2(n_1076),
.A3(n_1052),
.B(n_1074),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_960),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1014),
.B(n_1032),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_SL g1135 ( 
.A1(n_986),
.A2(n_1036),
.B(n_964),
.C(n_976),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1012),
.B(n_1013),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1075),
.A2(n_975),
.B(n_1088),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_1074),
.A2(n_1018),
.A3(n_995),
.B(n_1045),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_976),
.A2(n_1082),
.B(n_1099),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1084),
.A2(n_1095),
.B(n_1006),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1024),
.B(n_1022),
.C(n_1042),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1019),
.B(n_988),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_SL g1143 ( 
.A1(n_1036),
.A2(n_1038),
.B(n_1078),
.C(n_1073),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1086),
.A2(n_985),
.B(n_1066),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1095),
.A2(n_1020),
.B(n_1023),
.Y(n_1145)
);

NOR2xp67_ASAP7_75t_L g1146 ( 
.A(n_996),
.B(n_1102),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1012),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1093),
.A2(n_1009),
.B(n_1007),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1001),
.Y(n_1149)
);

OA21x2_ASAP7_75t_L g1150 ( 
.A1(n_1031),
.A2(n_1035),
.B(n_1002),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1014),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_969),
.B(n_1102),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_990),
.A2(n_998),
.B(n_1010),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1090),
.A2(n_1015),
.B(n_1097),
.Y(n_1154)
);

AO22x1_ASAP7_75t_L g1155 ( 
.A1(n_1034),
.A2(n_1062),
.B1(n_1013),
.B2(n_1012),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1008),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_1001),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1072),
.Y(n_1158)
);

AO32x2_ASAP7_75t_L g1159 ( 
.A1(n_970),
.A2(n_1064),
.A3(n_993),
.B1(n_1033),
.B2(n_1088),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1016),
.A2(n_1013),
.B1(n_1000),
.B2(n_1063),
.Y(n_1160)
);

O2A1O1Ixp5_ASAP7_75t_L g1161 ( 
.A1(n_1037),
.A2(n_1043),
.B(n_970),
.C(n_991),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1004),
.A2(n_1013),
.B1(n_1059),
.B2(n_1051),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1091),
.A2(n_1094),
.B(n_1098),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1056),
.B(n_1063),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1094),
.A2(n_1080),
.B(n_1081),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1067),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1077),
.A2(n_1081),
.B1(n_1094),
.B2(n_1030),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_969),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1081),
.B(n_1005),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1081),
.A2(n_1030),
.B(n_1005),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1030),
.B(n_1050),
.Y(n_1171)
);

OA21x2_ASAP7_75t_L g1172 ( 
.A1(n_1068),
.A2(n_1100),
.B(n_1070),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1071),
.A2(n_940),
.A3(n_1085),
.B(n_987),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_973),
.A2(n_645),
.B(n_979),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1071),
.A2(n_940),
.A3(n_1085),
.B(n_987),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1100),
.A2(n_1070),
.B(n_1057),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_973),
.A2(n_645),
.B(n_979),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_974),
.A2(n_1100),
.B(n_1029),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_984),
.B(n_1019),
.Y(n_1179)
);

BUFx10_ASAP7_75t_L g1180 ( 
.A(n_1062),
.Y(n_1180)
);

O2A1O1Ixp5_ASAP7_75t_SL g1181 ( 
.A1(n_974),
.A2(n_1084),
.B(n_692),
.C(n_961),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1070),
.A2(n_1029),
.B(n_994),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1070),
.A2(n_1029),
.B(n_994),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_974),
.A2(n_783),
.B(n_967),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_975),
.A2(n_783),
.B1(n_516),
.B2(n_800),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1070),
.A2(n_1029),
.B(n_994),
.Y(n_1186)
);

CKINVDCx11_ASAP7_75t_R g1187 ( 
.A(n_965),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_968),
.A2(n_783),
.B1(n_784),
.B2(n_800),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1071),
.A2(n_940),
.A3(n_1085),
.B(n_987),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_968),
.A2(n_783),
.B1(n_784),
.B2(n_761),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_975),
.A2(n_783),
.B1(n_516),
.B2(n_800),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_968),
.B(n_783),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_984),
.B(n_1019),
.Y(n_1193)
);

AO21x1_ASAP7_75t_L g1194 ( 
.A1(n_974),
.A2(n_783),
.B(n_967),
.Y(n_1194)
);

CKINVDCx11_ASAP7_75t_R g1195 ( 
.A(n_965),
.Y(n_1195)
);

NOR2xp67_ASAP7_75t_L g1196 ( 
.A(n_1079),
.B(n_728),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1012),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_963),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_972),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1012),
.B(n_1013),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_996),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1100),
.A2(n_783),
.B(n_1057),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1070),
.A2(n_1029),
.B(n_994),
.Y(n_1203)
);

AO21x1_ASAP7_75t_L g1204 ( 
.A1(n_974),
.A2(n_783),
.B(n_967),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1100),
.A2(n_783),
.B(n_1057),
.Y(n_1205)
);

NOR2x1_ASAP7_75t_L g1206 ( 
.A(n_970),
.B(n_728),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_R g1207 ( 
.A(n_966),
.B(n_618),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_1012),
.B(n_1013),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_960),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_999),
.B(n_1048),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1070),
.A2(n_1029),
.B(n_994),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_960),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_999),
.B(n_728),
.Y(n_1213)
);

AO22x2_ASAP7_75t_L g1214 ( 
.A1(n_968),
.A2(n_1044),
.B1(n_1041),
.B2(n_1039),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_973),
.A2(n_645),
.B(n_979),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1071),
.A2(n_940),
.A3(n_1085),
.B(n_987),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1070),
.A2(n_1029),
.B(n_994),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_973),
.A2(n_645),
.B(n_979),
.Y(n_1218)
);

OAI22x1_ASAP7_75t_L g1219 ( 
.A1(n_968),
.A2(n_783),
.B1(n_516),
.B2(n_550),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_968),
.B(n_783),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1012),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_984),
.B(n_1019),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_984),
.B(n_1019),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_973),
.A2(n_645),
.B(n_979),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_973),
.A2(n_645),
.B(n_979),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_973),
.A2(n_645),
.B(n_979),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1070),
.A2(n_1029),
.B(n_994),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_960),
.Y(n_1228)
);

AO21x1_ASAP7_75t_L g1229 ( 
.A1(n_974),
.A2(n_783),
.B(n_967),
.Y(n_1229)
);

BUFx12f_ASAP7_75t_L g1230 ( 
.A(n_965),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_979),
.A2(n_978),
.B(n_1100),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_968),
.A2(n_783),
.B(n_800),
.C(n_642),
.Y(n_1232)
);

NOR2x1_ASAP7_75t_SL g1233 ( 
.A(n_1012),
.B(n_1013),
.Y(n_1233)
);

OAI22x1_ASAP7_75t_L g1234 ( 
.A1(n_968),
.A2(n_783),
.B1(n_516),
.B2(n_550),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_975),
.A2(n_783),
.B1(n_516),
.B2(n_800),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_960),
.Y(n_1236)
);

AO22x2_ASAP7_75t_L g1237 ( 
.A1(n_968),
.A2(n_1044),
.B1(n_1041),
.B2(n_1039),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_984),
.B(n_1019),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_999),
.B(n_728),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_968),
.A2(n_783),
.B(n_800),
.C(n_642),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_996),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_980),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1207),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1187),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1185),
.A2(n_1191),
.B1(n_1235),
.B2(n_1192),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1185),
.A2(n_1235),
.B1(n_1191),
.B2(n_1220),
.Y(n_1246)
);

BUFx10_ASAP7_75t_L g1247 ( 
.A(n_1116),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1190),
.A2(n_1234),
.B1(n_1219),
.B2(n_1188),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1188),
.A2(n_1108),
.B1(n_1214),
.B2(n_1237),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1232),
.A2(n_1240),
.B1(n_1115),
.B2(n_1126),
.Y(n_1250)
);

INVx6_ASAP7_75t_L g1251 ( 
.A(n_1118),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1121),
.A2(n_1115),
.B1(n_1126),
.B2(n_1162),
.Y(n_1252)
);

AOI22x1_ASAP7_75t_L g1253 ( 
.A1(n_1124),
.A2(n_1214),
.B1(n_1237),
.B2(n_1202),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1195),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1114),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1118),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1121),
.A2(n_1205),
.B1(n_1202),
.B2(n_1204),
.Y(n_1257)
);

OAI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1179),
.A2(n_1193),
.B1(n_1223),
.B2(n_1222),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1205),
.A2(n_1184),
.B1(n_1229),
.B2(n_1194),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1179),
.A2(n_1222),
.B1(n_1223),
.B2(n_1193),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1209),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1238),
.A2(n_1141),
.B1(n_1130),
.B2(n_1142),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1230),
.Y(n_1263)
);

OAI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1238),
.A2(n_1162),
.B1(n_1142),
.B2(n_1239),
.Y(n_1264)
);

BUFx8_ASAP7_75t_L g1265 ( 
.A(n_1242),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1167),
.A2(n_1110),
.B1(n_1105),
.B2(n_1210),
.Y(n_1266)
);

INVx6_ASAP7_75t_L g1267 ( 
.A(n_1114),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1167),
.A2(n_1152),
.B1(n_1196),
.B2(n_1160),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1201),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1160),
.A2(n_1168),
.B1(n_1206),
.B2(n_1213),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1158),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1141),
.A2(n_1131),
.B1(n_1180),
.B2(n_1137),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1122),
.A2(n_1146),
.B1(n_1169),
.B2(n_1170),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1212),
.A2(n_1236),
.B1(n_1228),
.B2(n_1156),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1111),
.Y(n_1275)
);

CKINVDCx6p67_ASAP7_75t_R g1276 ( 
.A(n_1103),
.Y(n_1276)
);

INVx4_ASAP7_75t_L g1277 ( 
.A(n_1120),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1134),
.B(n_1241),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1123),
.Y(n_1279)
);

BUFx8_ASAP7_75t_L g1280 ( 
.A(n_1171),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1166),
.A2(n_1149),
.B1(n_1178),
.B2(n_1125),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1180),
.A2(n_1170),
.B1(n_1159),
.B2(n_1112),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1157),
.B(n_1155),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1178),
.A2(n_1125),
.B1(n_1112),
.B2(n_1199),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1127),
.A2(n_1113),
.B1(n_1151),
.B2(n_1153),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1169),
.A2(n_1198),
.B1(n_1163),
.B2(n_1208),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1159),
.A2(n_1233),
.B1(n_1119),
.B2(n_1117),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1144),
.A2(n_1150),
.B1(n_1139),
.B2(n_1231),
.Y(n_1288)
);

BUFx10_ASAP7_75t_L g1289 ( 
.A(n_1136),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1164),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1119),
.A2(n_1136),
.B1(n_1200),
.B2(n_1164),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1120),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1120),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1208),
.A2(n_1200),
.B1(n_1154),
.B2(n_1165),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1143),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1147),
.Y(n_1296)
);

CKINVDCx6p67_ASAP7_75t_R g1297 ( 
.A(n_1208),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1147),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1159),
.A2(n_1117),
.B1(n_1231),
.B2(n_1109),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1109),
.A2(n_1150),
.B1(n_1104),
.B2(n_1172),
.Y(n_1300)
);

CKINVDCx6p67_ASAP7_75t_R g1301 ( 
.A(n_1197),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1172),
.A2(n_1145),
.B1(n_1197),
.B2(n_1221),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1221),
.B(n_1132),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1221),
.A2(n_1148),
.B1(n_1176),
.B2(n_1128),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1176),
.Y(n_1305)
);

OAI21xp33_ASAP7_75t_L g1306 ( 
.A1(n_1181),
.A2(n_1129),
.B(n_1140),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1135),
.A2(n_1218),
.B1(n_1215),
.B2(n_1174),
.Y(n_1307)
);

CKINVDCx11_ASAP7_75t_R g1308 ( 
.A(n_1161),
.Y(n_1308)
);

INVx5_ASAP7_75t_L g1309 ( 
.A(n_1138),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1173),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1177),
.A2(n_1226),
.B1(n_1225),
.B2(n_1224),
.Y(n_1311)
);

BUFx4_ASAP7_75t_R g1312 ( 
.A(n_1173),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1175),
.A2(n_1216),
.B1(n_1189),
.B2(n_1106),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1138),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1175),
.A2(n_1189),
.B1(n_1216),
.B2(n_1106),
.Y(n_1315)
);

INVx8_ASAP7_75t_L g1316 ( 
.A(n_1175),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1216),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1107),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1182),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1183),
.A2(n_1186),
.B1(n_1203),
.B2(n_1211),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1217),
.A2(n_783),
.B1(n_1190),
.B2(n_1185),
.Y(n_1321)
);

BUFx8_ASAP7_75t_SL g1322 ( 
.A(n_1227),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1118),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1185),
.A2(n_1191),
.B1(n_1235),
.B2(n_783),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1185),
.A2(n_1191),
.B1(n_1235),
.B2(n_783),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1118),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1190),
.A2(n_1188),
.B1(n_783),
.B2(n_1232),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1133),
.Y(n_1328)
);

CKINVDCx11_ASAP7_75t_R g1329 ( 
.A(n_1187),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1187),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1114),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1190),
.A2(n_783),
.B1(n_1188),
.B2(n_450),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1118),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1185),
.A2(n_1191),
.B1(n_1235),
.B2(n_783),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1190),
.A2(n_1188),
.B1(n_783),
.B2(n_1232),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1188),
.A2(n_1235),
.B1(n_1185),
.B2(n_1191),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1185),
.A2(n_1191),
.B1(n_1235),
.B2(n_783),
.Y(n_1337)
);

OAI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1188),
.A2(n_1235),
.B1(n_1185),
.B2(n_1191),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1185),
.A2(n_1191),
.B1(n_1235),
.B2(n_783),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1207),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1190),
.A2(n_1188),
.B1(n_783),
.B2(n_1232),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1120),
.Y(n_1342)
);

OAI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1190),
.A2(n_783),
.B(n_1188),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1187),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1219),
.A2(n_783),
.B1(n_1234),
.B2(n_1220),
.Y(n_1345)
);

OAI21xp33_ASAP7_75t_L g1346 ( 
.A1(n_1190),
.A2(n_783),
.B(n_1188),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1190),
.A2(n_1188),
.B1(n_783),
.B2(n_1232),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1190),
.A2(n_783),
.B1(n_1191),
.B2(n_1185),
.Y(n_1348)
);

CKINVDCx6p67_ASAP7_75t_R g1349 ( 
.A(n_1187),
.Y(n_1349)
);

INVx6_ASAP7_75t_L g1350 ( 
.A(n_1118),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1185),
.A2(n_1191),
.B1(n_1235),
.B2(n_783),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1120),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1213),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1185),
.A2(n_1191),
.B1(n_1235),
.B2(n_783),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1324),
.B(n_1337),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1310),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1329),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1269),
.Y(n_1358)
);

NAND2x1p5_ASAP7_75t_L g1359 ( 
.A(n_1295),
.B(n_1309),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1324),
.B(n_1337),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1353),
.B(n_1290),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1260),
.B(n_1343),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1320),
.A2(n_1311),
.B(n_1288),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1317),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1312),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_SL g1366 ( 
.A(n_1248),
.B(n_1348),
.C(n_1351),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1307),
.A2(n_1306),
.B(n_1319),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1316),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1318),
.A2(n_1336),
.B(n_1338),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1316),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1316),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1320),
.A2(n_1288),
.B(n_1304),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1303),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1261),
.Y(n_1375)
);

OAI211xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1248),
.A2(n_1354),
.B(n_1325),
.C(n_1334),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1328),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1322),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1313),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1283),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1304),
.A2(n_1284),
.B(n_1285),
.Y(n_1382)
);

OAI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1327),
.A2(n_1335),
.B(n_1341),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1313),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1305),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1259),
.A2(n_1253),
.B(n_1284),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1347),
.A2(n_1354),
.B(n_1351),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1315),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1315),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1309),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1325),
.B(n_1334),
.Y(n_1391)
);

BUFx10_ASAP7_75t_L g1392 ( 
.A(n_1251),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1309),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1346),
.A2(n_1332),
.B1(n_1339),
.B2(n_1338),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1278),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1285),
.A2(n_1294),
.B(n_1259),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1286),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1314),
.Y(n_1398)
);

INVx4_ASAP7_75t_SL g1399 ( 
.A(n_1267),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1336),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1299),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1265),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1262),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1268),
.Y(n_1404)
);

INVx4_ASAP7_75t_SL g1405 ( 
.A(n_1267),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1339),
.A2(n_1250),
.B1(n_1321),
.B2(n_1249),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1257),
.B(n_1252),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1281),
.A2(n_1262),
.B(n_1273),
.Y(n_1408)
);

INVxp67_ASAP7_75t_SL g1409 ( 
.A(n_1281),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1308),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1258),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1258),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1300),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1264),
.A2(n_1270),
.B1(n_1266),
.B2(n_1260),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1300),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1247),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1257),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1302),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1264),
.B(n_1345),
.Y(n_1419)
);

OAI21xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1291),
.A2(n_1274),
.B(n_1287),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1302),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1267),
.B(n_1350),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1287),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1265),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1282),
.B(n_1272),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1274),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1282),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1279),
.A2(n_1331),
.B(n_1255),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1330),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1297),
.Y(n_1430)
);

OAI211xp5_ASAP7_75t_L g1431 ( 
.A1(n_1394),
.A2(n_1383),
.B(n_1420),
.C(n_1414),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1375),
.Y(n_1432)
);

NAND4xp25_ASAP7_75t_L g1433 ( 
.A(n_1406),
.B(n_1326),
.C(n_1323),
.D(n_1256),
.Y(n_1433)
);

AND2x2_ASAP7_75t_SL g1434 ( 
.A(n_1425),
.B(n_1298),
.Y(n_1434)
);

AND2x2_ASAP7_75t_SL g1435 ( 
.A(n_1425),
.B(n_1298),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1416),
.B(n_1361),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1420),
.A2(n_1352),
.B(n_1296),
.C(n_1292),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1392),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1375),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1401),
.B(n_1333),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1387),
.A2(n_1342),
.B(n_1277),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1395),
.B(n_1247),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1374),
.B(n_1352),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1381),
.B(n_1280),
.Y(n_1444)
);

NOR2x1_ASAP7_75t_SL g1445 ( 
.A(n_1422),
.B(n_1344),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1418),
.B(n_1276),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1377),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1368),
.B(n_1271),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1428),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1366),
.A2(n_1275),
.B1(n_1340),
.B2(n_1243),
.C(n_1244),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1418),
.B(n_1301),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1376),
.A2(n_1280),
.B1(n_1350),
.B2(n_1251),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1370),
.B(n_1293),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1414),
.A2(n_1289),
.B(n_1251),
.Y(n_1454)
);

AO21x1_ASAP7_75t_L g1455 ( 
.A1(n_1419),
.A2(n_1350),
.B(n_1349),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1358),
.B(n_1355),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1363),
.A2(n_1263),
.B(n_1254),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1355),
.A2(n_1360),
.B(n_1419),
.C(n_1408),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1379),
.B(n_1384),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1360),
.B(n_1362),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1404),
.B(n_1380),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1462)
);

NAND4xp25_ASAP7_75t_L g1463 ( 
.A(n_1404),
.B(n_1398),
.C(n_1417),
.D(n_1412),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1388),
.B(n_1389),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1410),
.A2(n_1373),
.B1(n_1378),
.B2(n_1398),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1422),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1428),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1363),
.A2(n_1382),
.B(n_1372),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1380),
.B(n_1400),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1389),
.B(n_1365),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1408),
.A2(n_1396),
.B(n_1382),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1407),
.A2(n_1396),
.B(n_1373),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1421),
.B(n_1413),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1372),
.A2(n_1359),
.B(n_1390),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1385),
.B(n_1369),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1410),
.A2(n_1391),
.B1(n_1397),
.B2(n_1400),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1357),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1427),
.A2(n_1403),
.B1(n_1417),
.B2(n_1409),
.C(n_1412),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1415),
.B(n_1427),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1391),
.A2(n_1407),
.B1(n_1410),
.B2(n_1403),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1392),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1468),
.B(n_1367),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1467),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1468),
.B(n_1367),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1475),
.B(n_1385),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1449),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1468),
.B(n_1367),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1471),
.B(n_1369),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1474),
.B(n_1371),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1474),
.B(n_1364),
.Y(n_1490)
);

NAND2x1_ASAP7_75t_L g1491 ( 
.A(n_1466),
.B(n_1393),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1431),
.A2(n_1410),
.B1(n_1423),
.B2(n_1378),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1432),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1472),
.A2(n_1433),
.B1(n_1480),
.B2(n_1460),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1442),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1478),
.A2(n_1411),
.B1(n_1423),
.B2(n_1463),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1473),
.B(n_1439),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1447),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1450),
.A2(n_1386),
.B1(n_1426),
.B2(n_1378),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1473),
.B(n_1356),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1443),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1434),
.A2(n_1435),
.B1(n_1461),
.B2(n_1386),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1470),
.B(n_1428),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1483),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1482),
.B(n_1484),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1482),
.B(n_1459),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1482),
.B(n_1462),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1503),
.B(n_1456),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1482),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1490),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1484),
.B(n_1487),
.Y(n_1511)
);

OAI221xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1496),
.A2(n_1458),
.B1(n_1437),
.B2(n_1476),
.C(n_1452),
.Y(n_1512)
);

INVx3_ASAP7_75t_SL g1513 ( 
.A(n_1486),
.Y(n_1513)
);

NOR2x1_ASAP7_75t_L g1514 ( 
.A(n_1491),
.B(n_1483),
.Y(n_1514)
);

AOI21xp33_ASAP7_75t_L g1515 ( 
.A1(n_1492),
.A2(n_1458),
.B(n_1437),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1494),
.A2(n_1386),
.B1(n_1455),
.B2(n_1435),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1489),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1498),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1484),
.B(n_1462),
.Y(n_1519)
);

INVxp67_ASAP7_75t_L g1520 ( 
.A(n_1498),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1503),
.B(n_1464),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1501),
.B(n_1464),
.Y(n_1522)
);

BUFx2_ASAP7_75t_SL g1523 ( 
.A(n_1490),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1484),
.B(n_1470),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1487),
.B(n_1479),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1489),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1493),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1494),
.B(n_1440),
.C(n_1446),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1503),
.B(n_1479),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1493),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1491),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1493),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1491),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1487),
.B(n_1457),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1492),
.A2(n_1386),
.B1(n_1455),
.B2(n_1434),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1487),
.B(n_1457),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1493),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1501),
.B(n_1457),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1496),
.A2(n_1469),
.B1(n_1465),
.B2(n_1426),
.C(n_1436),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1486),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1528),
.B(n_1502),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1510),
.Y(n_1542)
);

AND2x2_ASAP7_75t_SL g1543 ( 
.A(n_1516),
.B(n_1488),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1506),
.B(n_1507),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1527),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1527),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1518),
.B(n_1500),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1527),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1521),
.B(n_1497),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1531),
.B(n_1489),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1531),
.B(n_1489),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1530),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1512),
.A2(n_1499),
.B1(n_1502),
.B2(n_1440),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1521),
.B(n_1497),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1519),
.B(n_1495),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1530),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1521),
.B(n_1497),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1529),
.B(n_1497),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1532),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1540),
.B(n_1495),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1528),
.A2(n_1499),
.B1(n_1454),
.B2(n_1422),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1540),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1519),
.B(n_1489),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1532),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1514),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1529),
.B(n_1485),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1519),
.B(n_1489),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1537),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1513),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1562),
.B(n_1539),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1549),
.B(n_1529),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1544),
.B(n_1555),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1542),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1545),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1542),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1544),
.B(n_1517),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1549),
.B(n_1508),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1555),
.B(n_1517),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1550),
.B(n_1514),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1553),
.B(n_1515),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1554),
.B(n_1508),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1560),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1541),
.B(n_1539),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1545),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1546),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1546),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1550),
.B(n_1517),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1550),
.B(n_1526),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1554),
.B(n_1508),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1543),
.B(n_1553),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1557),
.B(n_1510),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1543),
.B(n_1519),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1550),
.B(n_1526),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1543),
.B(n_1525),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1548),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1569),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1548),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1561),
.A2(n_1512),
.B1(n_1516),
.B2(n_1535),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1569),
.B(n_1525),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1542),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1551),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1547),
.B(n_1525),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1552),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1547),
.B(n_1525),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1561),
.B(n_1522),
.Y(n_1605)
);

NAND3xp33_ASAP7_75t_L g1606 ( 
.A(n_1565),
.B(n_1515),
.C(n_1535),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1551),
.B(n_1526),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1552),
.Y(n_1608)
);

NOR3x1_ASAP7_75t_L g1609 ( 
.A(n_1565),
.B(n_1444),
.C(n_1430),
.Y(n_1609)
);

NAND2x1p5_ASAP7_75t_L g1610 ( 
.A(n_1551),
.B(n_1514),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1551),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1611),
.B(n_1563),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1572),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1611),
.B(n_1563),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1601),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1574),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1572),
.Y(n_1617)
);

AOI32xp33_ASAP7_75t_L g1618 ( 
.A1(n_1590),
.A2(n_1536),
.A3(n_1534),
.B1(n_1511),
.B2(n_1505),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1583),
.B(n_1524),
.Y(n_1619)
);

NAND4xp25_ASAP7_75t_L g1620 ( 
.A(n_1580),
.B(n_1446),
.C(n_1441),
.D(n_1451),
.Y(n_1620)
);

AOI22x1_ASAP7_75t_L g1621 ( 
.A1(n_1596),
.A2(n_1357),
.B1(n_1477),
.B2(n_1610),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1574),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1570),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1601),
.B(n_1567),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1601),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1605),
.B(n_1592),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1594),
.B(n_1557),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1610),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1584),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1599),
.B(n_1558),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1601),
.B(n_1567),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1582),
.B(n_1524),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1584),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1585),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1598),
.A2(n_1606),
.B(n_1610),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1577),
.B(n_1558),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1606),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1577),
.B(n_1581),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1585),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1573),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1581),
.B(n_1566),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1573),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1586),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1589),
.B(n_1477),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1609),
.B(n_1524),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1579),
.A2(n_1488),
.B1(n_1466),
.B2(n_1534),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1616),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1616),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1615),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1637),
.A2(n_1509),
.B1(n_1513),
.B2(n_1571),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1613),
.B(n_1617),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1623),
.B(n_1609),
.Y(n_1652)
);

OAI211xp5_ASAP7_75t_L g1653 ( 
.A1(n_1635),
.A2(n_1536),
.B(n_1534),
.C(n_1488),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1615),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_SL g1655 ( 
.A(n_1621),
.B(n_1429),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1621),
.A2(n_1402),
.B1(n_1424),
.B2(n_1513),
.C(n_1523),
.Y(n_1656)
);

AOI21xp33_ASAP7_75t_SL g1657 ( 
.A1(n_1644),
.A2(n_1513),
.B(n_1428),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1620),
.A2(n_1488),
.B1(n_1536),
.B2(n_1534),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1622),
.Y(n_1659)
);

OAI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1618),
.A2(n_1402),
.B1(n_1424),
.B2(n_1513),
.C(n_1523),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1619),
.B(n_1578),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1613),
.B(n_1579),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1626),
.A2(n_1617),
.B1(n_1645),
.B2(n_1643),
.C(n_1634),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1626),
.B(n_1578),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1627),
.A2(n_1579),
.B1(n_1536),
.B2(n_1466),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_L g1666 ( 
.A(n_1646),
.B(n_1402),
.C(n_1424),
.D(n_1607),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1633),
.A2(n_1608),
.B1(n_1586),
.B2(n_1595),
.C(n_1597),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1628),
.A2(n_1453),
.B1(n_1523),
.B2(n_1579),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1638),
.B(n_1576),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1622),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1627),
.B(n_1589),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1662),
.Y(n_1672)
);

AOI211x1_ASAP7_75t_SL g1673 ( 
.A1(n_1652),
.A2(n_1642),
.B(n_1640),
.C(n_1632),
.Y(n_1673)
);

NAND2x1p5_ASAP7_75t_L g1674 ( 
.A(n_1668),
.B(n_1628),
.Y(n_1674)
);

OAI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1655),
.A2(n_1628),
.B1(n_1625),
.B2(n_1638),
.C(n_1629),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1656),
.A2(n_1625),
.B(n_1629),
.Y(n_1676)
);

AOI322xp5_ASAP7_75t_L g1677 ( 
.A1(n_1663),
.A2(n_1658),
.A3(n_1664),
.B1(n_1671),
.B2(n_1667),
.C1(n_1650),
.C2(n_1661),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1666),
.B(n_1656),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1653),
.A2(n_1639),
.B1(n_1641),
.B2(n_1612),
.C(n_1614),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1647),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1651),
.B(n_1612),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1648),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1669),
.A2(n_1614),
.B1(n_1624),
.B2(n_1631),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1654),
.Y(n_1684)
);

OAI32xp33_ASAP7_75t_L g1685 ( 
.A1(n_1660),
.A2(n_1636),
.A3(n_1641),
.B1(n_1630),
.B2(n_1639),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1667),
.A2(n_1642),
.B(n_1640),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1649),
.B(n_1636),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1662),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1659),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1670),
.B(n_1630),
.Y(n_1690)
);

AOI322xp5_ASAP7_75t_L g1691 ( 
.A1(n_1665),
.A2(n_1505),
.A3(n_1511),
.B1(n_1576),
.B2(n_1624),
.C1(n_1631),
.C2(n_1604),
.Y(n_1691)
);

OAI322xp33_ASAP7_75t_L g1692 ( 
.A1(n_1686),
.A2(n_1657),
.A3(n_1660),
.B1(n_1571),
.B2(n_1591),
.C1(n_1573),
.C2(n_1575),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1689),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1681),
.B(n_1587),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1687),
.Y(n_1695)
);

INVxp67_ASAP7_75t_SL g1696 ( 
.A(n_1674),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1674),
.B(n_1587),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1672),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1684),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1688),
.B(n_1588),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1680),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1695),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1699),
.B(n_1676),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1696),
.A2(n_1675),
.B1(n_1673),
.B2(n_1677),
.C(n_1678),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1698),
.B(n_1683),
.Y(n_1705)
);

NOR3xp33_ASAP7_75t_L g1706 ( 
.A(n_1693),
.B(n_1675),
.C(n_1682),
.Y(n_1706)
);

NAND4xp25_ASAP7_75t_L g1707 ( 
.A(n_1700),
.B(n_1691),
.C(n_1690),
.D(n_1685),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1693),
.B(n_1690),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1697),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1701),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1704),
.A2(n_1697),
.B1(n_1679),
.B2(n_1694),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1709),
.A2(n_1692),
.B1(n_1694),
.B2(n_1595),
.C(n_1608),
.Y(n_1712)
);

O2A1O1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1703),
.A2(n_1607),
.B(n_1588),
.C(n_1593),
.Y(n_1713)
);

NAND4xp25_ASAP7_75t_L g1714 ( 
.A(n_1707),
.B(n_1430),
.C(n_1453),
.D(n_1448),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1708),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1715),
.A2(n_1706),
.B(n_1705),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1711),
.A2(n_1702),
.B1(n_1710),
.B2(n_1593),
.Y(n_1717)
);

NAND4xp25_ASAP7_75t_L g1718 ( 
.A(n_1714),
.B(n_1453),
.C(n_1448),
.D(n_1602),
.Y(n_1718)
);

OAI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1712),
.A2(n_1575),
.B1(n_1600),
.B2(n_1597),
.C(n_1603),
.Y(n_1719)
);

OAI211xp5_ASAP7_75t_L g1720 ( 
.A1(n_1713),
.A2(n_1575),
.B(n_1600),
.C(n_1531),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1715),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1721),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1716),
.B(n_1720),
.Y(n_1723)
);

NOR3xp33_ASAP7_75t_L g1724 ( 
.A(n_1717),
.B(n_1448),
.C(n_1603),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1718),
.Y(n_1725)
);

OA22x2_ASAP7_75t_L g1726 ( 
.A1(n_1719),
.A2(n_1603),
.B1(n_1533),
.B2(n_1504),
.Y(n_1726)
);

NAND4xp75_ASAP7_75t_L g1727 ( 
.A(n_1723),
.B(n_1533),
.C(n_1538),
.D(n_1399),
.Y(n_1727)
);

NAND3x1_ASAP7_75t_L g1728 ( 
.A(n_1722),
.B(n_1559),
.C(n_1556),
.Y(n_1728)
);

NOR3xp33_ASAP7_75t_SL g1729 ( 
.A(n_1725),
.B(n_1392),
.C(n_1399),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1729),
.A2(n_1724),
.B1(n_1726),
.B2(n_1392),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1730),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1731),
.A2(n_1727),
.B1(n_1728),
.B2(n_1533),
.Y(n_1732)
);

XOR2xp5_ASAP7_75t_L g1733 ( 
.A(n_1731),
.B(n_1445),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1733),
.A2(n_1591),
.B(n_1556),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1732),
.B(n_1399),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1531),
.B1(n_1533),
.B2(n_1504),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1734),
.A2(n_1504),
.B1(n_1399),
.B2(n_1405),
.Y(n_1737)
);

AO21x2_ASAP7_75t_L g1738 ( 
.A1(n_1737),
.A2(n_1568),
.B(n_1564),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1738),
.B(n_1736),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1739),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_R g1741 ( 
.A1(n_1740),
.A2(n_1405),
.B1(n_1399),
.B2(n_1518),
.C(n_1520),
.Y(n_1741)
);

AOI211xp5_ASAP7_75t_L g1742 ( 
.A1(n_1741),
.A2(n_1481),
.B(n_1438),
.C(n_1405),
.Y(n_1742)
);


endmodule