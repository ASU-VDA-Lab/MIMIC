module real_aes_4258_n_3 (n_0, n_2, n_1, n_3);
input n_0;
input n_2;
input n_1;
output n_3;
wire n_4;
wire n_5;
wire n_7;
wire n_8;
wire n_6;
wire n_9;
wire n_10;
INVx2_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
HB1xp67_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
AND2x4_ASAP7_75t_L g7 ( .A(n_1), .B(n_8), .Y(n_7) );
HB1xp67_ASAP7_75t_L g6 ( .A(n_2), .Y(n_6) );
INVx1_ASAP7_75t_L g8 ( .A(n_2), .Y(n_8) );
A2O1A1Ixp33_ASAP7_75t_L g3 ( .A1(n_4), .A2(n_6), .B(n_7), .C(n_9), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_5), .Y(n_4) );
HB1xp67_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
endmodule