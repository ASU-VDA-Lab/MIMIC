module fake_jpeg_418_n_216 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_16),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_66),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_54),
.B1(n_65),
.B2(n_63),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_54),
.B1(n_79),
.B2(n_83),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_94),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_63),
.B1(n_68),
.B2(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_79),
.B1(n_74),
.B2(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_68),
.B1(n_57),
.B2(n_77),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_73),
.B1(n_74),
.B2(n_62),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_102),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_103),
.Y(n_139)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_59),
.B1(n_26),
.B2(n_27),
.Y(n_141)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_87),
.B1(n_99),
.B2(n_93),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_118),
.B1(n_100),
.B2(n_78),
.Y(n_122)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_115),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_59),
.B(n_69),
.Y(n_136)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_87),
.B1(n_73),
.B2(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_56),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_137),
.B(n_7),
.C(n_9),
.D(n_10),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_141),
.B1(n_1),
.B2(n_2),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_127),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_96),
.B(n_76),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_132),
.B(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_138),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_75),
.B(n_70),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_52),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_59),
.C(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_0),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_107),
.B1(n_109),
.B2(n_5),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_141),
.B1(n_12),
.B2(n_13),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_164),
.B1(n_155),
.B2(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_147),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_2),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_7),
.B(n_8),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_11),
.B(n_12),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_156),
.A2(n_163),
.B(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_9),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_50),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_136),
.C(n_137),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_171),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_144),
.B1(n_18),
.B2(n_19),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_17),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_30),
.C(n_44),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_20),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_173),
.B(n_183),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_14),
.B(n_15),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_178),
.B(n_28),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_47),
.B(n_32),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_31),
.C(n_41),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_166),
.A2(n_167),
.B1(n_181),
.B2(n_142),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_189),
.B1(n_190),
.B2(n_192),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_182),
.B(n_156),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_187),
.B(n_188),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_166),
.A2(n_33),
.B1(n_37),
.B2(n_36),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_193),
.B1(n_178),
.B2(n_171),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_168),
.B1(n_166),
.B2(n_180),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_200),
.B1(n_198),
.B2(n_197),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_175),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_201),
.Y(n_203)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_184),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_179),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_177),
.B1(n_176),
.B2(n_190),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_183),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_194),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_202),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_174),
.B1(n_201),
.B2(n_172),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_209),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_211),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_203),
.B(n_34),
.Y(n_213)
);

AO21x2_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_35),
.B(n_42),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_21),
.B(n_22),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_22),
.Y(n_216)
);


endmodule