module fake_jpeg_883_n_689 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_689);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_689;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_672;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_112),
.Y(n_134)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_65),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_66),
.B(n_118),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_79),
.Y(n_183)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_80),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_83),
.Y(n_220)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g221 ( 
.A(n_84),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_85),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_86),
.B(n_17),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g217 ( 
.A(n_88),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_89),
.Y(n_185)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_96),
.Y(n_201)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

BUFx12f_ASAP7_75t_SL g98 ( 
.A(n_32),
.Y(n_98)
);

CKINVDCx9p33_ASAP7_75t_R g184 ( 
.A(n_98),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_103),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_104),
.Y(n_213)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_24),
.B(n_17),
.C(n_16),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_58),
.C(n_38),
.Y(n_179)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_24),
.B(n_17),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_20),
.Y(n_113)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_44),
.B(n_17),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_33),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_39),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_121),
.B(n_123),
.Y(n_192)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_30),
.Y(n_128)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_133),
.B(n_186),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_135),
.B(n_171),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_57),
.B(n_54),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_136),
.A2(n_211),
.B(n_2),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_59),
.A2(n_33),
.B1(n_51),
.B2(n_41),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_145),
.A2(n_172),
.B1(n_197),
.B2(n_209),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_85),
.A2(n_56),
.B1(n_45),
.B2(n_40),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_147),
.A2(n_152),
.B1(n_153),
.B2(n_174),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_61),
.A2(n_33),
.B1(n_51),
.B2(n_41),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_99),
.A2(n_31),
.B1(n_51),
.B2(n_41),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_30),
.B(n_57),
.C(n_46),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g268 ( 
.A1(n_157),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_160),
.B(n_180),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_31),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_89),
.A2(n_56),
.B1(n_45),
.B2(n_40),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_91),
.A2(n_56),
.B1(n_45),
.B2(n_40),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_62),
.A2(n_58),
.B1(n_38),
.B2(n_31),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_176),
.A2(n_178),
.B1(n_182),
.B2(n_198),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_127),
.A2(n_38),
.B1(n_58),
.B2(n_34),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_179),
.B(n_8),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_88),
.B(n_118),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_72),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_34),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_114),
.B(n_36),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_203),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_125),
.B(n_36),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_195),
.B(n_1),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_67),
.A2(n_74),
.B1(n_78),
.B2(n_69),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_94),
.A2(n_35),
.B1(n_54),
.B2(n_50),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_104),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_115),
.B(n_35),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_206),
.B(n_214),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_83),
.A2(n_92),
.B1(n_46),
.B2(n_54),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_208),
.A2(n_219),
.B1(n_222),
.B2(n_5),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_107),
.A2(n_57),
.B1(n_50),
.B2(n_47),
.Y(n_209)
);

HAxp5_ASAP7_75t_SL g211 ( 
.A(n_96),
.B(n_14),
.CON(n_211),
.SN(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_101),
.B(n_50),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_102),
.A2(n_47),
.B1(n_46),
.B2(n_14),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_112),
.A2(n_47),
.B1(n_13),
.B2(n_11),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_159),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_225),
.B(n_228),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_159),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_226),
.Y(n_345)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_227),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_184),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_230),
.B(n_241),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_134),
.B(n_1),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_231),
.B(n_256),
.Y(n_322)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_232),
.Y(n_330)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_130),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_233),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_13),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_236),
.Y(n_357)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_216),
.Y(n_237)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_237),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g238 ( 
.A(n_216),
.Y(n_238)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_238),
.Y(n_362)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_141),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_242),
.Y(n_307)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_155),
.Y(n_243)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_243),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_146),
.Y(n_244)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_244),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_172),
.A2(n_147),
.B1(n_174),
.B2(n_187),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_245),
.A2(n_257),
.B1(n_284),
.B2(n_153),
.Y(n_310)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_143),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_246),
.B(n_255),
.Y(n_346)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_130),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_247),
.Y(n_347)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_161),
.Y(n_248)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_248),
.Y(n_338)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_142),
.Y(n_249)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_249),
.Y(n_336)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_158),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_250),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g251 ( 
.A(n_215),
.B(n_1),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_251),
.A2(n_254),
.B(n_264),
.Y(n_312)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_252),
.Y(n_339)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_253),
.Y(n_361)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_156),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_150),
.B(n_2),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_191),
.A2(n_13),
.B1(n_11),
.B2(n_4),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_169),
.Y(n_258)
);

INVx6_ASAP7_75t_SL g313 ( 
.A(n_258),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_181),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_259),
.A2(n_273),
.B1(n_274),
.B2(n_287),
.Y(n_352)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_260),
.Y(n_358)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_189),
.Y(n_261)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_261),
.Y(n_365)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_262),
.B(n_265),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_175),
.B(n_137),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_263),
.B(n_266),
.Y(n_329)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_223),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_138),
.B(n_2),
.Y(n_266)
);

AO22x1_ASAP7_75t_L g334 ( 
.A1(n_268),
.A2(n_303),
.B1(n_212),
.B2(n_213),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_192),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_269),
.B(n_277),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_146),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_270),
.B(n_271),
.Y(n_360)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_142),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_272),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_131),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_275),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_132),
.B(n_6),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_193),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_278),
.Y(n_315)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_154),
.Y(n_280)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_154),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_281),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_198),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_282),
.A2(n_298),
.B1(n_217),
.B2(n_224),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_183),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_283),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_163),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_173),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_285),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_286),
.B(n_295),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_131),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_166),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_173),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_289),
.Y(n_348)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_290),
.Y(n_363)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_291),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_196),
.A2(n_9),
.B1(n_10),
.B2(n_165),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_296),
.Y(n_356)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_162),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_162),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_139),
.B(n_10),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_167),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_177),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_299),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g298 ( 
.A1(n_182),
.A2(n_10),
.B1(n_208),
.B2(n_178),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_140),
.A2(n_218),
.B1(n_200),
.B2(n_166),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_300),
.A2(n_301),
.B1(n_304),
.B2(n_169),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_148),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_157),
.B(n_211),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_148),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_210),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_151),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_229),
.A2(n_205),
.B1(n_204),
.B2(n_201),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_306),
.A2(n_320),
.B1(n_333),
.B2(n_284),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_310),
.A2(n_317),
.B1(n_319),
.B2(n_327),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_219),
.B1(n_185),
.B2(n_163),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_279),
.A2(n_240),
.B1(n_286),
.B2(n_267),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_244),
.A2(n_201),
.B1(n_205),
.B2(n_204),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_324),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_286),
.A2(n_199),
.B1(n_185),
.B2(n_213),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_303),
.A2(n_224),
.B1(n_199),
.B2(n_164),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_334),
.B(n_351),
.Y(n_385)
);

OR2x2_ASAP7_75t_SL g335 ( 
.A(n_303),
.B(n_217),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_335),
.A2(n_236),
.B(n_292),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_343),
.A2(n_359),
.B1(n_295),
.B2(n_258),
.Y(n_388)
);

AO22x1_ASAP7_75t_L g344 ( 
.A1(n_303),
.A2(n_149),
.B1(n_151),
.B2(n_164),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_350),
.B(n_301),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_256),
.B(n_170),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_266),
.B(n_170),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_366),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_251),
.A2(n_239),
.B1(n_298),
.B2(n_235),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_251),
.B(n_263),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_367),
.Y(n_420)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_308),
.Y(n_368)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_368),
.Y(n_431)
);

MAJx2_ASAP7_75t_L g369 ( 
.A(n_319),
.B(n_302),
.C(n_234),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_384),
.C(n_390),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_370),
.A2(n_349),
.B(n_324),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g371 ( 
.A1(n_359),
.A2(n_231),
.B(n_268),
.C(n_295),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_371),
.A2(n_331),
.B(n_348),
.C(n_328),
.Y(n_444)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_373),
.Y(n_432)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_374),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_375),
.B(n_391),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_322),
.B(n_252),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_377),
.B(n_378),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_313),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_379),
.A2(n_410),
.B1(n_413),
.B2(n_393),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_313),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_382),
.Y(n_419)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_341),
.Y(n_381)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_322),
.B(n_260),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_365),
.Y(n_383)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_383),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_335),
.B(n_262),
.C(n_290),
.Y(n_384)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_396),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_388),
.A2(n_397),
.B1(n_408),
.B2(n_345),
.Y(n_436)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_325),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_389),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_329),
.B(n_248),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_243),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_317),
.A2(n_226),
.B(n_283),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_392),
.A2(n_372),
.B(n_409),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_308),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_394),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_355),
.B(n_281),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_400),
.C(n_358),
.Y(n_428)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_334),
.A2(n_249),
.B1(n_291),
.B2(n_233),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_342),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_399),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_250),
.C(n_299),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_310),
.A2(n_261),
.B1(n_253),
.B2(n_232),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_401),
.A2(n_409),
.B1(n_411),
.B2(n_414),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_403),
.Y(n_441)
);

INVxp33_ASAP7_75t_L g403 ( 
.A(n_342),
.Y(n_403)
);

INVx3_ASAP7_75t_SL g404 ( 
.A(n_325),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_404),
.Y(n_429)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_412),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_351),
.B(n_304),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_407),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_280),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_334),
.A2(n_247),
.B1(n_272),
.B2(n_271),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_344),
.A2(n_275),
.B1(n_237),
.B2(n_238),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_323),
.A2(n_276),
.B1(n_242),
.B2(n_294),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_344),
.A2(n_227),
.B1(n_293),
.B2(n_343),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_358),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_323),
.A2(n_332),
.B1(n_314),
.B2(n_309),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_312),
.A2(n_366),
.B1(n_327),
.B2(n_360),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_385),
.A2(n_352),
.B(n_356),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_415),
.A2(n_425),
.B(n_437),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_332),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_424),
.B(n_433),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_372),
.A2(n_357),
.B1(n_360),
.B2(n_326),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_428),
.B(n_364),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_376),
.A2(n_309),
.B1(n_315),
.B2(n_336),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_430),
.A2(n_435),
.B1(n_454),
.B2(n_396),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_367),
.B(n_390),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_376),
.A2(n_315),
.B1(n_336),
.B2(n_349),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_436),
.A2(n_445),
.B1(n_450),
.B2(n_408),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_373),
.B(n_346),
.Y(n_438)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_442),
.C(n_444),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_386),
.B(n_338),
.C(n_346),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_440),
.B(n_446),
.C(n_364),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_374),
.B(n_331),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_443),
.A2(n_370),
.B(n_393),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_385),
.A2(n_388),
.B1(n_401),
.B2(n_392),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_386),
.B(n_395),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_414),
.A2(n_348),
.B1(n_354),
.B2(n_337),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_406),
.B(n_363),
.Y(n_452)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_452),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_407),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_453),
.B(n_412),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_397),
.A2(n_336),
.B1(n_328),
.B2(n_337),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_369),
.Y(n_455)
);

XNOR2x2_ASAP7_75t_L g510 ( 
.A(n_455),
.B(n_446),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_457),
.A2(n_466),
.B(n_470),
.Y(n_501)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_458),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_460),
.A2(n_421),
.B1(n_416),
.B2(n_454),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_423),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_461),
.B(n_462),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_423),
.Y(n_462)
);

NOR2x1_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_384),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_477),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_445),
.A2(n_371),
.B1(n_411),
.B2(n_379),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_465),
.A2(n_469),
.B1(n_473),
.B2(n_479),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_SL g466 ( 
.A(n_417),
.B(n_400),
.C(n_381),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_451),
.Y(n_467)
);

INVx11_ASAP7_75t_L g504 ( 
.A(n_467),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_415),
.A2(n_405),
.B1(n_383),
.B2(n_387),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_444),
.A2(n_378),
.B(n_380),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_471),
.A2(n_420),
.B1(n_434),
.B2(n_432),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_439),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_472),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_415),
.A2(n_404),
.B1(n_389),
.B2(n_399),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_451),
.Y(n_474)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_417),
.B(n_338),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_484),
.C(n_487),
.Y(n_497)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_448),
.Y(n_476)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_476),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_442),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_402),
.B(n_321),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_478),
.A2(n_486),
.B(n_424),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_427),
.A2(n_404),
.B1(n_368),
.B2(n_347),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_481),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_439),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_488),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_427),
.A2(n_337),
.B1(n_347),
.B2(n_361),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_483),
.A2(n_436),
.B1(n_460),
.B2(n_454),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_363),
.Y(n_485)
);

CKINVDCx14_ASAP7_75t_R g506 ( 
.A(n_485),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_437),
.A2(n_321),
.B(n_345),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_316),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_452),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_435),
.A2(n_354),
.B1(n_347),
.B2(n_307),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_489),
.A2(n_447),
.B1(n_429),
.B2(n_426),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_428),
.C(n_446),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_438),
.B(n_307),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_491),
.B(n_492),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_441),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_470),
.A2(n_443),
.B(n_422),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_494),
.A2(n_505),
.B(n_516),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_499),
.A2(n_509),
.B1(n_515),
.B2(n_519),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_522),
.C(n_525),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_503),
.A2(n_480),
.B(n_456),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g505 ( 
.A1(n_459),
.A2(n_435),
.B(n_430),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_471),
.A2(n_430),
.B1(n_450),
.B2(n_421),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_455),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_511),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_465),
.A2(n_432),
.B1(n_434),
.B2(n_420),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_477),
.A2(n_416),
.B1(n_433),
.B2(n_419),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_468),
.A2(n_441),
.B1(n_418),
.B2(n_419),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_459),
.A2(n_418),
.B(n_449),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_491),
.Y(n_517)
);

INVx11_ASAP7_75t_L g551 ( 
.A(n_517),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_468),
.A2(n_440),
.B1(n_428),
.B2(n_447),
.Y(n_521)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_521),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_475),
.B(n_487),
.C(n_484),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_478),
.A2(n_440),
.B1(n_431),
.B2(n_318),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_523),
.A2(n_509),
.B1(n_469),
.B2(n_473),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_458),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_463),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_475),
.B(n_431),
.C(n_330),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_457),
.A2(n_325),
.B(n_330),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_526),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_480),
.B(n_354),
.Y(n_527)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_527),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_488),
.A2(n_311),
.B1(n_318),
.B2(n_463),
.Y(n_528)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_528),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_530),
.B(n_547),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_461),
.Y(n_532)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_532),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_506),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_536),
.B(n_543),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_514),
.B(n_462),
.Y(n_538)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_538),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_529),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_539),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_540),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_500),
.B(n_490),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_541),
.B(n_542),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_500),
.B(n_464),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_529),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_496),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_544),
.B(n_549),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g577 ( 
.A(n_545),
.B(n_501),
.Y(n_577)
);

AO32x1_ASAP7_75t_L g547 ( 
.A1(n_503),
.A2(n_486),
.A3(n_464),
.B1(n_455),
.B2(n_485),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_496),
.B(n_467),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_548),
.B(n_550),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_524),
.B(n_474),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_502),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_506),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_552),
.A2(n_559),
.B1(n_560),
.B2(n_562),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_529),
.B(n_492),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_553),
.B(n_554),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_521),
.B(n_498),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_555),
.A2(n_528),
.B(n_527),
.Y(n_590)
);

BUFx12_ASAP7_75t_L g558 ( 
.A(n_526),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_558),
.Y(n_591)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_502),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_518),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_518),
.B(n_476),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_561),
.B(n_563),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_520),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_498),
.B(n_481),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_535),
.A2(n_494),
.B1(n_493),
.B2(n_499),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_564),
.A2(n_571),
.B1(n_580),
.B2(n_586),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_530),
.A2(n_516),
.B(n_505),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_570),
.A2(n_551),
.B1(n_546),
.B2(n_504),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_535),
.A2(n_493),
.B1(n_523),
.B2(n_515),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_541),
.B(n_522),
.C(n_497),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_572),
.B(n_582),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_534),
.B(n_522),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_574),
.B(n_575),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_534),
.B(n_497),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_577),
.B(n_547),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_542),
.B(n_497),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_578),
.B(n_579),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_533),
.B(n_466),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_538),
.A2(n_523),
.B1(n_520),
.B2(n_513),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_533),
.B(n_525),
.C(n_501),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_545),
.B(n_525),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_584),
.B(n_590),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_562),
.A2(n_556),
.B1(n_560),
.B2(n_532),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_555),
.B(n_510),
.C(n_495),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_589),
.B(n_557),
.C(n_556),
.Y(n_593)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_583),
.Y(n_592)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_592),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_593),
.B(n_584),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_581),
.B(n_539),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_595),
.B(n_596),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_566),
.A2(n_548),
.B1(n_552),
.B2(n_536),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_583),
.B(n_576),
.Y(n_597)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_597),
.Y(n_635)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_587),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_598),
.B(n_601),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_576),
.B(n_563),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_600),
.Y(n_633)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_587),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_569),
.B(n_561),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_602),
.B(n_604),
.Y(n_631)
);

AND2x2_ASAP7_75t_SL g604 ( 
.A(n_564),
.B(n_531),
.Y(n_604)
);

FAx1_ASAP7_75t_L g605 ( 
.A(n_565),
.B(n_547),
.CI(n_510),
.CON(n_605),
.SN(n_605)
);

O2A1O1Ixp33_ASAP7_75t_L g628 ( 
.A1(n_605),
.A2(n_614),
.B(n_537),
.C(n_551),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_574),
.B(n_557),
.C(n_546),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_606),
.B(n_615),
.C(n_582),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_607),
.B(n_606),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_573),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_608),
.B(n_609),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_581),
.Y(n_609)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_585),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_611),
.A2(n_613),
.B1(n_504),
.B2(n_559),
.Y(n_632)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_567),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_575),
.B(n_540),
.C(n_531),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g618 ( 
.A1(n_612),
.A2(n_565),
.B1(n_566),
.B2(n_570),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_618),
.B(n_622),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_620),
.B(n_594),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_605),
.A2(n_590),
.B(n_589),
.Y(n_621)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_621),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_610),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_623),
.B(n_603),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_612),
.A2(n_537),
.B1(n_588),
.B2(n_591),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_624),
.B(n_625),
.Y(n_640)
);

FAx1_ASAP7_75t_SL g625 ( 
.A(n_605),
.B(n_577),
.CI(n_607),
.CON(n_625),
.SN(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_596),
.A2(n_586),
.B(n_571),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_626),
.A2(n_602),
.B1(n_597),
.B2(n_600),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_627),
.B(n_629),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_628),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_599),
.B(n_579),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_593),
.B(n_572),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_630),
.B(n_632),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_638),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_622),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g659 ( 
.A(n_639),
.B(n_642),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g642 ( 
.A(n_630),
.B(n_623),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_627),
.B(n_615),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_644),
.B(n_649),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_634),
.B(n_604),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g652 ( 
.A(n_646),
.B(n_651),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_SL g647 ( 
.A1(n_626),
.A2(n_613),
.B1(n_604),
.B2(n_592),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_647),
.B(n_650),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_620),
.B(n_594),
.Y(n_649)
);

FAx1_ASAP7_75t_SL g651 ( 
.A(n_618),
.B(n_580),
.CI(n_504),
.CON(n_651),
.SN(n_651)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_641),
.A2(n_617),
.B(n_628),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_653),
.A2(n_662),
.B(n_663),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_648),
.B(n_619),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_654),
.B(n_658),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_642),
.B(n_603),
.C(n_636),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_656),
.B(n_657),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_643),
.B(n_624),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_648),
.B(n_633),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_637),
.A2(n_616),
.B(n_631),
.Y(n_662)
);

CKINVDCx14_ASAP7_75t_R g663 ( 
.A(n_640),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_639),
.B(n_649),
.C(n_644),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_664),
.B(n_621),
.C(n_635),
.Y(n_669)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_661),
.B(n_629),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_665),
.B(n_668),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_659),
.B(n_645),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_669),
.B(n_670),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g670 ( 
.A(n_659),
.B(n_578),
.C(n_568),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_655),
.Y(n_671)
);

AO21x1_ASAP7_75t_L g679 ( 
.A1(n_671),
.A2(n_666),
.B(n_665),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_656),
.A2(n_651),
.B(n_625),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_673),
.A2(n_652),
.B(n_664),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_675),
.B(n_676),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_672),
.B(n_661),
.C(n_660),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_667),
.A2(n_625),
.B(n_550),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_678),
.B(n_679),
.Y(n_682)
);

OAI321xp33_ASAP7_75t_L g680 ( 
.A1(n_674),
.A2(n_677),
.A3(n_669),
.B1(n_508),
.B2(n_507),
.C(n_512),
.Y(n_680)
);

A2O1A1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_680),
.A2(n_495),
.B(n_489),
.C(n_511),
.Y(n_684)
);

A2O1A1O1Ixp25_ASAP7_75t_L g683 ( 
.A1(n_682),
.A2(n_670),
.B(n_568),
.C(n_508),
.D(n_507),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_683),
.A2(n_684),
.B(n_519),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_685),
.A2(n_519),
.B1(n_681),
.B2(n_483),
.C(n_479),
.Y(n_686)
);

NAND2x1_ASAP7_75t_SL g687 ( 
.A(n_686),
.B(n_558),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_687),
.B(n_558),
.Y(n_688)
);

OAI21xp33_ASAP7_75t_L g689 ( 
.A1(n_688),
.A2(n_558),
.B(n_311),
.Y(n_689)
);


endmodule