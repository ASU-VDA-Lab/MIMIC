module real_aes_6778_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_175;
wire n_168;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g527 ( .A(n_1), .Y(n_527) );
INVx1_ASAP7_75t_L g149 ( .A(n_2), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_3), .A2(n_37), .B1(n_174), .B2(n_473), .Y(n_496) );
AOI21xp33_ASAP7_75t_L g181 ( .A1(n_4), .A2(n_165), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_5), .B(n_163), .Y(n_539) );
AND2x6_ASAP7_75t_L g142 ( .A(n_6), .B(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_7), .A2(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_8), .B(n_38), .Y(n_439) );
INVx1_ASAP7_75t_L g187 ( .A(n_9), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_10), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g134 ( .A(n_11), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_12), .B(n_155), .Y(n_482) );
INVx1_ASAP7_75t_L g258 ( .A(n_13), .Y(n_258) );
INVx1_ASAP7_75t_L g521 ( .A(n_14), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_15), .B(n_130), .Y(n_510) );
AO32x2_ASAP7_75t_L g494 ( .A1(n_16), .A2(n_129), .A3(n_163), .B1(n_475), .B2(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_17), .B(n_174), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_18), .B(n_170), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_19), .B(n_130), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_20), .A2(n_49), .B1(n_174), .B2(n_473), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_21), .B(n_165), .Y(n_215) );
OAI222xp33_ASAP7_75t_L g444 ( .A1(n_22), .A2(n_445), .B1(n_728), .B2(n_729), .C1(n_734), .C2(n_738), .Y(n_444) );
INVx1_ASAP7_75t_L g728 ( .A(n_22), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_23), .A2(n_74), .B1(n_155), .B2(n_174), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_24), .B(n_174), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_25), .B(n_177), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_26), .A2(n_256), .B(n_257), .C(n_259), .Y(n_255) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_27), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_28), .B(n_160), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_29), .B(n_153), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_30), .A2(n_100), .B1(n_113), .B2(n_739), .Y(n_99) );
INVx1_ASAP7_75t_L g202 ( .A(n_31), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_32), .B(n_160), .Y(n_466) );
INVx2_ASAP7_75t_L g140 ( .A(n_33), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_34), .B(n_174), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_35), .B(n_160), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_36), .A2(n_142), .B(n_145), .C(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_38), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g200 ( .A(n_39), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_40), .B(n_153), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_41), .B(n_174), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_42), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_43), .A2(n_84), .B1(n_222), .B2(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_44), .B(n_174), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_45), .B(n_174), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_46), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_47), .B(n_526), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_48), .B(n_165), .Y(n_246) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_50), .A2(n_60), .B1(n_155), .B2(n_174), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_51), .A2(n_145), .B1(n_155), .B2(n_198), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_52), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_53), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_54), .B(n_174), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g136 ( .A(n_55), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_56), .B(n_174), .Y(n_547) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_57), .A2(n_173), .B(n_185), .C(n_186), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_58), .Y(n_235) );
INVx1_ASAP7_75t_L g183 ( .A(n_59), .Y(n_183) );
INVx1_ASAP7_75t_L g143 ( .A(n_61), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_62), .B(n_174), .Y(n_528) );
INVx1_ASAP7_75t_L g133 ( .A(n_63), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
AO32x2_ASAP7_75t_L g470 ( .A1(n_65), .A2(n_163), .A3(n_238), .B1(n_471), .B2(n_475), .Y(n_470) );
INVx1_ASAP7_75t_L g546 ( .A(n_66), .Y(n_546) );
INVx1_ASAP7_75t_L g461 ( .A(n_67), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_SL g169 ( .A1(n_68), .A2(n_170), .B(n_171), .C(n_173), .Y(n_169) );
INVxp67_ASAP7_75t_L g172 ( .A(n_69), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_70), .B(n_155), .Y(n_462) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_72), .Y(n_205) );
INVx1_ASAP7_75t_L g228 ( .A(n_73), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_75), .A2(n_142), .B(n_145), .C(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_76), .B(n_473), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_77), .B(n_155), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_78), .B(n_150), .Y(n_218) );
INVx2_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_80), .B(n_170), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_81), .B(n_155), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_82), .A2(n_142), .B(n_145), .C(n_148), .Y(n_144) );
INVx2_ASAP7_75t_L g109 ( .A(n_83), .Y(n_109) );
OR2x2_ASAP7_75t_L g436 ( .A(n_83), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g449 ( .A(n_83), .B(n_438), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_85), .A2(n_98), .B1(n_155), .B2(n_156), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_86), .A2(n_120), .B1(n_121), .B2(n_434), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_86), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_87), .B(n_160), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_88), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_89), .A2(n_142), .B(n_145), .C(n_241), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_90), .Y(n_248) );
INVx1_ASAP7_75t_L g168 ( .A(n_91), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g254 ( .A(n_92), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_93), .B(n_150), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_94), .B(n_155), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_95), .B(n_163), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_96), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_97), .A2(n_165), .B(n_166), .Y(n_164) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx3_ASAP7_75t_SL g739 ( .A(n_102), .Y(n_739) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g438 ( .A(n_108), .B(n_439), .Y(n_438) );
OR2x2_ASAP7_75t_L g727 ( .A(n_109), .B(n_438), .Y(n_727) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_109), .B(n_437), .Y(n_737) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_443), .Y(n_113) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_114), .A2(n_440), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_435), .B(n_440), .Y(n_118) );
INVx1_ASAP7_75t_L g434 ( .A(n_121), .Y(n_434) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_122), .A2(n_447), .B1(n_450), .B2(n_725), .Y(n_446) );
INVx1_ASAP7_75t_L g732 ( .A(n_122), .Y(n_732) );
NAND2x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_350), .Y(n_122) );
NOR5xp2_ASAP7_75t_L g123 ( .A(n_124), .B(n_273), .C(n_305), .D(n_320), .E(n_337), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_189), .B(n_210), .C(n_261), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_126), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_126), .B(n_325), .Y(n_388) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_127), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_127), .B(n_207), .Y(n_274) );
AND2x2_ASAP7_75t_L g315 ( .A(n_127), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_127), .B(n_284), .Y(n_319) );
OR2x2_ASAP7_75t_L g356 ( .A(n_127), .B(n_195), .Y(n_356) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g194 ( .A(n_128), .B(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g264 ( .A(n_128), .Y(n_264) );
OR2x2_ASAP7_75t_L g427 ( .A(n_128), .B(n_267), .Y(n_427) );
AO21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_135), .B(n_157), .Y(n_128) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_129), .A2(n_196), .B(n_204), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_129), .B(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g223 ( .A(n_129), .Y(n_223) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_130), .Y(n_163) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_131), .B(n_132), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
OAI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_144), .Y(n_135) );
OAI22xp33_ASAP7_75t_L g196 ( .A1(n_137), .A2(n_175), .B1(n_197), .B2(n_203), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_137), .A2(n_228), .B(n_229), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
AND2x4_ASAP7_75t_L g165 ( .A(n_138), .B(n_142), .Y(n_165) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g526 ( .A(n_139), .Y(n_526) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_140), .Y(n_156) );
INVx1_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx3_ASAP7_75t_L g151 ( .A(n_141), .Y(n_151) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
INVx1_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_141), .Y(n_199) );
INVx4_ASAP7_75t_SL g175 ( .A(n_142), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_142), .A2(n_460), .B(n_463), .Y(n_459) );
BUFx3_ASAP7_75t_L g475 ( .A(n_142), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_142), .A2(n_480), .B(n_484), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_142), .A2(n_520), .B(n_524), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_142), .A2(n_533), .B(n_536), .Y(n_532) );
INVx5_ASAP7_75t_L g167 ( .A(n_145), .Y(n_167) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
BUFx3_ASAP7_75t_L g222 ( .A(n_146), .Y(n_222) );
INVx1_ASAP7_75t_L g473 ( .A(n_146), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_152), .C(n_154), .Y(n_148) );
O2A1O1Ixp5_ASAP7_75t_SL g460 ( .A1(n_150), .A2(n_173), .B(n_461), .C(n_462), .Y(n_460) );
INVx2_ASAP7_75t_L g497 ( .A(n_150), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_150), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_150), .A2(n_543), .B(n_544), .Y(n_542) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_151), .B(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_151), .B(n_187), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g471 ( .A1(n_151), .A2(n_153), .B1(n_472), .B2(n_474), .Y(n_471) );
INVx2_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
INVx4_ASAP7_75t_L g244 ( .A(n_153), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_153), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_153), .A2(n_497), .B1(n_513), .B2(n_514), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_154), .A2(n_521), .B(n_522), .C(n_523), .Y(n_520) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_159), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_159), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g238 ( .A(n_160), .Y(n_238) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_160), .A2(n_251), .B(n_260), .Y(n_250) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_160), .A2(n_459), .B(n_466), .Y(n_458) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_160), .A2(n_479), .B(n_487), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_161), .A2(n_330), .B1(n_331), .B2(n_334), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_161), .B(n_264), .Y(n_413) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_179), .Y(n_161) );
AND2x2_ASAP7_75t_L g209 ( .A(n_162), .B(n_195), .Y(n_209) );
AND2x2_ASAP7_75t_L g266 ( .A(n_162), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g271 ( .A(n_162), .Y(n_271) );
INVx3_ASAP7_75t_L g284 ( .A(n_162), .Y(n_284) );
OR2x2_ASAP7_75t_L g304 ( .A(n_162), .B(n_267), .Y(n_304) );
AND2x2_ASAP7_75t_L g323 ( .A(n_162), .B(n_180), .Y(n_323) );
BUFx2_ASAP7_75t_L g355 ( .A(n_162), .Y(n_355) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_176), .Y(n_162) );
INVx4_ASAP7_75t_L g178 ( .A(n_163), .Y(n_178) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_163), .A2(n_532), .B(n_539), .Y(n_531) );
BUFx2_ASAP7_75t_L g252 ( .A(n_165), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_169), .C(n_175), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_167), .A2(n_175), .B(n_183), .C(n_184), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_167), .A2(n_175), .B(n_254), .C(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g483 ( .A(n_170), .Y(n_483) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_174), .Y(n_245) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_177), .A2(n_181), .B(n_188), .Y(n_180) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_178), .B(n_225), .Y(n_224) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_178), .B(n_475), .C(n_512), .Y(n_511) );
AO21x1_ASAP7_75t_L g601 ( .A1(n_178), .A2(n_512), .B(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_L g270 ( .A(n_179), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_SL g179 ( .A(n_180), .Y(n_179) );
BUFx2_ASAP7_75t_L g193 ( .A(n_180), .Y(n_193) );
INVx2_ASAP7_75t_L g208 ( .A(n_180), .Y(n_208) );
OR2x2_ASAP7_75t_L g286 ( .A(n_180), .B(n_267), .Y(n_286) );
AND2x2_ASAP7_75t_L g316 ( .A(n_180), .B(n_195), .Y(n_316) );
AND2x2_ASAP7_75t_L g333 ( .A(n_180), .B(n_264), .Y(n_333) );
AND2x2_ASAP7_75t_L g373 ( .A(n_180), .B(n_284), .Y(n_373) );
AND2x2_ASAP7_75t_SL g409 ( .A(n_180), .B(n_209), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_185), .A2(n_485), .B(n_486), .Y(n_484) );
O2A1O1Ixp5_ASAP7_75t_L g545 ( .A1(n_185), .A2(n_525), .B(n_546), .C(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp33_ASAP7_75t_SL g190 ( .A(n_191), .B(n_206), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_194), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_192), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
OAI21xp33_ASAP7_75t_L g347 ( .A1(n_193), .A2(n_209), .B(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_193), .B(n_195), .Y(n_403) );
AND2x2_ASAP7_75t_L g339 ( .A(n_194), .B(n_340), .Y(n_339) );
INVx3_ASAP7_75t_L g267 ( .A(n_195), .Y(n_267) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_195), .Y(n_365) );
OAI22xp5_ASAP7_75t_SL g198 ( .A1(n_199), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_198) );
INVx2_ASAP7_75t_L g201 ( .A(n_199), .Y(n_201) );
INVx4_ASAP7_75t_L g256 ( .A(n_199), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_206), .B(n_264), .Y(n_432) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_207), .A2(n_375), .B1(n_376), .B2(n_381), .Y(n_374) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
AND2x2_ASAP7_75t_L g265 ( .A(n_208), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g303 ( .A(n_208), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g340 ( .A(n_208), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_209), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g394 ( .A(n_209), .Y(n_394) );
CKINVDCx16_ASAP7_75t_R g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_236), .Y(n_211) );
INVx4_ASAP7_75t_L g280 ( .A(n_212), .Y(n_280) );
AND2x2_ASAP7_75t_L g358 ( .A(n_212), .B(n_325), .Y(n_358) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
INVx3_ASAP7_75t_L g277 ( .A(n_213), .Y(n_277) );
AND2x2_ASAP7_75t_L g291 ( .A(n_213), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g295 ( .A(n_213), .Y(n_295) );
INVx2_ASAP7_75t_L g309 ( .A(n_213), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_213), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g366 ( .A(n_213), .B(n_361), .Y(n_366) );
AND2x2_ASAP7_75t_L g431 ( .A(n_213), .B(n_401), .Y(n_431) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_216), .B(n_223), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_220), .A2(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g259 ( .A(n_222), .Y(n_259) );
INVx1_ASAP7_75t_L g233 ( .A(n_223), .Y(n_233) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_223), .A2(n_519), .B(n_529), .Y(n_518) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_223), .A2(n_541), .B(n_548), .Y(n_540) );
AND2x2_ASAP7_75t_L g272 ( .A(n_226), .B(n_250), .Y(n_272) );
INVx2_ASAP7_75t_L g292 ( .A(n_226), .Y(n_292) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_233), .B(n_234), .Y(n_226) );
INVx1_ASAP7_75t_L g297 ( .A(n_236), .Y(n_297) );
AND2x2_ASAP7_75t_L g343 ( .A(n_236), .B(n_291), .Y(n_343) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_249), .Y(n_236) );
INVx2_ASAP7_75t_L g282 ( .A(n_237), .Y(n_282) );
INVx1_ASAP7_75t_L g290 ( .A(n_237), .Y(n_290) );
AND2x2_ASAP7_75t_L g308 ( .A(n_237), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_237), .B(n_292), .Y(n_346) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_247), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_246), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_245), .Y(n_241) );
AND2x2_ASAP7_75t_L g325 ( .A(n_249), .B(n_282), .Y(n_325) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g278 ( .A(n_250), .Y(n_278) );
AND2x2_ASAP7_75t_L g361 ( .A(n_250), .B(n_292), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_256), .B(n_258), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_256), .A2(n_464), .B(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g523 ( .A(n_256), .Y(n_523) );
OAI21xp5_ASAP7_75t_SL g261 ( .A1(n_262), .A2(n_268), .B(n_272), .Y(n_261) );
INVx1_ASAP7_75t_SL g306 ( .A(n_262), .Y(n_306) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_263), .B(n_270), .Y(n_363) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g312 ( .A(n_264), .B(n_267), .Y(n_312) );
AND2x2_ASAP7_75t_L g341 ( .A(n_264), .B(n_285), .Y(n_341) );
OR2x2_ASAP7_75t_L g344 ( .A(n_264), .B(n_304), .Y(n_344) );
AOI222xp33_ASAP7_75t_L g408 ( .A1(n_265), .A2(n_357), .B1(n_409), .B2(n_410), .C1(n_412), .C2(n_414), .Y(n_408) );
BUFx2_ASAP7_75t_L g322 ( .A(n_267), .Y(n_322) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g311 ( .A(n_270), .B(n_312), .Y(n_311) );
INVx3_ASAP7_75t_SL g328 ( .A(n_270), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_270), .B(n_322), .Y(n_382) );
AND2x2_ASAP7_75t_L g317 ( .A(n_272), .B(n_277), .Y(n_317) );
INVx1_ASAP7_75t_L g336 ( .A(n_272), .Y(n_336) );
OAI221xp5_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_275), .B1(n_279), .B2(n_283), .C(n_287), .Y(n_273) );
OR2x2_ASAP7_75t_L g345 ( .A(n_275), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g330 ( .A(n_277), .B(n_300), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_277), .B(n_290), .Y(n_370) );
AND2x2_ASAP7_75t_L g375 ( .A(n_277), .B(n_325), .Y(n_375) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_277), .Y(n_385) );
NAND2x1_ASAP7_75t_SL g396 ( .A(n_277), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g281 ( .A(n_278), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g301 ( .A(n_278), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_278), .B(n_296), .Y(n_327) );
INVx1_ASAP7_75t_L g393 ( .A(n_278), .Y(n_393) );
INVx1_ASAP7_75t_L g368 ( .A(n_279), .Y(n_368) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g380 ( .A(n_280), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g392 ( .A(n_280), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g397 ( .A(n_281), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_281), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g300 ( .A(n_282), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_282), .B(n_292), .Y(n_313) );
INVx1_ASAP7_75t_L g379 ( .A(n_282), .Y(n_379) );
INVx1_ASAP7_75t_L g400 ( .A(n_283), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_293), .B(n_302), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
AND2x2_ASAP7_75t_L g433 ( .A(n_289), .B(n_366), .Y(n_433) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g401 ( .A(n_290), .B(n_361), .Y(n_401) );
AOI32xp33_ASAP7_75t_L g314 ( .A1(n_291), .A2(n_297), .A3(n_315), .B1(n_317), .B2(n_318), .Y(n_314) );
AOI322xp5_ASAP7_75t_L g416 ( .A1(n_291), .A2(n_323), .A3(n_406), .B1(n_417), .B2(n_418), .C1(n_419), .C2(n_421), .Y(n_416) );
INVx2_ASAP7_75t_L g296 ( .A(n_292), .Y(n_296) );
INVx1_ASAP7_75t_L g406 ( .A(n_292), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B1(n_298), .B2(n_299), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_294), .B(n_300), .Y(n_349) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_295), .B(n_361), .Y(n_411) );
INVx1_ASAP7_75t_L g298 ( .A(n_296), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_296), .B(n_325), .Y(n_415) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_304), .B(n_399), .Y(n_398) );
OAI221xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_307), .B1(n_310), .B2(n_313), .C(n_314), .Y(n_305) );
OR2x2_ASAP7_75t_L g326 ( .A(n_307), .B(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g335 ( .A(n_307), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g360 ( .A(n_308), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g364 ( .A(n_318), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OAI221xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_324), .B1(n_326), .B2(n_328), .C(n_329), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_322), .A2(n_353), .B1(n_357), .B2(n_358), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_323), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_323), .Y(n_428) );
INVx1_ASAP7_75t_L g422 ( .A(n_325), .Y(n_422) );
INVx1_ASAP7_75t_SL g357 ( .A(n_326), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_328), .B(n_356), .Y(n_418) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_333), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g399 ( .A(n_333), .Y(n_399) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
OAI221xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_342), .B1(n_344), .B2(n_345), .C(n_347), .Y(n_337) );
NOR2xp33_ASAP7_75t_SL g338 ( .A(n_339), .B(n_341), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_339), .A2(n_357), .B1(n_403), .B2(n_404), .Y(n_402) );
CKINVDCx14_ASAP7_75t_R g342 ( .A(n_343), .Y(n_342) );
OAI21xp33_ASAP7_75t_L g421 ( .A1(n_344), .A2(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR3xp33_ASAP7_75t_SL g350 ( .A(n_351), .B(n_383), .C(n_407), .Y(n_350) );
NAND4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_359), .C(n_367), .D(n_374), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g430 ( .A(n_355), .Y(n_430) );
INVx3_ASAP7_75t_SL g424 ( .A(n_356), .Y(n_424) );
OR2x2_ASAP7_75t_L g429 ( .A(n_356), .B(n_430), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B1(n_364), .B2(n_366), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_361), .B(n_379), .Y(n_420) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI21xp5_ASAP7_75t_SL g367 ( .A1(n_368), .A2(n_369), .B(n_371), .Y(n_367) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI211xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_386), .B(n_389), .C(n_402), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g417 ( .A(n_388), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_394), .B1(n_395), .B2(n_398), .C1(n_400), .C2(n_401), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND4xp25_ASAP7_75t_SL g426 ( .A(n_399), .B(n_427), .C(n_428), .D(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND3xp33_ASAP7_75t_SL g407 ( .A(n_408), .B(n_416), .C(n_425), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_431), .B1(n_432), .B2(n_433), .Y(n_425) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g441 ( .A(n_436), .Y(n_441) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_SL g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g731 ( .A(n_448), .Y(n_731) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g733 ( .A(n_450), .Y(n_733) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_646), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_595), .C(n_637), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_504), .B(n_549), .C(n_571), .Y(n_452) );
OAI211xp5_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_467), .B(n_488), .C(n_499), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_455), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g658 ( .A(n_455), .B(n_575), .Y(n_658) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g560 ( .A(n_456), .B(n_491), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_456), .B(n_478), .Y(n_677) );
INVx1_ASAP7_75t_L g695 ( .A(n_456), .Y(n_695) );
AND2x2_ASAP7_75t_L g704 ( .A(n_456), .B(n_592), .Y(n_704) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g587 ( .A(n_457), .B(n_478), .Y(n_587) );
AND2x2_ASAP7_75t_L g645 ( .A(n_457), .B(n_592), .Y(n_645) );
INVx1_ASAP7_75t_L g689 ( .A(n_457), .Y(n_689) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g566 ( .A(n_458), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g574 ( .A(n_458), .Y(n_574) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_458), .Y(n_614) );
INVxp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_476), .Y(n_468) );
AND2x2_ASAP7_75t_L g553 ( .A(n_469), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g586 ( .A(n_469), .Y(n_586) );
OR2x2_ASAP7_75t_L g712 ( .A(n_469), .B(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_469), .B(n_478), .Y(n_716) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g491 ( .A(n_470), .Y(n_491) );
INVx1_ASAP7_75t_L g502 ( .A(n_470), .Y(n_502) );
AND2x2_ASAP7_75t_L g575 ( .A(n_470), .B(n_493), .Y(n_575) );
AND2x2_ASAP7_75t_L g615 ( .A(n_470), .B(n_494), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_475), .A2(n_542), .B(n_545), .Y(n_541) );
INVxp67_ASAP7_75t_L g657 ( .A(n_476), .Y(n_657) );
AND2x4_ASAP7_75t_L g682 ( .A(n_476), .B(n_575), .Y(n_682) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_SL g573 ( .A(n_477), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g492 ( .A(n_478), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g561 ( .A(n_478), .B(n_494), .Y(n_561) );
INVx1_ASAP7_75t_L g567 ( .A(n_478), .Y(n_567) );
INVx2_ASAP7_75t_L g593 ( .A(n_478), .Y(n_593) );
AND2x2_ASAP7_75t_L g609 ( .A(n_478), .B(n_610), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_483), .Y(n_480) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_489), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g564 ( .A(n_491), .Y(n_564) );
AND2x2_ASAP7_75t_L g672 ( .A(n_491), .B(n_493), .Y(n_672) );
AND2x2_ASAP7_75t_L g589 ( .A(n_492), .B(n_574), .Y(n_589) );
AND2x2_ASAP7_75t_L g688 ( .A(n_492), .B(n_689), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g610 ( .A(n_493), .B(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g713 ( .A(n_493), .B(n_574), .Y(n_713) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g503 ( .A(n_494), .Y(n_503) );
AND2x2_ASAP7_75t_L g592 ( .A(n_494), .B(n_593), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_497), .A2(n_525), .B(n_527), .C(n_528), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_497), .A2(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
AND2x2_ASAP7_75t_L g638 ( .A(n_501), .B(n_573), .Y(n_638) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_502), .B(n_574), .Y(n_623) );
INVx2_ASAP7_75t_L g622 ( .A(n_503), .Y(n_622) );
OAI222xp33_ASAP7_75t_L g626 ( .A1(n_503), .A2(n_566), .B1(n_627), .B2(n_629), .C1(n_630), .C2(n_633), .Y(n_626) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g551 ( .A(n_508), .Y(n_551) );
OR2x2_ASAP7_75t_L g662 ( .A(n_508), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx3_ASAP7_75t_L g584 ( .A(n_509), .Y(n_584) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_509), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g641 ( .A(n_509), .B(n_555), .Y(n_641) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g602 ( .A(n_510), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_515), .A2(n_605), .B1(n_644), .B2(n_645), .Y(n_643) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_530), .Y(n_515) );
INVx3_ASAP7_75t_L g577 ( .A(n_516), .Y(n_577) );
OR2x2_ASAP7_75t_L g710 ( .A(n_516), .B(n_586), .Y(n_710) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g583 ( .A(n_517), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g599 ( .A(n_517), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g607 ( .A(n_517), .B(n_555), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_517), .B(n_531), .Y(n_663) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g554 ( .A(n_518), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g558 ( .A(n_518), .B(n_531), .Y(n_558) );
AND2x2_ASAP7_75t_L g634 ( .A(n_518), .B(n_581), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_518), .B(n_540), .Y(n_674) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_530), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g590 ( .A(n_530), .B(n_551), .Y(n_590) );
AND2x2_ASAP7_75t_L g594 ( .A(n_530), .B(n_584), .Y(n_594) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_540), .Y(n_530) );
INVx3_ASAP7_75t_L g555 ( .A(n_531), .Y(n_555) );
AND2x2_ASAP7_75t_L g580 ( .A(n_531), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g715 ( .A(n_531), .B(n_698), .Y(n_715) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_540), .Y(n_569) );
INVx2_ASAP7_75t_L g581 ( .A(n_540), .Y(n_581) );
AND2x2_ASAP7_75t_L g625 ( .A(n_540), .B(n_601), .Y(n_625) );
INVx1_ASAP7_75t_L g668 ( .A(n_540), .Y(n_668) );
OR2x2_ASAP7_75t_L g699 ( .A(n_540), .B(n_601), .Y(n_699) );
AND2x2_ASAP7_75t_L g719 ( .A(n_540), .B(n_555), .Y(n_719) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_552), .B(n_556), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g557 ( .A(n_551), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_551), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g676 ( .A(n_553), .Y(n_676) );
INVx2_ASAP7_75t_SL g570 ( .A(n_554), .Y(n_570) );
AND2x2_ASAP7_75t_L g690 ( .A(n_554), .B(n_584), .Y(n_690) );
INVx2_ASAP7_75t_L g636 ( .A(n_555), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_555), .B(n_668), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B1(n_562), .B2(n_568), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_558), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g724 ( .A(n_558), .Y(n_724) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g649 ( .A(n_560), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_560), .B(n_592), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_561), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g665 ( .A(n_561), .B(n_614), .Y(n_665) );
INVx2_ASAP7_75t_L g721 ( .A(n_561), .Y(n_721) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g591 ( .A(n_564), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_564), .B(n_609), .Y(n_642) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_566), .B(n_586), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g703 ( .A(n_569), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_SL g653 ( .A1(n_570), .A2(n_654), .B(n_656), .C(n_659), .Y(n_653) );
OR2x2_ASAP7_75t_L g680 ( .A(n_570), .B(n_584), .Y(n_680) );
OAI221xp5_ASAP7_75t_SL g571 ( .A1(n_572), .A2(n_576), .B1(n_578), .B2(n_585), .C(n_588), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_573), .B(n_575), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_573), .B(n_622), .Y(n_629) );
AND2x2_ASAP7_75t_L g671 ( .A(n_573), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g707 ( .A(n_573), .Y(n_707) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_574), .Y(n_598) );
INVx1_ASAP7_75t_L g611 ( .A(n_574), .Y(n_611) );
NOR2xp67_ASAP7_75t_L g631 ( .A(n_577), .B(n_632), .Y(n_631) );
INVxp67_ASAP7_75t_L g685 ( .A(n_577), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_577), .B(n_625), .Y(n_701) );
INVx2_ASAP7_75t_L g687 ( .A(n_578), .Y(n_687) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g628 ( .A(n_580), .B(n_599), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_580), .A2(n_596), .B(n_638), .C(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g606 ( .A(n_581), .B(n_601), .Y(n_606) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_585), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
OR2x2_ASAP7_75t_L g654 ( .A(n_586), .B(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_591), .B2(n_594), .Y(n_588) );
INVx1_ASAP7_75t_L g708 ( .A(n_590), .Y(n_708) );
INVx1_ASAP7_75t_L g655 ( .A(n_592), .Y(n_655) );
INVx1_ASAP7_75t_L g706 ( .A(n_594), .Y(n_706) );
AOI211xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_599), .B(n_603), .C(n_626), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g618 ( .A(n_598), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g669 ( .A(n_599), .Y(n_669) );
AND2x2_ASAP7_75t_L g718 ( .A(n_599), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .B(n_616), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g632 ( .A(n_606), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_606), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g624 ( .A(n_607), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g700 ( .A(n_607), .Y(n_700) );
OAI32xp33_ASAP7_75t_L g711 ( .A1(n_607), .A2(n_659), .A3(n_666), .B1(n_707), .B2(n_712), .Y(n_711) );
NOR2xp33_ASAP7_75t_SL g608 ( .A(n_609), .B(n_612), .Y(n_608) );
INVx1_ASAP7_75t_SL g679 ( .A(n_609), .Y(n_679) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g619 ( .A(n_615), .Y(n_619) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_620), .B(n_624), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_618), .A2(n_666), .B1(n_692), .B2(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_622), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g659 ( .A(n_625), .Y(n_659) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2x1p5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g652 ( .A(n_636), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B(n_643), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_645), .A2(n_687), .B1(n_688), .B2(n_690), .C(n_691), .Y(n_686) );
NAND5xp2_ASAP7_75t_L g646 ( .A(n_647), .B(n_670), .C(n_686), .D(n_696), .E(n_714), .Y(n_646) );
AOI211xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_650), .B(n_653), .C(n_660), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g717 ( .A(n_654), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_664), .B2(n_666), .Y(n_660) );
INVx1_ASAP7_75t_SL g693 ( .A(n_663), .Y(n_693) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI322xp33_ASAP7_75t_L g675 ( .A1(n_666), .A2(n_676), .A3(n_677), .B1(n_678), .B2(n_679), .C1(n_680), .C2(n_681), .Y(n_675) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx1_ASAP7_75t_L g678 ( .A(n_668), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_668), .B(n_693), .Y(n_692) );
AOI211xp5_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_673), .B(n_675), .C(n_683), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g705 ( .A1(n_679), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_705) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g722 ( .A(n_689), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_704), .B1(n_705), .B2(n_709), .C(n_711), .Y(n_696) );
OAI211xp5_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_700), .B(n_701), .C(n_702), .Y(n_697) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g723 ( .A(n_699), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_718), .C(n_720), .Y(n_714) );
AOI21xp33_ASAP7_75t_SL g720 ( .A1(n_721), .A2(n_722), .B(n_723), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_725), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
endmodule