module fake_jpeg_1399_n_440 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_45),
.B(n_57),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_46),
.B(n_48),
.Y(n_91)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_31),
.Y(n_47)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_52),
.B(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_8),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_85),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_55),
.Y(n_100)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_63),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_7),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_64),
.B(n_69),
.Y(n_121)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_65),
.Y(n_117)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_77),
.B(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_1),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_7),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_1),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_41),
.C(n_17),
.Y(n_119)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_77),
.B1(n_72),
.B2(n_86),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_93),
.A2(n_99),
.B1(n_110),
.B2(n_111),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_18),
.B1(n_34),
.B2(n_33),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_61),
.A2(n_34),
.B1(n_16),
.B2(n_36),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_65),
.C(n_76),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_34),
.B1(n_40),
.B2(n_36),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_73),
.A2(n_34),
.B1(n_49),
.B2(n_84),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_66),
.A2(n_17),
.B1(n_40),
.B2(n_44),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_46),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_79),
.B1(n_87),
.B2(n_51),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_44),
.B1(n_23),
.B2(n_25),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_47),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_68),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_45),
.A2(n_26),
.B1(n_41),
.B2(n_37),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_91),
.B1(n_119),
.B2(n_115),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_138),
.A2(n_140),
.B1(n_159),
.B2(n_160),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_67),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_139),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_55),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_141),
.Y(n_215)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_157),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_107),
.B(n_92),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_144),
.B(n_136),
.C(n_89),
.Y(n_211)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_104),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_154),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

AO22x2_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_81),
.B1(n_75),
.B2(n_74),
.Y(n_156)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_97),
.A2(n_78),
.B(n_65),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_102),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_97),
.A2(n_58),
.B1(n_54),
.B2(n_63),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_95),
.A2(n_62),
.B1(n_60),
.B2(n_70),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_105),
.A2(n_56),
.B(n_71),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_162),
.A2(n_134),
.B(n_108),
.Y(n_212)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_100),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_165),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_50),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_167),
.B(n_169),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_80),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_172),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_112),
.B(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_11),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_112),
.A2(n_43),
.B1(n_20),
.B2(n_37),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_101),
.B(n_10),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_177),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_90),
.B1(n_103),
.B2(n_106),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_175),
.A2(n_165),
.B1(n_106),
.B2(n_109),
.Y(n_209)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_94),
.B(n_1),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_124),
.A2(n_43),
.B1(n_20),
.B2(n_37),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_178),
.A2(n_180),
.B1(n_160),
.B2(n_131),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_2),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_182),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_103),
.A2(n_37),
.B1(n_29),
.B2(n_2),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_133),
.B(n_3),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_96),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_188),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_96),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_136),
.CI(n_124),
.CON(n_193),
.SN(n_193)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_193),
.A2(n_212),
.B(n_161),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_156),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_139),
.B(n_134),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_211),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_152),
.A2(n_120),
.B1(n_109),
.B2(n_114),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_165),
.B1(n_162),
.B2(n_180),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_102),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_220),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_139),
.B(n_120),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_148),
.B(n_114),
.C(n_89),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_145),
.C(n_149),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_169),
.B1(n_138),
.B2(n_182),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_223),
.B(n_235),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_159),
.B1(n_150),
.B2(n_156),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_224),
.A2(n_233),
.B1(n_190),
.B2(n_218),
.Y(n_283)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_249),
.Y(n_274)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_227),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_156),
.B1(n_144),
.B2(n_151),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_228),
.A2(n_230),
.B1(n_256),
.B2(n_197),
.Y(n_271)
);

AOI22x1_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_156),
.B1(n_144),
.B2(n_161),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_231),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_188),
.A2(n_153),
.B1(n_167),
.B2(n_146),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_141),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_252),
.C(n_257),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_198),
.A2(n_141),
.B1(n_132),
.B2(n_181),
.Y(n_235)
);

XOR2x2_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_256),
.Y(n_267)
);

BUFx8_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_238),
.A2(n_253),
.B1(n_255),
.B2(n_192),
.Y(n_273)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_197),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_240),
.B(n_243),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_170),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_254),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_164),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_176),
.B(n_147),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_251),
.Y(n_287)
);

OAI22x1_ASAP7_75t_SL g247 ( 
.A1(n_205),
.A2(n_142),
.B1(n_155),
.B2(n_166),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_247),
.A2(n_4),
.B(n_5),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_163),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_258),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_191),
.A2(n_149),
.B1(n_171),
.B2(n_37),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_215),
.B1(n_212),
.B2(n_213),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_197),
.A2(n_171),
.B(n_29),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_191),
.B(n_171),
.C(n_29),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_198),
.A2(n_29),
.B1(n_4),
.B2(n_5),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_186),
.B(n_3),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_193),
.A2(n_214),
.B1(n_207),
.B2(n_187),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_185),
.B(n_4),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_259),
.A2(n_260),
.B1(n_280),
.B2(n_285),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_229),
.A2(n_193),
.B1(n_207),
.B2(n_220),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_184),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_194),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

XNOR2x2_ASAP7_75t_SL g266 ( 
.A(n_226),
.B(n_185),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g303 ( 
.A1(n_266),
.A2(n_232),
.B(n_251),
.C(n_252),
.D(n_247),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_236),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_202),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_272),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_211),
.C(n_221),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_275),
.C(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_271),
.B(n_228),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_195),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_273),
.A2(n_238),
.B1(n_253),
.B2(n_255),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_195),
.C(n_222),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_229),
.A2(n_210),
.B1(n_209),
.B2(n_216),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_230),
.B1(n_235),
.B2(n_250),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_199),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_277),
.B(n_284),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_213),
.C(n_216),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_242),
.A2(n_190),
.B1(n_218),
.B2(n_217),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_283),
.A2(n_286),
.B1(n_288),
.B2(n_276),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_199),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_242),
.A2(n_217),
.B1(n_192),
.B2(n_6),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_231),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_289),
.B1(n_286),
.B2(n_285),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_223),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_280),
.Y(n_344)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_297),
.A2(n_281),
.B1(n_290),
.B2(n_287),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_244),
.C(n_249),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_313),
.C(n_270),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_282),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_308),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_303),
.A2(n_322),
.B(n_262),
.C(n_266),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_232),
.Y(n_305)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_225),
.Y(n_307)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_311),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_310),
.A2(n_321),
.B(n_288),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_274),
.B(n_238),
.C(n_12),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_261),
.B(n_12),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_314),
.B(n_319),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_265),
.B(n_14),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_318),
.Y(n_346)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_14),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_304),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_290),
.A2(n_281),
.B1(n_260),
.B2(n_259),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_290),
.B(n_271),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_323),
.A2(n_342),
.B1(n_321),
.B2(n_310),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_329),
.C(n_298),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_312),
.B(n_265),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_331),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_327),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_307),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_328),
.A2(n_334),
.B1(n_343),
.B2(n_347),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_275),
.C(n_262),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_SL g331 ( 
.A(n_299),
.B(n_267),
.C(n_287),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_299),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_267),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_344),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_337),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_300),
.A2(n_266),
.B1(n_279),
.B2(n_289),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_338),
.A2(n_322),
.B1(n_295),
.B2(n_317),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_297),
.A2(n_304),
.B1(n_311),
.B2(n_315),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_302),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_318),
.Y(n_350)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_350),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_334),
.Y(n_351)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_362),
.Y(n_375)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_355),
.A2(n_357),
.B1(n_358),
.B2(n_361),
.Y(n_376)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_364),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_346),
.B(n_305),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_360),
.B(n_363),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_320),
.B1(n_303),
.B2(n_296),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_316),
.Y(n_363)
);

XNOR2x1_ASAP7_75t_SL g364 ( 
.A(n_336),
.B(n_313),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_308),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_365),
.B(n_368),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_342),
.A2(n_293),
.B1(n_294),
.B2(n_306),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_366),
.B(n_333),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_309),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_348),
.Y(n_368)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_324),
.Y(n_379)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_379),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_329),
.C(n_344),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_380),
.B(n_381),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_360),
.B(n_330),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_337),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_384),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_350),
.Y(n_383)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_351),
.B(n_348),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_338),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_333),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_349),
.C(n_364),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_388),
.B(n_391),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_376),
.A2(n_354),
.B(n_369),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_392),
.A2(n_401),
.B(n_386),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_375),
.A2(n_362),
.B(n_355),
.Y(n_394)
);

AOI21x1_ASAP7_75t_SL g402 ( 
.A1(n_394),
.A2(n_396),
.B(n_392),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_349),
.C(n_352),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_395),
.B(n_398),
.C(n_377),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_387),
.A2(n_367),
.B(n_323),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_366),
.C(n_368),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_387),
.A2(n_327),
.B(n_341),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_406),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_396),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_405),
.B(n_408),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_389),
.A2(n_377),
.B1(n_386),
.B2(n_341),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_382),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_401),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_399),
.B(n_372),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_372),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_410),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_400),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_378),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_411),
.B(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_412),
.B(n_384),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_414),
.B(n_418),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_413),
.A2(n_390),
.B(n_395),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_422),
.B(n_406),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_419),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_403),
.A2(n_388),
.B(n_393),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_374),
.C(n_357),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_423),
.B(n_358),
.Y(n_429)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_421),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_424),
.B(n_425),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_415),
.B(n_412),
.C(n_404),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_426),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_420),
.A2(n_416),
.B(n_414),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_429),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_427),
.Y(n_432)
);

AO21x1_ASAP7_75t_L g436 ( 
.A1(n_432),
.A2(n_420),
.B(n_402),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_427),
.C(n_430),
.Y(n_435)
);

OAI321xp33_ASAP7_75t_L g437 ( 
.A1(n_435),
.A2(n_436),
.A3(n_434),
.B1(n_431),
.B2(n_332),
.C(n_339),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_330),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_339),
.B(n_332),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_331),
.Y(n_440)
);


endmodule