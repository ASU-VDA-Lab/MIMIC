module fake_jpeg_21774_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_29),
.B1(n_24),
.B2(n_18),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx9p33_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_32),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_47),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_42),
.B1(n_41),
.B2(n_32),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_17),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_22),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_22),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_22),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_33),
.B1(n_52),
.B2(n_35),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_70),
.B1(n_83),
.B2(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_60),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_65),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_66),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_67),
.B(n_75),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_27),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_72),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_36),
.B1(n_22),
.B2(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_36),
.B(n_31),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_28),
.C(n_16),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_20),
.B1(n_27),
.B2(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_27),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_41),
.B1(n_42),
.B2(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_30),
.B1(n_17),
.B2(n_25),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_30),
.B1(n_25),
.B2(n_28),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_82),
.B1(n_68),
.B2(n_70),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_101),
.B1(n_53),
.B2(n_60),
.Y(n_118)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_97),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_27),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_21),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_112),
.A3(n_117),
.B1(n_96),
.B2(n_93),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_62),
.B1(n_75),
.B2(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_76),
.B1(n_85),
.B2(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_119),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_67),
.B(n_64),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_64),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_122),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_76),
.C(n_59),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_89),
.C(n_86),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_129),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_124),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_66),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_89),
.C(n_88),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_69),
.B1(n_20),
.B2(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_15),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_13),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_95),
.CI(n_98),
.CON(n_131),
.SN(n_131)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_137),
.Y(n_162)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_147),
.Y(n_153)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_145),
.B1(n_112),
.B2(n_138),
.C(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_86),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_121),
.C(n_116),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_146),
.B(n_10),
.Y(n_160)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_88),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_129),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_155),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_157),
.C(n_143),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_156),
.A2(n_163),
.B1(n_134),
.B2(n_149),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_111),
.Y(n_157)
);

OAI322xp33_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_126),
.A3(n_112),
.B1(n_117),
.B2(n_124),
.C1(n_130),
.C2(n_128),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_146),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_140),
.B(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_130),
.B1(n_74),
.B2(n_90),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_143),
.B1(n_133),
.B2(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_168),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_167),
.B(n_171),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_144),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_172),
.C(n_152),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_90),
.B(n_9),
.Y(n_182)
);

OAI322xp33_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_157),
.A3(n_154),
.B1(n_164),
.B2(n_163),
.C1(n_156),
.C2(n_150),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_177),
.C(n_184),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_162),
.C(n_154),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_182),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_171),
.A2(n_53),
.B1(n_1),
.B2(n_2),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_0),
.C(n_1),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_174),
.B(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_180),
.A2(n_175),
.B(n_1),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_189),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_179),
.C2(n_187),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_195),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_188),
.Y(n_198)
);

AOI221xp5_ASAP7_75t_L g201 ( 
.A1(n_198),
.A2(n_199),
.B1(n_6),
.B2(n_7),
.C(n_194),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_191),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_194),
.B1(n_188),
.B2(n_8),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_6),
.Y(n_204)
);


endmodule