module real_jpeg_9578_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_321, n_11, n_14, n_7, n_322, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_321;
input n_11;
input n_14;
input n_7;
input n_322;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_1),
.A2(n_48),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_1),
.B(n_48),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_1),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_1),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_1),
.A2(n_34),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_34),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_38),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_1),
.A2(n_31),
.B(n_35),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_1),
.A2(n_25),
.B1(n_27),
.B2(n_110),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_2),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_97),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_97),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_2),
.A2(n_25),
.B1(n_27),
.B2(n_97),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_25),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_4),
.A2(n_37),
.B1(n_48),
.B2(n_49),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_4),
.A2(n_37),
.B1(n_63),
.B2(n_64),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_5),
.A2(n_25),
.B1(n_27),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_5),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_58),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_6),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_7),
.A2(n_25),
.B1(n_27),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_7),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_56),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_56),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_48),
.B(n_61),
.C(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_8),
.B(n_48),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_9),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_10),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_10),
.A2(n_24),
.B1(n_63),
.B2(n_64),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_10),
.A2(n_24),
.B1(n_48),
.B2(n_49),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_13),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_85),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_85),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_13),
.A2(n_25),
.B1(n_27),
.B2(n_85),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_14),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_144),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_14),
.A2(n_34),
.B1(n_35),
.B2(n_144),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_14),
.A2(n_25),
.B1(n_27),
.B2(n_144),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_16),
.A2(n_63),
.B1(n_64),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_16),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_16),
.A2(n_48),
.B1(n_49),
.B2(n_90),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_16),
.A2(n_34),
.B1(n_35),
.B2(n_90),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_16),
.A2(n_25),
.B1(n_27),
.B2(n_90),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_17),
.A2(n_63),
.B1(n_64),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_17),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_17),
.A2(n_48),
.B1(n_49),
.B2(n_126),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_17),
.A2(n_34),
.B1(n_35),
.B2(n_126),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_17),
.A2(n_25),
.B1(n_27),
.B2(n_126),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_72),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_71),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_39),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_36),
.B2(n_38),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_23),
.A2(n_28),
.B1(n_38),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_25),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_30),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_25),
.A2(n_30),
.B(n_110),
.C(n_174),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_28),
.A2(n_38),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_29),
.A2(n_33),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_29),
.A2(n_33),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_29),
.A2(n_33),
.B1(n_207),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_29),
.A2(n_33),
.B1(n_232),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_29),
.A2(n_33),
.B1(n_250),
.B2(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_29),
.A2(n_33),
.B1(n_55),
.B2(n_271),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_45),
.Y(n_46)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_67),
.C(n_69),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_40),
.A2(n_41),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_53),
.C(n_59),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_42),
.A2(n_43),
.B1(n_59),
.B2(n_297),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_43)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_47),
.B(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_44),
.A2(n_47),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_44),
.A2(n_47),
.B1(n_135),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_44),
.A2(n_47),
.B1(n_152),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_44),
.A2(n_47),
.B1(n_192),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_44),
.A2(n_47),
.B1(n_203),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_44),
.A2(n_47),
.B1(n_229),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_44),
.A2(n_47),
.B1(n_247),
.B2(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_44),
.A2(n_47),
.B1(n_51),
.B2(n_264),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_46),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_47),
.B(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_48),
.B(n_50),
.Y(n_139)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_49),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_53),
.A2(n_54),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_59),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_59),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_66),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_62),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_60),
.A2(n_62),
.B1(n_96),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_60),
.A2(n_62),
.B1(n_123),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_60),
.A2(n_62),
.B1(n_131),
.B2(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_60),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_60),
.A2(n_62),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_60),
.A2(n_62),
.B1(n_215),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_60),
.A2(n_62),
.B1(n_224),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_60),
.A2(n_62),
.B1(n_66),
.B2(n_256),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_62),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_62),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_65),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_63),
.B(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_67),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_312),
.B(n_318),
.Y(n_72)
);

OAI321xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_289),
.A3(n_307),
.B1(n_310),
.B2(n_311),
.C(n_321),
.Y(n_73)
);

AOI321xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_240),
.A3(n_277),
.B1(n_283),
.B2(n_288),
.C(n_322),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_197),
.C(n_236),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_167),
.B(n_196),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_146),
.B(n_166),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_128),
.B(n_145),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_117),
.B(n_127),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_103),
.B(n_116),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_91),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_91),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_86),
.A2(n_87),
.B1(n_143),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_107),
.B1(n_108),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_102),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_102),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_111),
.B(n_115),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_109),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_108),
.B1(n_125),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_107),
.A2(n_108),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_107),
.A2(n_108),
.B1(n_178),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_107),
.A2(n_108),
.B1(n_212),
.B2(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_107),
.A2(n_108),
.B(n_222),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_129),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.CI(n_124),
.CON(n_120),
.SN(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.CI(n_136),
.CON(n_129),
.SN(n_129)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_148),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_159),
.B2(n_160),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_162),
.C(n_164),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_158),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_156),
.C(n_158),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_161),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_162),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_169),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_182),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_171),
.B(n_181),
.C(n_182),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_176),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_179),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_190),
.B2(n_191),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_190),
.C(n_193),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_198),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_217),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_199),
.B(n_217),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_210),
.C(n_216),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_209),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_208),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_208),
.C(n_209),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_216),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_213),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_234),
.B2(n_235),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_220),
.B(n_225),
.C(n_235),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_223),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_230),
.C(n_233),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_228),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_238),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_259),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_241),
.B(n_259),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_252),
.C(n_258),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_242),
.A2(n_243),
.B1(n_252),
.B2(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_248),
.C(n_251),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_248),
.B1(n_249),
.B2(n_251),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_246),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_252),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_254),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_253),
.A2(n_270),
.B(n_273),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_255),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_255),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_275),
.B2(n_276),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_267),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_267),
.C(n_276),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_265),
.B(n_266),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_265),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_291),
.C(n_299),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_266),
.B(n_291),
.CI(n_299),
.CON(n_309),
.SN(n_309)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_273),
.B2(n_274),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_270),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_275),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_284),
.B(n_287),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_279),
.B(n_280),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_300),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_300),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_292),
.A2(n_293),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_297),
.C(n_298),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_302),
.C(n_306),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_296),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_308),
.B(n_309),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_309),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_317),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_317),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_314),
.Y(n_316)
);


endmodule