module fake_jpeg_16933_n_40 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_40);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

INVx8_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_2),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_1),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_17),
.A2(n_5),
.B1(n_18),
.B2(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_16),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.Y(n_33)
);

AO22x1_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_22),
.B1(n_13),
.B2(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_19),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_21),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_23),
.B(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

MAJx2_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_28),
.C(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_36),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_31),
.B(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_15),
.B1(n_32),
.B2(n_35),
.Y(n_40)
);


endmodule