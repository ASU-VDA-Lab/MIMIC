module fake_jpeg_31960_n_193 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_193);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_18),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_56),
.Y(n_71)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_25),
.B1(n_28),
.B2(n_23),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_40),
.B1(n_27),
.B2(n_26),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_56),
.C(n_42),
.Y(n_58)
);

XNOR2x1_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_17),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_34),
.B(n_37),
.C(n_33),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_59),
.B(n_61),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_36),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_37),
.B(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_74),
.Y(n_91)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_75),
.B1(n_35),
.B2(n_26),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_35),
.B1(n_32),
.B2(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_60),
.Y(n_107)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_22),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_20),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_35),
.B(n_17),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_99),
.B(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_101),
.B1(n_32),
.B2(n_80),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_28),
.B1(n_25),
.B2(n_35),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_75),
.B1(n_71),
.B2(n_69),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_59),
.A2(n_27),
.B1(n_28),
.B2(n_23),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_17),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_58),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_110),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_117),
.B1(n_124),
.B2(n_15),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_113),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_65),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_118),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_104),
.B1(n_96),
.B2(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_20),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_125),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_66),
.B(n_85),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_122),
.A2(n_97),
.B1(n_90),
.B2(n_106),
.Y(n_128)
);

XOR2x2_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_29),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_67),
.B1(n_72),
.B2(n_17),
.Y(n_124)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_32),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_62),
.C(n_79),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_62),
.C(n_87),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_15),
.B1(n_30),
.B2(n_16),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_100),
.B(n_93),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_132),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_93),
.B(n_87),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_135),
.C(n_143),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_83),
.C(n_67),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_138),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_112),
.Y(n_138)
);

AO221x1_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_114),
.B1(n_120),
.B2(n_125),
.C(n_126),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_39),
.C(n_15),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_144),
.A2(n_109),
.B(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_122),
.B(n_116),
.Y(n_147)
);

HAxp5_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_29),
.CON(n_162),
.SN(n_162)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_127),
.C(n_115),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_133),
.C(n_136),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_21),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_39),
.B(n_29),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_157),
.B(n_21),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_136),
.B1(n_143),
.B2(n_30),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_144),
.C(n_140),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_162),
.B1(n_166),
.B2(n_155),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_39),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_39),
.C(n_16),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_145),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_171),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_156),
.B1(n_147),
.B2(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_173),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_150),
.C(n_154),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_175),
.C(n_164),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_157),
.B1(n_9),
.B2(n_10),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_162),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_8),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_21),
.C(n_6),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_163),
.B(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_178),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_169),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_14),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_11),
.Y(n_183)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_169),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_183),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_184),
.B(n_180),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_187),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_188),
.B(n_185),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_189),
.C(n_4),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_3),
.Y(n_193)
);


endmodule