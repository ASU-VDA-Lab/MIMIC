module fake_jpeg_692_n_70 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_70);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_70;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_67;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_6),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_28),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_2),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_27),
.Y(n_37)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_25),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_21),
.A2(n_14),
.B1(n_16),
.B2(n_13),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_14),
.B1(n_16),
.B2(n_9),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_6),
.B1(n_10),
.B2(n_23),
.Y(n_34)
);

NOR2xp67_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_46),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_47),
.B(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_38),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_36),
.C(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_62),
.B(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_65),
.Y(n_68)
);

AOI21x1_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_40),
.B(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_69),
.B(n_56),
.Y(n_70)
);


endmodule