module real_aes_2670_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_0), .B(n_502), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_1), .A2(n_504), .B(n_505), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_2), .B(n_796), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_3), .A2(n_4), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_3), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_4), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_5), .B(n_220), .Y(n_539) );
INVx1_ASAP7_75t_L g152 ( .A(n_6), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_7), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_8), .B(n_220), .Y(n_588) );
INVx1_ASAP7_75t_L g190 ( .A(n_9), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g796 ( .A(n_10), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_11), .Y(n_158) );
NAND2xp33_ASAP7_75t_L g580 ( .A(n_12), .B(n_217), .Y(n_580) );
INVx2_ASAP7_75t_L g134 ( .A(n_13), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g113 ( .A1(n_14), .A2(n_114), .B1(n_115), .B2(n_118), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_14), .Y(n_118) );
AOI221x1_ASAP7_75t_L g524 ( .A1(n_15), .A2(n_29), .B1(n_502), .B2(n_504), .C(n_525), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_16), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_17), .B(n_502), .Y(n_576) );
AOI22xp5_ASAP7_75t_SL g111 ( .A1(n_18), .A2(n_112), .B1(n_113), .B2(n_119), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_18), .Y(n_119) );
INVx1_ASAP7_75t_L g218 ( .A(n_19), .Y(n_218) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_20), .A2(n_187), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_21), .B(n_182), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_22), .A2(n_82), .B1(n_818), .B2(n_819), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_22), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_23), .B(n_220), .Y(n_513) );
AO21x1_ASAP7_75t_L g534 ( .A1(n_24), .A2(n_502), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g108 ( .A(n_25), .Y(n_108) );
INVx1_ASAP7_75t_L g215 ( .A(n_26), .Y(n_215) );
INVx1_ASAP7_75t_SL g202 ( .A(n_27), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_28), .B(n_145), .Y(n_260) );
AOI33xp33_ASAP7_75t_L g240 ( .A1(n_30), .A2(n_55), .A3(n_138), .B1(n_163), .B2(n_241), .B3(n_242), .Y(n_240) );
NAND2x1_ASAP7_75t_L g555 ( .A(n_31), .B(n_220), .Y(n_555) );
NAND2x1_ASAP7_75t_L g587 ( .A(n_32), .B(n_217), .Y(n_587) );
INVx1_ASAP7_75t_L g143 ( .A(n_33), .Y(n_143) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_34), .A2(n_89), .B(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g184 ( .A(n_34), .B(n_89), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_35), .B(n_167), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_36), .B(n_217), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_37), .B(n_220), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_38), .B(n_217), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_39), .A2(n_504), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g151 ( .A(n_40), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g162 ( .A(n_40), .Y(n_162) );
AND2x2_ASAP7_75t_L g171 ( .A(n_40), .B(n_141), .Y(n_171) );
OR2x6_ASAP7_75t_L g106 ( .A(n_41), .B(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_42), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_43), .B(n_502), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_44), .B(n_167), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_45), .A2(n_132), .B1(n_209), .B2(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_46), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_47), .B(n_145), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_48), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_49), .B(n_217), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_50), .B(n_187), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_51), .B(n_145), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_52), .A2(n_504), .B(n_586), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_53), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_54), .B(n_217), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_56), .B(n_145), .Y(n_179) );
INVx1_ASAP7_75t_L g139 ( .A(n_57), .Y(n_139) );
INVx1_ASAP7_75t_L g147 ( .A(n_57), .Y(n_147) );
AND2x2_ASAP7_75t_L g181 ( .A(n_58), .B(n_182), .Y(n_181) );
AOI221xp5_ASAP7_75t_L g188 ( .A1(n_59), .A2(n_77), .B1(n_160), .B2(n_167), .C(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_60), .B(n_167), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_61), .B(n_220), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_62), .B(n_132), .Y(n_165) );
AOI21xp5_ASAP7_75t_SL g227 ( .A1(n_63), .A2(n_160), .B(n_228), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_64), .A2(n_504), .B(n_554), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_65), .Y(n_786) );
INVx1_ASAP7_75t_L g212 ( .A(n_66), .Y(n_212) );
AO21x1_ASAP7_75t_L g536 ( .A1(n_67), .A2(n_504), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_68), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g178 ( .A(n_69), .Y(n_178) );
XOR2xp5_ASAP7_75t_L g814 ( .A(n_70), .B(n_85), .Y(n_814) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_71), .B(n_502), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_72), .A2(n_160), .B(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g549 ( .A(n_73), .B(n_183), .Y(n_549) );
INVx1_ASAP7_75t_L g141 ( .A(n_74), .Y(n_141) );
INVx1_ASAP7_75t_L g149 ( .A(n_74), .Y(n_149) );
AND2x2_ASAP7_75t_L g590 ( .A(n_75), .B(n_131), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_76), .B(n_167), .Y(n_243) );
AND2x2_ASAP7_75t_L g204 ( .A(n_78), .B(n_131), .Y(n_204) );
INVx1_ASAP7_75t_L g213 ( .A(n_79), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_80), .A2(n_160), .B(n_201), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_81), .A2(n_160), .B(n_235), .C(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g819 ( .A(n_82), .Y(n_819) );
INVx1_ASAP7_75t_L g109 ( .A(n_83), .Y(n_109) );
AND2x2_ASAP7_75t_L g499 ( .A(n_84), .B(n_131), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_85), .A2(n_104), .B1(n_789), .B2(n_800), .C(n_809), .Y(n_103) );
AND2x2_ASAP7_75t_SL g225 ( .A(n_85), .B(n_131), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_86), .B(n_502), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_87), .A2(n_160), .B1(n_238), .B2(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g535 ( .A(n_88), .B(n_209), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_90), .B(n_217), .Y(n_514) );
AND2x2_ASAP7_75t_L g558 ( .A(n_91), .B(n_131), .Y(n_558) );
INVx1_ASAP7_75t_L g229 ( .A(n_92), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_93), .B(n_220), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_94), .A2(n_504), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_95), .B(n_217), .Y(n_526) );
AND2x2_ASAP7_75t_L g244 ( .A(n_96), .B(n_131), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_97), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_98), .B(n_220), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_99), .A2(n_136), .B(n_142), .C(n_150), .Y(n_135) );
BUFx2_ASAP7_75t_L g797 ( .A(n_100), .Y(n_797) );
BUFx2_ASAP7_75t_SL g806 ( .A(n_100), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_101), .A2(n_504), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_102), .B(n_145), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_110), .B1(n_786), .B2(n_787), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_105), .B(n_491), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g788 ( .A(n_106), .B(n_491), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
XOR2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_120), .Y(n_110) );
INVxp33_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_489), .B1(n_490), .B2(n_492), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_368), .C(n_435), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_328), .Y(n_123) );
NOR3x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_279), .C(n_308), .Y(n_124) );
OAI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_193), .B1(n_232), .B2(n_247), .C(n_264), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_SL g442 ( .A1(n_126), .A2(n_206), .B(n_443), .C(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_127), .A2(n_414), .B1(n_417), .B2(n_419), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_127), .B(n_233), .Y(n_488) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_172), .Y(n_127) );
BUFx2_ASAP7_75t_L g407 ( .A(n_128), .Y(n_407) );
INVx1_ASAP7_75t_SL g420 ( .A(n_128), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_128), .B(n_275), .Y(n_462) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g245 ( .A(n_129), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g290 ( .A(n_129), .B(n_186), .Y(n_290) );
INVx1_ASAP7_75t_L g301 ( .A(n_129), .Y(n_301) );
INVx2_ASAP7_75t_L g305 ( .A(n_129), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_129), .B(n_276), .Y(n_432) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_155), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B1(n_153), .B2(n_154), .Y(n_130) );
INVx3_ASAP7_75t_L g154 ( .A(n_131), .Y(n_154) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_132), .B(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_133), .Y(n_187) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_134), .B(n_184), .Y(n_183) );
AND2x4_ASAP7_75t_L g209 ( .A(n_134), .B(n_184), .Y(n_209) );
INVxp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_137), .A2(n_178), .B(n_179), .C(n_180), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g189 ( .A1(n_137), .A2(n_180), .B(n_190), .C(n_191), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_SL g201 ( .A1(n_137), .A2(n_180), .B(n_202), .C(n_203), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_137), .A2(n_144), .B1(n_212), .B2(n_213), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_137), .A2(n_180), .B(n_229), .C(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g262 ( .A(n_137), .Y(n_262) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
AND2x2_ASAP7_75t_L g168 ( .A(n_138), .B(n_169), .Y(n_168) );
INVxp33_ASAP7_75t_L g241 ( .A(n_138), .Y(n_241) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g164 ( .A(n_139), .B(n_152), .Y(n_164) );
AND2x4_ASAP7_75t_L g220 ( .A(n_139), .B(n_148), .Y(n_220) );
INVx3_ASAP7_75t_L g163 ( .A(n_140), .Y(n_163) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x6_ASAP7_75t_L g217 ( .A(n_141), .B(n_146), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g502 ( .A(n_145), .B(n_151), .Y(n_502) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx5_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_154), .A2(n_174), .B(n_181), .Y(n_173) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_154), .A2(n_174), .B(n_181), .Y(n_276) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_154), .A2(n_543), .B(n_549), .Y(n_542) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_154), .A2(n_552), .B(n_558), .Y(n_551) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_154), .A2(n_552), .B(n_558), .Y(n_564) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_154), .A2(n_543), .B(n_549), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .B1(n_165), .B2(n_166), .Y(n_155) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVxp67_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_164), .Y(n_160) );
NOR2x1p5_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVx1_ASAP7_75t_L g242 ( .A(n_163), .Y(n_242) );
AND2x6_ASAP7_75t_L g504 ( .A(n_164), .B(n_171), .Y(n_504) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_170), .Y(n_167) );
INVx1_ASAP7_75t_L g255 ( .A(n_168), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_170), .Y(n_256) );
BUFx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g381 ( .A(n_172), .B(n_382), .Y(n_381) );
NOR2x1_ASAP7_75t_L g172 ( .A(n_173), .B(n_185), .Y(n_172) );
INVx2_ASAP7_75t_L g284 ( .A(n_173), .Y(n_284) );
AND2x2_ASAP7_75t_L g304 ( .A(n_173), .B(n_305), .Y(n_304) );
NOR2xp67_ASAP7_75t_L g429 ( .A(n_173), .B(n_305), .Y(n_429) );
AND2x2_ASAP7_75t_L g454 ( .A(n_173), .B(n_297), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_180), .B(n_209), .Y(n_221) );
INVx1_ASAP7_75t_L g238 ( .A(n_180), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_180), .A2(n_260), .B(n_261), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_180), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_180), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_180), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_180), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_180), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_180), .A2(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_180), .A2(n_579), .B(n_580), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_180), .A2(n_587), .B(n_588), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_182), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_182), .A2(n_501), .B(n_503), .Y(n_500) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_182), .A2(n_524), .B(n_528), .Y(n_523) );
OA21x2_ASAP7_75t_L g594 ( .A1(n_182), .A2(n_524), .B(n_528), .Y(n_594) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g246 ( .A(n_186), .Y(n_246) );
INVx1_ASAP7_75t_L g268 ( .A(n_186), .Y(n_268) );
INVxp67_ASAP7_75t_L g307 ( .A(n_186), .Y(n_307) );
AND2x4_ASAP7_75t_L g347 ( .A(n_186), .B(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_186), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_186), .B(n_298), .Y(n_433) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_192), .Y(n_186) );
INVx2_ASAP7_75t_SL g235 ( .A(n_187), .Y(n_235) );
INVx1_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_205), .Y(n_194) );
AND2x2_ASAP7_75t_L g321 ( .A(n_195), .B(n_293), .Y(n_321) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_196), .Y(n_249) );
AND2x2_ASAP7_75t_L g277 ( .A(n_196), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g288 ( .A(n_196), .Y(n_288) );
INVx1_ASAP7_75t_L g312 ( .A(n_196), .Y(n_312) );
AND2x2_ASAP7_75t_L g315 ( .A(n_196), .B(n_207), .Y(n_315) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_196), .Y(n_337) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_204), .Y(n_196) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_197), .A2(n_584), .B(n_590), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
NOR2x1_ASAP7_75t_L g205 ( .A(n_206), .B(n_222), .Y(n_205) );
AND2x2_ASAP7_75t_L g302 ( .A(n_206), .B(n_224), .Y(n_302) );
NAND2x1_ASAP7_75t_L g335 ( .A(n_206), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g438 ( .A(n_206), .Y(n_438) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g278 ( .A(n_207), .Y(n_278) );
AND2x2_ASAP7_75t_L g293 ( .A(n_207), .B(n_252), .Y(n_293) );
NOR2x1_ASAP7_75t_SL g362 ( .A(n_207), .B(n_224), .Y(n_362) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_210), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_209), .A2(n_227), .B(n_231), .Y(n_226) );
INVx1_ASAP7_75t_SL g509 ( .A(n_209), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_209), .B(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_209), .A2(n_576), .B(n_577), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_214), .B(n_221), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B1(n_218), .B2(n_219), .Y(n_214) );
INVxp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVxp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_222), .B(n_386), .Y(n_399) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g324 ( .A(n_223), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx4_ASAP7_75t_L g263 ( .A(n_224), .Y(n_263) );
AND2x4_ASAP7_75t_L g270 ( .A(n_224), .B(n_271), .Y(n_270) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_224), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_224), .B(n_287), .Y(n_387) );
AND2x2_ASAP7_75t_L g415 ( .A(n_224), .B(n_252), .Y(n_415) );
OR2x6_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
NAND2x1_ASAP7_75t_SL g232 ( .A(n_233), .B(n_245), .Y(n_232) );
OR2x2_ASAP7_75t_L g443 ( .A(n_233), .B(n_355), .Y(n_443) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x4_ASAP7_75t_L g283 ( .A(n_234), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g348 ( .A(n_234), .Y(n_348) );
AND2x2_ASAP7_75t_L g382 ( .A(n_234), .B(n_305), .Y(n_382) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_244), .Y(n_234) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_235), .A2(n_236), .B(n_244), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_237), .B(n_243), .Y(n_236) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g355 ( .A(n_245), .Y(n_355) );
AND2x2_ASAP7_75t_L g363 ( .A(n_245), .B(n_296), .Y(n_363) );
AND2x2_ASAP7_75t_L g480 ( .A(n_245), .B(n_283), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g434 ( .A(n_249), .B(n_375), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_249), .B(n_274), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_250), .A2(n_311), .B(n_314), .Y(n_310) );
AND2x2_ASAP7_75t_L g380 ( .A(n_250), .B(n_286), .Y(n_380) );
INVx2_ASAP7_75t_SL g467 ( .A(n_250), .Y(n_467) );
AND2x4_ASAP7_75t_SL g250 ( .A(n_251), .B(n_263), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g271 ( .A(n_252), .Y(n_271) );
INVx2_ASAP7_75t_L g318 ( .A(n_252), .Y(n_318) );
AND2x4_ASAP7_75t_L g325 ( .A(n_252), .B(n_278), .Y(n_325) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_258), .Y(n_252) );
NOR3xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .C(n_257), .Y(n_254) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_263), .Y(n_281) );
AND2x4_ASAP7_75t_L g357 ( .A(n_263), .B(n_271), .Y(n_357) );
OR2x2_ASAP7_75t_L g483 ( .A(n_263), .B(n_484), .Y(n_483) );
NAND4xp25_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .C(n_272), .D(n_277), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g330 ( .A(n_266), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g427 ( .A(n_266), .Y(n_427) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_267), .B(n_275), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_267), .B(n_332), .Y(n_461) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_270), .B(n_286), .Y(n_339) );
INVx2_ASAP7_75t_L g441 ( .A(n_270), .Y(n_441) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_270), .B(n_311), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_270), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g343 ( .A(n_274), .B(n_290), .Y(n_343) );
AND2x2_ASAP7_75t_L g411 ( .A(n_274), .B(n_347), .Y(n_411) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g296 ( .A(n_275), .B(n_297), .Y(n_296) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_276), .Y(n_350) );
AND2x2_ASAP7_75t_L g401 ( .A(n_276), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_276), .B(n_298), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_277), .B(n_441), .Y(n_448) );
INVx1_ASAP7_75t_SL g484 ( .A(n_277), .Y(n_484) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
AND2x2_ASAP7_75t_L g375 ( .A(n_278), .B(n_318), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_289), .B(n_291), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
AND2x2_ASAP7_75t_L g341 ( .A(n_283), .B(n_290), .Y(n_341) );
AND2x2_ASAP7_75t_L g449 ( .A(n_283), .B(n_300), .Y(n_449) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g323 ( .A(n_286), .Y(n_323) );
AND2x2_ASAP7_75t_L g356 ( .A(n_286), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g361 ( .A(n_286), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_286), .B(n_325), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_286), .B(n_461), .C(n_462), .Y(n_460) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B1(n_302), .B2(n_303), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g386 ( .A(n_293), .Y(n_386) );
AND2x2_ASAP7_75t_L g320 ( .A(n_294), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g342 ( .A(n_294), .B(n_315), .Y(n_342) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_294), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
INVx1_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
AND2x2_ASAP7_75t_L g306 ( .A(n_297), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g395 ( .A(n_301), .B(n_347), .Y(n_395) );
INVx1_ASAP7_75t_L g453 ( .A(n_301), .Y(n_453) );
INVx1_ASAP7_75t_L g309 ( .A(n_303), .Y(n_309) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_304), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g440 ( .A(n_304), .B(n_347), .Y(n_440) );
AND2x2_ASAP7_75t_L g406 ( .A(n_306), .B(n_407), .Y(n_406) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_306), .B(n_475), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B(n_319), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_311), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g367 ( .A(n_311), .B(n_316), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_311), .B(n_357), .Y(n_418) );
AND2x4_ASAP7_75t_SL g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_312), .B(n_375), .Y(n_405) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_312), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_314), .A2(n_341), .B1(n_342), .B2(n_343), .Y(n_340) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_315), .B(n_357), .Y(n_376) );
INVx1_ASAP7_75t_L g477 ( .A(n_315), .Y(n_477) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_322), .B(n_326), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_321), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g458 ( .A(n_324), .Y(n_458) );
INVx4_ASAP7_75t_L g360 ( .A(n_325), .Y(n_360) );
INVxp33_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g388 ( .A(n_327), .B(n_389), .Y(n_388) );
NOR2x1_ASAP7_75t_L g328 ( .A(n_329), .B(n_344), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B(n_340), .Y(n_329) );
INVx1_ASAP7_75t_L g378 ( .A(n_331), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_338), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g383 ( .A(n_335), .Y(n_383) );
INVx1_ASAP7_75t_L g416 ( .A(n_336), .Y(n_416) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_341), .A2(n_380), .B1(n_381), .B2(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g393 ( .A(n_342), .Y(n_393) );
NAND4xp25_ASAP7_75t_SL g344 ( .A(n_345), .B(n_351), .C(n_358), .D(n_364), .Y(n_344) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g366 ( .A(n_347), .Y(n_366) );
AND2x2_ASAP7_75t_L g478 ( .A(n_347), .B(n_475), .Y(n_478) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_356), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g485 ( .A(n_355), .B(n_422), .Y(n_485) );
INVx1_ASAP7_75t_L g482 ( .A(n_356), .Y(n_482) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_357), .Y(n_391) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_363), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_396), .Y(n_368) );
NOR3xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_384), .C(n_392), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_377), .B(n_379), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_374), .A2(n_406), .B1(n_409), .B2(n_411), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_377), .A2(n_385), .B1(n_388), .B2(n_390), .Y(n_384) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g389 ( .A(n_382), .Y(n_389) );
AND2x4_ASAP7_75t_L g400 ( .A(n_382), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_387), .Y(n_487) );
AOI31xp33_ASAP7_75t_L g486 ( .A1(n_390), .A2(n_463), .A3(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_412), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_398), .B(n_408), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_403), .B2(n_406), .Y(n_398) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_402), .Y(n_466) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_410), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_413), .B(n_423), .Y(n_412) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
AND2x2_ASAP7_75t_L g424 ( .A(n_415), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g463 ( .A(n_415), .Y(n_463) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_415), .A2(n_473), .B1(n_476), .B2(n_478), .Y(n_472) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_420), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_430), .B2(n_434), .Y(n_423) );
NOR2xp33_ASAP7_75t_SL g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx2_ASAP7_75t_SL g475 ( .A(n_432), .Y(n_475) );
INVx2_ASAP7_75t_L g456 ( .A(n_433), .Y(n_456) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_470), .Y(n_435) );
AOI211xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_442), .B(n_445), .C(n_459), .Y(n_436) );
OAI21xp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_441), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_446), .B(n_450), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B1(n_455), .B2(n_457), .Y(n_450) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AND2x2_ASAP7_75t_L g455 ( .A(n_453), .B(n_456), .Y(n_455) );
AO22x1_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B1(n_464), .B2(n_468), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_481), .C(n_486), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_472), .B(n_479), .Y(n_471) );
INVx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI21xp33_ASAP7_75t_R g481 ( .A1(n_482), .A2(n_483), .B(n_485), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_SL g816 ( .A(n_492), .Y(n_816) );
NOR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_673), .Y(n_492) );
AO211x2_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_518), .B(n_568), .C(n_641), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
AND3x2_ASAP7_75t_L g722 ( .A(n_496), .B(n_603), .C(n_619), .Y(n_722) );
AND2x4_ASAP7_75t_L g725 ( .A(n_496), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_508), .Y(n_496) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_497), .B(n_582), .Y(n_581) );
INVx4_ASAP7_75t_L g634 ( .A(n_497), .Y(n_634) );
AND2x2_ASAP7_75t_SL g719 ( .A(n_497), .B(n_628), .Y(n_719) );
AND2x2_ASAP7_75t_L g762 ( .A(n_497), .B(n_583), .Y(n_762) );
INVx5_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g611 ( .A(n_498), .Y(n_611) );
AND2x2_ASAP7_75t_L g630 ( .A(n_498), .B(n_574), .Y(n_630) );
AND2x2_ASAP7_75t_L g648 ( .A(n_498), .B(n_583), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_498), .B(n_582), .Y(n_708) );
NOR2x1_ASAP7_75t_SL g735 ( .A(n_498), .B(n_508), .Y(n_735) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_508), .B(n_574), .Y(n_573) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_516), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_509), .B(n_517), .Y(n_516) );
AO21x2_ASAP7_75t_L g607 ( .A1(n_509), .A2(n_510), .B(n_516), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
AO21x1_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_550), .B(n_559), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_520), .A2(n_617), .B1(n_621), .B2(n_622), .Y(n_616) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_529), .Y(n_520) );
AND2x2_ASAP7_75t_L g677 ( .A(n_521), .B(n_565), .Y(n_677) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g610 ( .A(n_522), .B(n_593), .Y(n_610) );
AND2x2_ASAP7_75t_L g682 ( .A(n_522), .B(n_567), .Y(n_682) );
AND2x2_ASAP7_75t_L g701 ( .A(n_522), .B(n_667), .Y(n_701) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g560 ( .A(n_523), .Y(n_560) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_523), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_529), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g661 ( .A(n_530), .B(n_562), .Y(n_661) );
AND2x4_ASAP7_75t_L g530 ( .A(n_531), .B(n_542), .Y(n_530) );
AND2x2_ASAP7_75t_L g565 ( .A(n_531), .B(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g598 ( .A(n_531), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_SL g658 ( .A(n_531), .B(n_594), .Y(n_658) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g751 ( .A(n_532), .Y(n_751) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g593 ( .A(n_533), .Y(n_593) );
OAI21x1_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_536), .B(n_540), .Y(n_533) );
INVx1_ASAP7_75t_L g541 ( .A(n_535), .Y(n_541) );
INVx2_ASAP7_75t_L g599 ( .A(n_542), .Y(n_599) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_542), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_548), .Y(n_543) );
INVx2_ASAP7_75t_L g595 ( .A(n_550), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_550), .B(n_727), .Y(n_753) );
AND2x2_ASAP7_75t_L g772 ( .A(n_550), .B(n_762), .Y(n_772) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_SL g640 ( .A(n_551), .B(n_599), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
AND2x2_ASAP7_75t_SL g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g639 ( .A(n_560), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_560), .B(n_609), .Y(n_644) );
INVx1_ASAP7_75t_SL g771 ( .A(n_560), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_561), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
INVx1_ASAP7_75t_L g597 ( .A(n_562), .Y(n_597) );
AND2x2_ASAP7_75t_L g783 ( .A(n_562), .B(n_784), .Y(n_783) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g659 ( .A(n_563), .B(n_566), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_563), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g713 ( .A(n_563), .B(n_567), .Y(n_713) );
AND2x2_ASAP7_75t_L g744 ( .A(n_563), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g609 ( .A(n_564), .B(n_567), .Y(n_609) );
INVxp67_ASAP7_75t_L g626 ( .A(n_564), .Y(n_626) );
BUFx3_ASAP7_75t_L g667 ( .A(n_564), .Y(n_667) );
AND2x2_ASAP7_75t_L g687 ( .A(n_565), .B(n_688), .Y(n_687) );
NAND2xp33_ASAP7_75t_L g700 ( .A(n_565), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_566), .B(n_593), .Y(n_656) );
AND2x2_ASAP7_75t_L g745 ( .A(n_566), .B(n_594), .Y(n_745) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g672 ( .A(n_567), .B(n_594), .Y(n_672) );
OR3x1_ASAP7_75t_L g568 ( .A(n_569), .B(n_616), .C(n_631), .Y(n_568) );
OAI321xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_581), .A3(n_591), .B1(n_596), .B2(n_600), .C(n_608), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_573), .Y(n_647) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_573), .Y(n_665) );
OR2x2_ASAP7_75t_L g669 ( .A(n_573), .B(n_581), .Y(n_669) );
BUFx3_ASAP7_75t_L g603 ( .A(n_574), .Y(n_603) );
AND2x2_ASAP7_75t_L g620 ( .A(n_574), .B(n_606), .Y(n_620) );
INVx1_ASAP7_75t_L g637 ( .A(n_574), .Y(n_637) );
INVx2_ASAP7_75t_L g653 ( .A(n_574), .Y(n_653) );
OR2x2_ASAP7_75t_L g692 ( .A(n_574), .B(n_582), .Y(n_692) );
INVx2_ASAP7_75t_L g680 ( .A(n_581), .Y(n_680) );
AND2x2_ASAP7_75t_L g604 ( .A(n_582), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g619 ( .A(n_582), .Y(n_619) );
AND2x4_ASAP7_75t_L g628 ( .A(n_582), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_582), .B(n_605), .Y(n_651) );
AND2x2_ASAP7_75t_L g758 ( .A(n_582), .B(n_653), .Y(n_758) );
INVx4_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_583), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_589), .Y(n_584) );
INVx1_ASAP7_75t_L g645 ( .A(n_591), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_592), .B(n_595), .Y(n_591) );
AND2x2_ASAP7_75t_L g732 ( .A(n_592), .B(n_659), .Y(n_732) );
INVx1_ASAP7_75t_SL g749 ( .A(n_592), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_592), .B(n_725), .Y(n_778) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OR2x2_ASAP7_75t_L g621 ( .A(n_593), .B(n_594), .Y(n_621) );
AND2x2_ASAP7_75t_L g714 ( .A(n_595), .B(n_610), .Y(n_714) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_599), .B(n_610), .Y(n_737) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_601), .A2(n_750), .B1(n_755), .B2(n_757), .Y(n_754) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
AND2x2_ASAP7_75t_L g679 ( .A(n_602), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g774 ( .A(n_602), .B(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g730 ( .A(n_603), .B(n_648), .Y(n_730) );
AND2x4_ASAP7_75t_L g684 ( .A(n_604), .B(n_630), .Y(n_684) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_606), .Y(n_782) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g615 ( .A(n_607), .Y(n_615) );
INVx1_ASAP7_75t_L g629 ( .A(n_607), .Y(n_629) );
NAND4xp25_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .C(n_611), .D(n_612), .Y(n_608) );
AND2x2_ASAP7_75t_L g766 ( .A(n_609), .B(n_751), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_609), .B(n_777), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_610), .B(n_686), .Y(n_685) );
OAI322xp33_ASAP7_75t_L g693 ( .A1(n_610), .A2(n_694), .A3(n_698), .B1(n_700), .B2(n_702), .C1(n_704), .C2(n_709), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_610), .B(n_659), .Y(n_709) );
INVx1_ASAP7_75t_L g777 ( .A(n_610), .Y(n_777) );
INVx2_ASAP7_75t_L g623 ( .A(n_611), .Y(n_623) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_614), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_615), .B(n_634), .Y(n_691) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_618), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx1_ASAP7_75t_L g664 ( .A(n_619), .Y(n_664) );
AND2x2_ASAP7_75t_L g736 ( .A(n_619), .B(n_647), .Y(n_736) );
AOI31xp33_ASAP7_75t_L g622 ( .A1(n_620), .A2(n_623), .A3(n_624), .B(n_627), .Y(n_622) );
AND2x2_ASAP7_75t_L g633 ( .A(n_620), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g761 ( .A(n_620), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_SL g768 ( .A(n_620), .B(n_648), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_620), .Y(n_769) );
INVx1_ASAP7_75t_SL g727 ( .A(n_621), .Y(n_727) );
NAND3xp33_ASAP7_75t_SL g755 ( .A(n_621), .B(n_749), .C(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g655 ( .A(n_626), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
AND2x2_ASAP7_75t_L g636 ( .A(n_628), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g697 ( .A(n_628), .Y(n_697) );
AOI322xp5_ASAP7_75t_L g779 ( .A1(n_628), .A2(n_658), .A3(n_661), .B1(n_780), .B2(n_781), .C1(n_783), .C2(n_785), .Y(n_779) );
AND2x2_ASAP7_75t_L g785 ( .A(n_628), .B(n_634), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_635), .B(n_638), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_634), .B(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g780 ( .A(n_634), .B(n_667), .Y(n_780) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g706 ( .A(n_637), .Y(n_706) );
AND2x2_ASAP7_75t_L g734 ( .A(n_637), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g781 ( .A(n_637), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g686 ( .A(n_640), .Y(n_686) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
O2A1O1Ixp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B(n_646), .C(n_649), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AND2x2_ASAP7_75t_L g703 ( .A(n_648), .B(n_653), .Y(n_703) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_654), .B(n_660), .C(n_662), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_650), .A2(n_676), .B1(n_678), .B2(n_681), .C(n_683), .Y(n_675) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g695 ( .A(n_652), .Y(n_695) );
OR2x2_ASAP7_75t_L g715 ( .A(n_652), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g760 ( .A(n_655), .Y(n_760) );
INVx1_ASAP7_75t_L g784 ( .A(n_656), .Y(n_784) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_658), .B(n_659), .Y(n_657) );
AND2x2_ASAP7_75t_L g666 ( .A(n_658), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_658), .B(n_728), .Y(n_740) );
INVx1_ASAP7_75t_L g720 ( .A(n_659), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B1(n_668), .B2(n_670), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_SL g728 ( .A(n_667), .Y(n_728) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND4xp75_ASAP7_75t_L g673 ( .A(n_674), .B(n_710), .C(n_738), .D(n_763), .Y(n_673) );
NOR2xp67_ASAP7_75t_L g674 ( .A(n_675), .B(n_693), .Y(n_674) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_SL g750 ( .A(n_682), .B(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_687), .B2(n_689), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_686), .B(n_749), .Y(n_748) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx2_ASAP7_75t_L g726 ( .A(n_692), .Y(n_726) );
OR2x2_ASAP7_75t_L g741 ( .A(n_692), .B(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g756 ( .A(n_701), .Y(n_756) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
OAI21xp5_ASAP7_75t_SL g747 ( .A1(n_703), .A2(n_748), .B(n_750), .Y(n_747) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR2x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_723), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B1(n_718), .B2(n_720), .C(n_721), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
OAI21xp33_ASAP7_75t_L g759 ( .A1(n_713), .A2(n_760), .B(n_761), .Y(n_759) );
INVx3_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
OAI322xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_727), .A3(n_728), .B1(n_729), .B2(n_731), .C1(n_733), .C2(n_737), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
NOR2x1_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g746 ( .A(n_734), .Y(n_746) );
INVx1_ASAP7_75t_L g742 ( .A(n_735), .Y(n_742) );
AND2x2_ASAP7_75t_L g757 ( .A(n_735), .B(n_758), .Y(n_757) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_752), .Y(n_738) );
OAI221xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B1(n_743), .B2(n_746), .C(n_747), .Y(n_739) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
OAI211xp5_ASAP7_75t_SL g752 ( .A1(n_746), .A2(n_753), .B(n_754), .C(n_759), .Y(n_752) );
INVx2_ASAP7_75t_SL g775 ( .A(n_762), .Y(n_775) );
NOR2x1_ASAP7_75t_L g763 ( .A(n_764), .B(n_773), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_767), .B1(n_769), .B2(n_770), .Y(n_764) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
OAI211xp5_ASAP7_75t_SL g773 ( .A1(n_774), .A2(n_776), .B(n_778), .C(n_779), .Y(n_773) );
BUFx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_798), .Y(n_791) );
INVxp67_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_794), .B(n_797), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_795), .A2(n_804), .B(n_807), .Y(n_803) );
OR2x2_ASAP7_75t_SL g824 ( .A(n_795), .B(n_797), .Y(n_824) );
INVx1_ASAP7_75t_L g821 ( .A(n_798), .Y(n_821) );
BUFx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
BUFx2_ASAP7_75t_L g808 ( .A(n_799), .Y(n_808) );
BUFx2_ASAP7_75t_R g811 ( .A(n_799), .Y(n_811) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
CKINVDCx11_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
CKINVDCx8_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
O2A1O1Ixp33_ASAP7_75t_SL g809 ( .A1(n_810), .A2(n_812), .B(n_820), .C(n_822), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
XNOR2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
XOR2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
endmodule