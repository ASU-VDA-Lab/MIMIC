module fake_netlist_1_6198_n_1284 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1284);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1284;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_271;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_265;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_272;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_266;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_267;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_270;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_264;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_584;
wire n_1130;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_269;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_274;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_262;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_263;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_261;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g261 ( .A(n_24), .Y(n_261) );
INVxp67_ASAP7_75t_L g262 ( .A(n_233), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_159), .Y(n_263) );
INVxp33_ASAP7_75t_L g264 ( .A(n_203), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_1), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_154), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_229), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_147), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_131), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_119), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_80), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_230), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_88), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_122), .B(n_195), .Y(n_274) );
INVxp33_ASAP7_75t_L g275 ( .A(n_169), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_45), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_225), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_259), .Y(n_278) );
INVxp33_ASAP7_75t_L g279 ( .A(n_249), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_192), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_43), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_79), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_156), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_62), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_191), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_12), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_103), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_34), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_189), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_151), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_118), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_83), .Y(n_292) );
INVxp33_ASAP7_75t_SL g293 ( .A(n_115), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_238), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_190), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_200), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_94), .Y(n_297) );
CKINVDCx16_ASAP7_75t_R g298 ( .A(n_144), .Y(n_298) );
INVxp33_ASAP7_75t_SL g299 ( .A(n_141), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_123), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_227), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_187), .Y(n_302) );
INVxp67_ASAP7_75t_SL g303 ( .A(n_60), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_0), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_95), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_185), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_51), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_250), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_107), .Y(n_309) );
BUFx5_ASAP7_75t_L g310 ( .A(n_175), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_213), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_63), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_8), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_215), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_105), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_136), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_67), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_176), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_29), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_63), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_31), .Y(n_322) );
CKINVDCx16_ASAP7_75t_R g323 ( .A(n_222), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_163), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_174), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_106), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_193), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_38), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_10), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_132), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_0), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_26), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_188), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_153), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_17), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_121), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_140), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_26), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_138), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_90), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_155), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_91), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_35), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_166), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_85), .Y(n_345) );
CKINVDCx14_ASAP7_75t_R g346 ( .A(n_16), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_28), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_207), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_41), .Y(n_349) );
INVxp33_ASAP7_75t_L g350 ( .A(n_33), .Y(n_350) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_78), .Y(n_351) );
INVxp33_ASAP7_75t_L g352 ( .A(n_208), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_142), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_245), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_194), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_134), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_205), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_167), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g359 ( .A(n_157), .Y(n_359) );
BUFx2_ASAP7_75t_SL g360 ( .A(n_46), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_31), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_210), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_74), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_76), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_46), .Y(n_365) );
INVxp67_ASAP7_75t_L g366 ( .A(n_241), .Y(n_366) );
NOR2xp67_ASAP7_75t_L g367 ( .A(n_100), .B(n_54), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_127), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_73), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_29), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_110), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_87), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_247), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_54), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_43), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_116), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_124), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_246), .Y(n_378) );
INVxp33_ASAP7_75t_L g379 ( .A(n_67), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_20), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_164), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_93), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_184), .Y(n_383) );
CKINVDCx16_ASAP7_75t_R g384 ( .A(n_55), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_239), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_99), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_42), .Y(n_387) );
INVxp33_ASAP7_75t_SL g388 ( .A(n_114), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_81), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_234), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_7), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_11), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_25), .Y(n_393) );
BUFx5_ASAP7_75t_L g394 ( .A(n_23), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_125), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_59), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_30), .Y(n_397) );
CKINVDCx6p67_ASAP7_75t_R g398 ( .A(n_9), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_49), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_310), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_286), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_286), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_286), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_298), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_394), .Y(n_405) );
OAI22x1_ASAP7_75t_R g406 ( .A1(n_392), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_346), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_309), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_350), .B(n_2), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_394), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_346), .Y(n_411) );
OA21x2_ASAP7_75t_L g412 ( .A1(n_297), .A2(n_77), .B(n_75), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_316), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_350), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_379), .B(n_3), .Y(n_415) );
INVx3_ASAP7_75t_L g416 ( .A(n_394), .Y(n_416) );
BUFx8_ASAP7_75t_L g417 ( .A(n_310), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_394), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_310), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_310), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_394), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_394), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_394), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_304), .Y(n_424) );
NAND2xp33_ASAP7_75t_L g425 ( .A(n_310), .B(n_82), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_285), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_304), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_380), .Y(n_428) );
INVxp67_ASAP7_75t_L g429 ( .A(n_315), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_379), .B(n_4), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_323), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_380), .B(n_4), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_351), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_266), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_264), .B(n_5), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_407), .B(n_264), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_429), .B(n_275), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_408), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g439 ( .A(n_415), .B(n_384), .C(n_343), .Y(n_439) );
INVx4_ASAP7_75t_L g440 ( .A(n_432), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_429), .B(n_275), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_414), .B(n_279), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_416), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_407), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_409), .A2(n_265), .B1(n_276), .B2(n_261), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_416), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_408), .Y(n_447) );
INVx5_ASAP7_75t_L g448 ( .A(n_416), .Y(n_448) );
INVx4_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_416), .Y(n_450) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_435), .B(n_274), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_426), .B(n_279), .Y(n_452) );
INVx5_ASAP7_75t_L g453 ( .A(n_416), .Y(n_453) );
INVx6_ASAP7_75t_L g454 ( .A(n_417), .Y(n_454) );
AO22x2_ASAP7_75t_L g455 ( .A1(n_432), .A2(n_360), .B1(n_332), .B2(n_303), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_414), .B(n_352), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_426), .B(n_435), .Y(n_457) );
NAND2xp33_ASAP7_75t_L g458 ( .A(n_435), .B(n_310), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_405), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_409), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_434), .B(n_348), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_417), .B(n_306), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_405), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_417), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_401), .B(n_336), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_409), .A2(n_284), .B1(n_318), .B2(n_281), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_404), .B(n_262), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_430), .A2(n_320), .B1(n_329), .B2(n_322), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_410), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_413), .B(n_366), .Y(n_470) );
BUFx4f_ASAP7_75t_L g471 ( .A(n_432), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g472 ( .A(n_432), .B(n_268), .Y(n_472) );
BUFx3_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_401), .B(n_312), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_430), .B(n_307), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_410), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_417), .B(n_431), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_433), .B(n_306), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_402), .B(n_335), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_418), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_400), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_481), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_460), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_444), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_442), .B(n_415), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_454), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_481), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_440), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_440), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_440), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_449), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_444), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_455), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_455), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_457), .B(n_430), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_437), .B(n_402), .Y(n_496) );
BUFx12f_ASAP7_75t_L g497 ( .A(n_451), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_455), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_456), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_441), .B(n_398), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_451), .A2(n_272), .B1(n_291), .B2(n_283), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_465), .B(n_403), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_465), .B(n_403), .Y(n_503) );
OAI22xp5_ASAP7_75t_SL g504 ( .A1(n_445), .A2(n_392), .B1(n_411), .B2(n_272), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_449), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_455), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_479), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_439), .B(n_425), .C(n_313), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_464), .B(n_400), .Y(n_509) );
NOR3xp33_ASAP7_75t_SL g510 ( .A(n_478), .B(n_313), .C(n_312), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_464), .B(n_400), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_465), .B(n_428), .Y(n_512) );
NOR2x2_ASAP7_75t_L g513 ( .A(n_451), .B(n_411), .Y(n_513) );
NOR2x2_ASAP7_75t_L g514 ( .A(n_475), .B(n_406), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_454), .Y(n_515) );
NOR3xp33_ASAP7_75t_SL g516 ( .A(n_467), .B(n_321), .C(n_288), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_449), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_479), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_475), .B(n_328), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_471), .B(n_419), .Y(n_520) );
AOI22x1_ASAP7_75t_L g521 ( .A1(n_472), .A2(n_419), .B1(n_420), .B2(n_418), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_479), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_452), .B(n_293), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_471), .B(n_419), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_474), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_443), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_461), .B(n_353), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_473), .B(n_424), .Y(n_528) );
OAI21xp33_ASAP7_75t_L g529 ( .A1(n_466), .A2(n_422), .B(n_421), .Y(n_529) );
INVx4_ASAP7_75t_L g530 ( .A(n_454), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_436), .B(n_356), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_472), .B(n_356), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_471), .A2(n_421), .B1(n_423), .B2(n_422), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_468), .A2(n_291), .B1(n_359), .B2(n_283), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_458), .B(n_425), .C(n_387), .Y(n_535) );
INVx2_ASAP7_75t_SL g536 ( .A(n_472), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_454), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_470), .B(n_349), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_473), .B(n_420), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_446), .B(n_371), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_446), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_443), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_450), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_477), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_450), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_462), .A2(n_359), .B1(n_376), .B2(n_373), .Y(n_546) );
INVx2_ASAP7_75t_SL g547 ( .A(n_448), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_448), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_459), .B(n_293), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_459), .A2(n_373), .B1(n_385), .B2(n_376), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_463), .B(n_420), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_463), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_469), .B(n_385), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_469), .B(n_370), .Y(n_554) );
INVxp33_ASAP7_75t_SL g555 ( .A(n_476), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_480), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_448), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_448), .A2(n_388), .B1(n_299), .B2(n_338), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_448), .A2(n_388), .B1(n_299), .B2(n_361), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_448), .B(n_423), .Y(n_561) );
AND2x6_ASAP7_75t_SL g562 ( .A(n_438), .B(n_406), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_453), .B(n_424), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_453), .B(n_427), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_453), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_453), .B(n_270), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_453), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_453), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_438), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_485), .B(n_427), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_501), .A2(n_550), .B1(n_534), .B2(n_497), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_553), .B(n_347), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_500), .B(n_363), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_488), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_488), .Y(n_575) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_486), .Y(n_576) );
AND2x6_ASAP7_75t_L g577 ( .A(n_493), .B(n_273), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_495), .B(n_365), .Y(n_578) );
BUFx2_ASAP7_75t_SL g579 ( .A(n_484), .Y(n_579) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_486), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_507), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_552), .A2(n_412), .B(n_277), .Y(n_582) );
NOR2xp33_ASAP7_75t_R g583 ( .A(n_497), .B(n_499), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_506), .A2(n_369), .B1(n_375), .B2(n_374), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_495), .B(n_391), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_492), .B(n_393), .Y(n_586) );
INVx5_ASAP7_75t_L g587 ( .A(n_536), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_494), .A2(n_397), .B1(n_399), .B2(n_396), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_489), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_525), .B(n_367), .Y(n_590) );
INVx3_ASAP7_75t_L g591 ( .A(n_490), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_490), .Y(n_592) );
OR2x6_ASAP7_75t_SL g593 ( .A(n_546), .B(n_263), .Y(n_593) );
AO22x1_ASAP7_75t_L g594 ( .A1(n_553), .A2(n_269), .B1(n_300), .B2(n_267), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_555), .B(n_317), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_562), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_498), .A2(n_278), .B(n_280), .C(n_271), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_518), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g599 ( .A1(n_483), .A2(n_282), .B(n_289), .C(n_287), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_489), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_509), .A2(n_412), .B(n_294), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_522), .Y(n_602) );
BUFx2_ASAP7_75t_L g603 ( .A(n_499), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_528), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_530), .B(n_325), .Y(n_605) );
BUFx3_ASAP7_75t_L g606 ( .A(n_563), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_519), .B(n_331), .Y(n_607) );
INVx3_ASAP7_75t_L g608 ( .A(n_491), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_496), .B(n_337), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_502), .B(n_342), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_491), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_505), .Y(n_612) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_486), .Y(n_613) );
OR2x6_ASAP7_75t_L g614 ( .A(n_504), .B(n_331), .Y(n_614) );
OAI21x1_ASAP7_75t_L g615 ( .A1(n_521), .A2(n_412), .B(n_302), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_503), .B(n_382), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_528), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_511), .A2(n_412), .B(n_295), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_557), .A2(n_290), .B(n_301), .C(n_296), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_544), .B(n_305), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_530), .B(n_314), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_505), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_517), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_513), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_529), .A2(n_508), .B1(n_512), .B2(n_554), .Y(n_625) );
OAI22xp5_ASAP7_75t_SL g626 ( .A1(n_514), .A2(n_326), .B1(n_327), .B2(n_324), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_517), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_549), .B(n_333), .Y(n_628) );
INVx4_ASAP7_75t_L g629 ( .A(n_528), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_537), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_486), .B(n_334), .Y(n_631) );
BUFx12f_ASAP7_75t_L g632 ( .A(n_514), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_532), .Y(n_633) );
INVx2_ASAP7_75t_SL g634 ( .A(n_531), .Y(n_634) );
AO31x2_ASAP7_75t_L g635 ( .A1(n_556), .A2(n_302), .A3(n_308), .B(n_297), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_520), .A2(n_341), .B(n_340), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_556), .A2(n_354), .B1(n_368), .B2(n_344), .Y(n_637) );
AND2x2_ASAP7_75t_SL g638 ( .A(n_513), .B(n_372), .Y(n_638) );
NOR2xp33_ASAP7_75t_R g639 ( .A(n_523), .B(n_5), .Y(n_639) );
CKINVDCx6p67_ASAP7_75t_R g640 ( .A(n_538), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_515), .B(n_378), .Y(n_641) );
INVx3_ASAP7_75t_SL g642 ( .A(n_566), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_559), .B(n_6), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_515), .B(n_273), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_535), .A2(n_386), .B1(n_390), .B2(n_381), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_523), .B(n_395), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_541), .Y(n_647) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_515), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_516), .B(n_510), .Y(n_649) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_547), .Y(n_650) );
BUFx3_ASAP7_75t_L g651 ( .A(n_564), .Y(n_651) );
INVx4_ASAP7_75t_L g652 ( .A(n_568), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_560), .B(n_292), .Y(n_653) );
OR2x6_ASAP7_75t_L g654 ( .A(n_524), .B(n_308), .Y(n_654) );
BUFx3_ASAP7_75t_L g655 ( .A(n_558), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_542), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_527), .B(n_6), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_540), .B(n_7), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_548), .B(n_292), .Y(n_659) );
NAND2x2_ASAP7_75t_L g660 ( .A(n_566), .B(n_319), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_543), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_482), .Y(n_662) );
AOI222xp33_ASAP7_75t_L g663 ( .A1(n_533), .A2(n_339), .B1(n_383), .B2(n_319), .C1(n_330), .C2(n_357), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_545), .Y(n_664) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_487), .Y(n_665) );
INVx4_ASAP7_75t_L g666 ( .A(n_568), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_533), .A2(n_345), .B1(n_357), .B2(n_355), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_526), .Y(n_668) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_487), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_526), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_565), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g672 ( .A1(n_567), .A2(n_383), .B1(n_339), .B2(n_355), .Y(n_672) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_539), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_551), .A2(n_358), .B(n_345), .Y(n_674) );
NAND3xp33_ASAP7_75t_SL g675 ( .A(n_561), .B(n_364), .C(n_362), .Y(n_675) );
CKINVDCx16_ASAP7_75t_R g676 ( .A(n_569), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_561), .B(n_9), .Y(n_677) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_569), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_506), .A2(n_364), .B1(n_362), .B2(n_377), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_501), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_485), .B(n_377), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_485), .B(n_10), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_495), .A2(n_389), .B(n_311), .C(n_309), .Y(n_683) );
AND2x4_ASAP7_75t_L g684 ( .A(n_525), .B(n_11), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_506), .A2(n_310), .B1(n_389), .B2(n_311), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_497), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_485), .B(n_12), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_555), .B(n_309), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_488), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g690 ( .A(n_536), .B(n_84), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_500), .B(n_13), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_488), .Y(n_692) );
OAI21x1_ASAP7_75t_L g693 ( .A1(n_615), .A2(n_311), .B(n_309), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_614), .A2(n_687), .B1(n_682), .B2(n_684), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_614), .A2(n_389), .B1(n_311), .B2(n_408), .Y(n_695) );
BUFx3_ASAP7_75t_L g696 ( .A(n_603), .Y(n_696) );
INVx1_ASAP7_75t_SL g697 ( .A(n_676), .Y(n_697) );
AND2x4_ASAP7_75t_L g698 ( .A(n_587), .B(n_14), .Y(n_698) );
OAI21x1_ASAP7_75t_L g699 ( .A1(n_582), .A2(n_389), .B(n_408), .Y(n_699) );
AO21x2_ASAP7_75t_L g700 ( .A1(n_582), .A2(n_408), .B(n_438), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_607), .Y(n_701) );
OAI21x1_ASAP7_75t_L g702 ( .A1(n_601), .A2(n_408), .B(n_438), .Y(n_702) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_678), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_570), .Y(n_704) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_676), .Y(n_705) );
INVx3_ASAP7_75t_L g706 ( .A(n_587), .Y(n_706) );
AO21x2_ASAP7_75t_L g707 ( .A1(n_683), .A2(n_408), .B(n_447), .Y(n_707) );
OR2x4_ASAP7_75t_L g708 ( .A(n_643), .B(n_14), .Y(n_708) );
INVx3_ASAP7_75t_L g709 ( .A(n_587), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_684), .A2(n_447), .B1(n_16), .B2(n_17), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_618), .A2(n_447), .B(n_89), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_638), .B(n_15), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_662), .Y(n_713) );
OAI21x1_ASAP7_75t_L g714 ( .A1(n_644), .A2(n_92), .B(n_86), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_583), .Y(n_715) );
AO32x2_ASAP7_75t_L g716 ( .A1(n_667), .A2(n_15), .A3(n_18), .B1(n_19), .B2(n_20), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_632), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_614), .A2(n_18), .B1(n_19), .B2(n_21), .Y(n_718) );
OR2x6_ASAP7_75t_L g719 ( .A(n_579), .B(n_21), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_647), .B(n_22), .Y(n_720) );
BUFx12f_ASAP7_75t_L g721 ( .A(n_596), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_581), .B(n_22), .Y(n_722) );
INVxp67_ASAP7_75t_SL g723 ( .A(n_662), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_586), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_633), .B(n_23), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_598), .B(n_24), .Y(n_726) );
OAI21x1_ASAP7_75t_L g727 ( .A1(n_674), .A2(n_97), .B(n_96), .Y(n_727) );
INVx1_ASAP7_75t_SL g728 ( .A(n_604), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_680), .A2(n_571), .B1(n_604), .B2(n_640), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_679), .A2(n_25), .B1(n_27), .B2(n_28), .Y(n_730) );
BUFx12f_ASAP7_75t_L g731 ( .A(n_624), .Y(n_731) );
OAI21x1_ASAP7_75t_L g732 ( .A1(n_674), .A2(n_101), .B(n_98), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_649), .A2(n_27), .B1(n_30), .B2(n_32), .Y(n_733) );
AND2x2_ASAP7_75t_SL g734 ( .A(n_629), .B(n_32), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_602), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_670), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_608), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_656), .Y(n_738) );
AOI22x1_ASAP7_75t_L g739 ( .A1(n_663), .A2(n_152), .B1(n_258), .B2(n_257), .Y(n_739) );
OR2x2_ASAP7_75t_L g740 ( .A(n_572), .B(n_33), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_661), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_679), .A2(n_588), .B1(n_625), .B2(n_593), .Y(n_742) );
OAI21x1_ASAP7_75t_L g743 ( .A1(n_690), .A2(n_104), .B(n_102), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_573), .B(n_34), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_691), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_745) );
OAI21x1_ASAP7_75t_L g746 ( .A1(n_690), .A2(n_109), .B(n_108), .Y(n_746) );
AND2x4_ASAP7_75t_L g747 ( .A(n_634), .B(n_36), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_664), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_681), .B(n_37), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_608), .Y(n_750) );
AND2x4_ASAP7_75t_L g751 ( .A(n_629), .B(n_38), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_677), .Y(n_752) );
CKINVDCx11_ASAP7_75t_R g753 ( .A(n_660), .Y(n_753) );
OAI21x1_ASAP7_75t_L g754 ( .A1(n_631), .A2(n_112), .B(n_111), .Y(n_754) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_578), .A2(n_39), .B1(n_40), .B2(n_41), .C(n_42), .Y(n_755) );
OAI21x1_ASAP7_75t_L g756 ( .A1(n_641), .A2(n_171), .B(n_256), .Y(n_756) );
BUFx3_ASAP7_75t_L g757 ( .A(n_606), .Y(n_757) );
OAI211xp5_ASAP7_75t_L g758 ( .A1(n_639), .A2(n_39), .B(n_40), .C(n_44), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_678), .B(n_44), .Y(n_759) );
OAI21xp5_ASAP7_75t_L g760 ( .A1(n_625), .A2(n_45), .B(n_47), .Y(n_760) );
NAND2x1p5_ASAP7_75t_L g761 ( .A(n_651), .B(n_47), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_588), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_762) );
BUFx2_ASAP7_75t_R g763 ( .A(n_595), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_611), .Y(n_764) );
INVx3_ASAP7_75t_L g765 ( .A(n_650), .Y(n_765) );
NAND2x1p5_ASAP7_75t_L g766 ( .A(n_678), .B(n_48), .Y(n_766) );
NAND2x1p5_ASAP7_75t_L g767 ( .A(n_652), .B(n_50), .Y(n_767) );
AND2x2_ASAP7_75t_SL g768 ( .A(n_649), .B(n_51), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_626), .A2(n_52), .B1(n_53), .B2(n_55), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_574), .Y(n_770) );
OAI21x1_ASAP7_75t_L g771 ( .A1(n_636), .A2(n_173), .B(n_255), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_575), .Y(n_772) );
AO21x2_ASAP7_75t_L g773 ( .A1(n_675), .A2(n_172), .B(n_254), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_612), .Y(n_774) );
OA21x2_ASAP7_75t_L g775 ( .A1(n_685), .A2(n_170), .B(n_253), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_622), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_589), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_623), .Y(n_778) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_626), .Y(n_779) );
OAI21x1_ASAP7_75t_L g780 ( .A1(n_668), .A2(n_168), .B(n_252), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_585), .B(n_52), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_658), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_597), .A2(n_53), .B(n_56), .Y(n_783) );
INVx1_ASAP7_75t_SL g784 ( .A(n_665), .Y(n_784) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_619), .A2(n_599), .B(n_646), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_590), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_628), .A2(n_165), .B(n_251), .Y(n_787) );
NAND3xp33_ASAP7_75t_L g788 ( .A(n_663), .B(n_56), .C(n_57), .Y(n_788) );
BUFx3_ASAP7_75t_L g789 ( .A(n_650), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_594), .Y(n_790) );
AND2x2_ASAP7_75t_SL g791 ( .A(n_617), .B(n_57), .Y(n_791) );
AND2x4_ASAP7_75t_L g792 ( .A(n_620), .B(n_58), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_642), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_600), .Y(n_794) );
INVx3_ASAP7_75t_SL g795 ( .A(n_659), .Y(n_795) );
OAI222xp33_ASAP7_75t_L g796 ( .A1(n_654), .A2(n_58), .B1(n_59), .B2(n_60), .C1(n_61), .C2(n_62), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_627), .Y(n_797) );
BUFx6f_ASAP7_75t_L g798 ( .A(n_576), .Y(n_798) );
AOI21xp33_ASAP7_75t_L g799 ( .A1(n_654), .A2(n_61), .B(n_64), .Y(n_799) );
OR2x2_ASAP7_75t_L g800 ( .A(n_620), .B(n_609), .Y(n_800) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_665), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_653), .A2(n_178), .B(n_244), .Y(n_802) );
AND2x4_ASAP7_75t_L g803 ( .A(n_590), .B(n_64), .Y(n_803) );
OR2x6_ASAP7_75t_L g804 ( .A(n_654), .B(n_65), .Y(n_804) );
OAI21xp5_ASAP7_75t_L g805 ( .A1(n_645), .A2(n_65), .B(n_66), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_689), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_657), .A2(n_66), .B1(n_68), .B2(n_69), .Y(n_807) );
INVx2_ASAP7_75t_SL g808 ( .A(n_659), .Y(n_808) );
OAI21xp33_ASAP7_75t_SL g809 ( .A1(n_688), .A2(n_68), .B(n_69), .Y(n_809) );
AO31x2_ASAP7_75t_L g810 ( .A1(n_645), .A2(n_70), .A3(n_71), .B(n_72), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_584), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_610), .B(n_73), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_692), .Y(n_813) );
A2O1A1Ixp33_ASAP7_75t_L g814 ( .A1(n_591), .A2(n_74), .B(n_113), .C(n_117), .Y(n_814) );
AND2x4_ASAP7_75t_L g815 ( .A(n_591), .B(n_260), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_665), .B(n_120), .Y(n_816) );
OAI21x1_ASAP7_75t_L g817 ( .A1(n_630), .A2(n_126), .B(n_128), .Y(n_817) );
BUFx2_ASAP7_75t_L g818 ( .A(n_652), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_669), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_616), .B(n_129), .Y(n_820) );
INVx3_ASAP7_75t_L g821 ( .A(n_650), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_637), .Y(n_822) );
AND2x4_ASAP7_75t_L g823 ( .A(n_592), .B(n_130), .Y(n_823) );
INVx2_ASAP7_75t_SL g824 ( .A(n_655), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_738), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_741), .Y(n_826) );
AND2x4_ASAP7_75t_L g827 ( .A(n_706), .B(n_592), .Y(n_827) );
AOI21x1_ASAP7_75t_L g828 ( .A1(n_693), .A2(n_621), .B(n_605), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_742), .A2(n_577), .B1(n_671), .B2(n_672), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_704), .B(n_577), .Y(n_830) );
CKINVDCx8_ASAP7_75t_R g831 ( .A(n_717), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_748), .Y(n_832) );
AO21x2_ASAP7_75t_L g833 ( .A1(n_700), .A2(n_635), .B(n_577), .Y(n_833) );
NAND2xp5_ASAP7_75t_SL g834 ( .A(n_791), .B(n_669), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_742), .A2(n_791), .B1(n_734), .B2(n_768), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_724), .B(n_577), .Y(n_836) );
OAI221xp5_ASAP7_75t_L g837 ( .A1(n_729), .A2(n_666), .B1(n_673), .B2(n_648), .C(n_613), .Y(n_837) );
AO31x2_ASAP7_75t_L g838 ( .A1(n_711), .A2(n_635), .A3(n_666), .B(n_648), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g839 ( .A1(n_708), .A2(n_673), .B1(n_648), .B2(n_613), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g840 ( .A1(n_734), .A2(n_673), .B1(n_613), .B2(n_580), .Y(n_840) );
OAI21x1_ASAP7_75t_L g841 ( .A1(n_702), .A2(n_635), .B(n_580), .Y(n_841) );
A2O1A1Ixp33_ASAP7_75t_L g842 ( .A1(n_812), .A2(n_785), .B(n_788), .C(n_783), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_720), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_736), .B(n_752), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_720), .Y(n_845) );
AOI221xp5_ASAP7_75t_L g846 ( .A1(n_785), .A2(n_133), .B1(n_135), .B2(n_137), .C(n_139), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_804), .A2(n_143), .B1(n_145), .B2(n_146), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_736), .B(n_735), .Y(n_848) );
AOI21xp33_ASAP7_75t_L g849 ( .A1(n_812), .A2(n_148), .B(n_149), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_705), .B(n_150), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g851 ( .A1(n_723), .A2(n_158), .B(n_160), .Y(n_851) );
OAI21xp33_ASAP7_75t_L g852 ( .A1(n_760), .A2(n_161), .B(n_162), .Y(n_852) );
INVx4_ASAP7_75t_SL g853 ( .A(n_719), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_722), .Y(n_854) );
OAI22xp5_ASAP7_75t_SL g855 ( .A1(n_779), .A2(n_177), .B1(n_179), .B2(n_180), .Y(n_855) );
AOI21xp5_ASAP7_75t_L g856 ( .A1(n_723), .A2(n_181), .B(n_182), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_804), .A2(n_183), .B1(n_186), .B2(n_196), .Y(n_857) );
OAI21xp5_ASAP7_75t_SL g858 ( .A1(n_769), .A2(n_197), .B(n_198), .Y(n_858) );
OAI22xp5_ASAP7_75t_SL g859 ( .A1(n_708), .A2(n_199), .B1(n_201), .B2(n_202), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_804), .A2(n_204), .B1(n_206), .B2(n_209), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_792), .A2(n_211), .B1(n_212), .B2(n_214), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_764), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_792), .A2(n_216), .B1(n_217), .B2(n_218), .Y(n_863) );
OAI221xp5_ASAP7_75t_L g864 ( .A1(n_694), .A2(n_219), .B1(n_220), .B2(n_221), .C(n_223), .Y(n_864) );
AND2x2_ASAP7_75t_SL g865 ( .A(n_715), .B(n_224), .Y(n_865) );
AO31x2_ASAP7_75t_L g866 ( .A1(n_802), .A2(n_710), .A3(n_787), .B(n_816), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_710), .A2(n_226), .B1(n_228), .B2(n_231), .Y(n_867) );
AOI22xp33_ASAP7_75t_SL g868 ( .A1(n_712), .A2(n_232), .B1(n_235), .B2(n_236), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_774), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_697), .B(n_237), .Y(n_870) );
AO22x1_ASAP7_75t_L g871 ( .A1(n_790), .A2(n_243), .B1(n_240), .B2(n_242), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_722), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_705), .B(n_697), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_694), .A2(n_747), .B1(n_719), .B2(n_800), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_696), .B(n_795), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_747), .A2(n_719), .B1(n_725), .B2(n_803), .Y(n_876) );
NAND2xp33_ASAP7_75t_R g877 ( .A(n_698), .B(n_751), .Y(n_877) );
INVx3_ASAP7_75t_L g878 ( .A(n_789), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_782), .B(n_725), .Y(n_879) );
INVx3_ASAP7_75t_L g880 ( .A(n_703), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_803), .A2(n_744), .B1(n_751), .B2(n_822), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_758), .A2(n_761), .B1(n_730), .B2(n_698), .Y(n_882) );
A2O1A1Ixp33_ASAP7_75t_L g883 ( .A1(n_783), .A2(n_760), .B(n_781), .C(n_805), .Y(n_883) );
AOI21xp33_ASAP7_75t_L g884 ( .A1(n_749), .A2(n_781), .B(n_808), .Y(n_884) );
CKINVDCx11_ASAP7_75t_R g885 ( .A(n_721), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_795), .A2(n_740), .B1(n_730), .B2(n_761), .Y(n_886) );
BUFx2_ASAP7_75t_L g887 ( .A(n_793), .Y(n_887) );
AOI222xp33_ASAP7_75t_L g888 ( .A1(n_769), .A2(n_762), .B1(n_755), .B2(n_805), .C1(n_811), .C2(n_796), .Y(n_888) );
OAI221xp5_ASAP7_75t_L g889 ( .A1(n_786), .A2(n_718), .B1(n_733), .B2(n_807), .C(n_745), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_731), .Y(n_890) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_762), .A2(n_767), .B1(n_811), .B2(n_728), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_767), .A2(n_718), .B1(n_728), .B2(n_733), .Y(n_892) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_818), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_776), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_713), .A2(n_778), .B1(n_726), .B2(n_766), .Y(n_895) );
INVxp67_ASAP7_75t_L g896 ( .A(n_757), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g897 ( .A(n_753), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_701), .A2(n_755), .B1(n_726), .B2(n_799), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_799), .A2(n_820), .B1(n_759), .B2(n_739), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_758), .A2(n_809), .B1(n_813), .B2(n_806), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_824), .B(n_706), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_815), .A2(n_823), .B1(n_750), .B2(n_737), .Y(n_902) );
AND2x4_ASAP7_75t_L g903 ( .A(n_709), .B(n_815), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_823), .A2(n_709), .B1(n_695), .B2(n_794), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_763), .B(n_716), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_770), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_695), .A2(n_772), .B1(n_777), .B2(n_797), .Y(n_907) );
OA21x2_ASAP7_75t_L g908 ( .A1(n_727), .A2(n_732), .B(n_780), .Y(n_908) );
OR2x2_ASAP7_75t_L g909 ( .A(n_765), .B(n_821), .Y(n_909) );
NAND2xp5_ASAP7_75t_SL g910 ( .A(n_703), .B(n_784), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_766), .A2(n_765), .B1(n_821), .B2(n_801), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_801), .A2(n_819), .B1(n_703), .B2(n_775), .Y(n_912) );
A2O1A1Ixp33_ASAP7_75t_L g913 ( .A1(n_814), .A2(n_743), .B(n_746), .C(n_771), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_707), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_763), .A2(n_819), .B1(n_798), .B2(n_775), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_716), .Y(n_916) );
AOI221xp5_ASAP7_75t_L g917 ( .A1(n_796), .A2(n_773), .B1(n_798), .B2(n_716), .C(n_810), .Y(n_917) );
AOI22xp33_ASAP7_75t_SL g918 ( .A1(n_817), .A2(n_714), .B1(n_754), .B2(n_756), .Y(n_918) );
AND2x4_ASAP7_75t_L g919 ( .A(n_798), .B(n_810), .Y(n_919) );
OA21x2_ASAP7_75t_L g920 ( .A1(n_810), .A2(n_693), .B(n_699), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_742), .A2(n_614), .B1(n_638), .B2(n_791), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_704), .A2(n_571), .B1(n_573), .B2(n_724), .C(n_742), .Y(n_922) );
AOI21xp33_ASAP7_75t_L g923 ( .A1(n_742), .A2(n_812), .B(n_785), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_694), .A2(n_804), .B1(n_742), .B2(n_501), .Y(n_924) );
AO21x2_ASAP7_75t_L g925 ( .A1(n_700), .A2(n_711), .B(n_699), .Y(n_925) );
AND2x4_ASAP7_75t_L g926 ( .A(n_706), .B(n_686), .Y(n_926) );
AND2x4_ASAP7_75t_L g927 ( .A(n_706), .B(n_686), .Y(n_927) );
AND2x4_ASAP7_75t_L g928 ( .A(n_706), .B(n_686), .Y(n_928) );
INVx11_ASAP7_75t_L g929 ( .A(n_721), .Y(n_929) );
BUFx6f_ASAP7_75t_L g930 ( .A(n_703), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_768), .B(n_638), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_704), .B(n_485), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_738), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_768), .B(n_638), .Y(n_934) );
AO21x2_ASAP7_75t_L g935 ( .A1(n_700), .A2(n_711), .B(n_699), .Y(n_935) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_768), .A2(n_501), .B1(n_791), .B2(n_734), .Y(n_936) );
OAI211xp5_ASAP7_75t_SL g937 ( .A1(n_769), .A2(n_516), .B(n_729), .C(n_510), .Y(n_937) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_739), .B(n_760), .C(n_758), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_738), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_694), .A2(n_804), .B1(n_734), .B2(n_742), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_738), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_742), .A2(n_614), .B1(n_638), .B2(n_791), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_738), .Y(n_943) );
BUFx3_ASAP7_75t_L g944 ( .A(n_793), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g945 ( .A1(n_704), .A2(n_571), .B1(n_573), .B2(n_724), .C(n_742), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_704), .B(n_485), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_906), .B(n_862), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_841), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_914), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_916), .Y(n_950) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_893), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_869), .B(n_894), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_920), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_940), .B(n_835), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_931), .B(n_934), .Y(n_955) );
INVx3_ASAP7_75t_L g956 ( .A(n_930), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_843), .B(n_845), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_940), .B(n_854), .Y(n_958) );
CKINVDCx8_ASAP7_75t_R g959 ( .A(n_853), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_838), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_872), .B(n_825), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_933), .B(n_943), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_838), .Y(n_963) );
OR2x2_ASAP7_75t_L g964 ( .A(n_924), .B(n_848), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_826), .B(n_832), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_838), .Y(n_966) );
INVx1_ASAP7_75t_SL g967 ( .A(n_903), .Y(n_967) );
INVx2_ASAP7_75t_L g968 ( .A(n_925), .Y(n_968) );
BUFx6f_ASAP7_75t_L g969 ( .A(n_930), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_939), .Y(n_970) );
AND2x2_ASAP7_75t_L g971 ( .A(n_941), .B(n_923), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_919), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_919), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_883), .B(n_842), .Y(n_974) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_926), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_921), .B(n_942), .Y(n_976) );
INVx3_ASAP7_75t_L g977 ( .A(n_930), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_922), .B(n_945), .Y(n_978) );
OR2x2_ASAP7_75t_L g979 ( .A(n_844), .B(n_874), .Y(n_979) );
INVx2_ASAP7_75t_SL g980 ( .A(n_926), .Y(n_980) );
INVx1_ASAP7_75t_SL g981 ( .A(n_903), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_936), .B(n_888), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_927), .Y(n_983) );
INVx3_ASAP7_75t_L g984 ( .A(n_880), .Y(n_984) );
INVx2_ASAP7_75t_SL g985 ( .A(n_927), .Y(n_985) );
BUFx3_ASAP7_75t_L g986 ( .A(n_928), .Y(n_986) );
OR2x2_ASAP7_75t_L g987 ( .A(n_881), .B(n_834), .Y(n_987) );
INVx5_ASAP7_75t_L g988 ( .A(n_880), .Y(n_988) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_928), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_888), .B(n_898), .Y(n_990) );
BUFx2_ASAP7_75t_L g991 ( .A(n_853), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_925), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_882), .B(n_865), .Y(n_993) );
HB1xp67_ASAP7_75t_L g994 ( .A(n_873), .Y(n_994) );
OAI222xp33_ASAP7_75t_L g995 ( .A1(n_891), .A2(n_892), .B1(n_886), .B2(n_840), .C1(n_889), .C2(n_876), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_895), .Y(n_996) );
OR2x2_ASAP7_75t_L g997 ( .A(n_879), .B(n_932), .Y(n_997) );
INVx3_ASAP7_75t_L g998 ( .A(n_833), .Y(n_998) );
AND2x4_ASAP7_75t_L g999 ( .A(n_910), .B(n_900), .Y(n_999) );
INVx3_ASAP7_75t_SL g1000 ( .A(n_890), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_833), .Y(n_1001) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_878), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_900), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_877), .Y(n_1004) );
BUFx3_ASAP7_75t_L g1005 ( .A(n_878), .Y(n_1005) );
INVx2_ASAP7_75t_SL g1006 ( .A(n_901), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_917), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_905), .B(n_902), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_847), .Y(n_1009) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_892), .Y(n_1010) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_896), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_829), .B(n_884), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_937), .A2(n_859), .B1(n_839), .B2(n_938), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_875), .Y(n_1014) );
INVxp67_ASAP7_75t_L g1015 ( .A(n_946), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1016 ( .A(n_836), .B(n_909), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_850), .B(n_863), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1018 ( .A(n_827), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_863), .B(n_858), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_830), .B(n_866), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_866), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_858), .B(n_867), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_867), .B(n_827), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_866), .Y(n_1024) );
OR2x2_ASAP7_75t_L g1025 ( .A(n_870), .B(n_904), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_935), .Y(n_1026) );
INVx2_ASAP7_75t_L g1027 ( .A(n_935), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_899), .B(n_912), .Y(n_1028) );
INVx2_ASAP7_75t_SL g1029 ( .A(n_944), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_859), .Y(n_1030) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_915), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_907), .B(n_911), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_887), .Y(n_1033) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_837), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_857), .B(n_860), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_852), .B(n_868), .Y(n_1036) );
HB1xp67_ASAP7_75t_L g1037 ( .A(n_855), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_913), .B(n_918), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_908), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_855), .B(n_861), .Y(n_1040) );
INVx2_ASAP7_75t_L g1041 ( .A(n_953), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_965), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_958), .B(n_846), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_990), .B(n_871), .Y(n_1044) );
NAND3xp33_ASAP7_75t_L g1045 ( .A(n_1013), .B(n_849), .C(n_864), .Y(n_1045) );
NAND3xp33_ASAP7_75t_L g1046 ( .A(n_1037), .B(n_851), .C(n_856), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_958), .B(n_828), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_954), .B(n_897), .Y(n_1048) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_982), .A2(n_831), .B1(n_885), .B2(n_929), .C(n_990), .Y(n_1049) );
OAI222xp33_ASAP7_75t_L g1050 ( .A1(n_993), .A2(n_1030), .B1(n_982), .B2(n_954), .C1(n_1019), .C2(n_1040), .Y(n_1050) );
HB1xp67_ASAP7_75t_L g1051 ( .A(n_951), .Y(n_1051) );
BUFx3_ASAP7_75t_L g1052 ( .A(n_986), .Y(n_1052) );
INVxp67_ASAP7_75t_L g1053 ( .A(n_1014), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_971), .B(n_1003), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_1030), .A2(n_1019), .B1(n_993), .B2(n_1040), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_978), .B(n_997), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_971), .B(n_1003), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_972), .B(n_973), .Y(n_1058) );
NOR3xp33_ASAP7_75t_L g1059 ( .A(n_1015), .B(n_995), .C(n_1029), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_972), .B(n_973), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_952), .B(n_962), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_952), .B(n_962), .Y(n_1062) );
HB1xp67_ASAP7_75t_L g1063 ( .A(n_994), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1064 ( .A(n_964), .B(n_979), .Y(n_1064) );
NAND2x1_ASAP7_75t_L g1065 ( .A(n_991), .B(n_1022), .Y(n_1065) );
OR2x2_ASAP7_75t_L g1066 ( .A(n_964), .B(n_979), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_950), .B(n_1008), .Y(n_1067) );
INVx5_ASAP7_75t_L g1068 ( .A(n_991), .Y(n_1068) );
OAI221xp5_ASAP7_75t_L g1069 ( .A1(n_1012), .A2(n_959), .B1(n_1033), .B2(n_1006), .C(n_1011), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_961), .B(n_947), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_970), .Y(n_1071) );
OAI221xp5_ASAP7_75t_L g1072 ( .A1(n_959), .A2(n_1006), .B1(n_1029), .B2(n_987), .C(n_957), .Y(n_1072) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_1010), .B(n_1007), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_970), .Y(n_1074) );
NAND2xp5_ASAP7_75t_SL g1075 ( .A(n_1036), .B(n_1022), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1008), .B(n_1010), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_957), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_975), .B(n_983), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1007), .B(n_1009), .Y(n_1079) );
INVx4_ASAP7_75t_L g1080 ( .A(n_988), .Y(n_1080) );
INVxp67_ASAP7_75t_L g1081 ( .A(n_989), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1016), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1083 ( .A(n_999), .B(n_1023), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_974), .B(n_949), .Y(n_1084) );
NAND2x1p5_ASAP7_75t_SL g1085 ( .A(n_1036), .B(n_1035), .Y(n_1085) );
OAI22xp33_ASAP7_75t_L g1086 ( .A1(n_1004), .A2(n_987), .B1(n_1017), .B2(n_1025), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_949), .B(n_1024), .Y(n_1087) );
NOR2xp33_ASAP7_75t_SL g1088 ( .A(n_1000), .B(n_995), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1016), .Y(n_1089) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_999), .B(n_1023), .Y(n_1090) );
OAI221xp5_ASAP7_75t_SL g1091 ( .A1(n_976), .A2(n_1025), .B1(n_1031), .B2(n_955), .C(n_1017), .Y(n_1091) );
NOR2xp33_ASAP7_75t_R g1092 ( .A(n_1000), .B(n_985), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_980), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_949), .B(n_1024), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_1020), .B(n_996), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g1096 ( .A1(n_1034), .A2(n_1028), .B1(n_1018), .B2(n_981), .C(n_967), .Y(n_1096) );
INVx1_ASAP7_75t_SL g1097 ( .A(n_1000), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1021), .B(n_996), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1021), .B(n_1001), .Y(n_1099) );
INVx4_ASAP7_75t_L g1100 ( .A(n_988), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1020), .B(n_1032), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_967), .A2(n_981), .B1(n_1028), .B2(n_1002), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1002), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1101), .B(n_1067), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_1064), .B(n_992), .Y(n_1105) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_1068), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g1107 ( .A(n_1063), .Y(n_1107) );
INVx2_ASAP7_75t_SL g1108 ( .A(n_1068), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1099), .Y(n_1109) );
NAND2x1_ASAP7_75t_L g1110 ( .A(n_1080), .B(n_960), .Y(n_1110) );
AOI31xp33_ASAP7_75t_SL g1111 ( .A1(n_1049), .A2(n_1038), .A3(n_966), .B(n_960), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1101), .B(n_966), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1067), .B(n_966), .Y(n_1113) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1041), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1099), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1098), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1117 ( .A1(n_1050), .A2(n_992), .B1(n_1026), .B2(n_1027), .C(n_968), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1041), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1054), .B(n_963), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1098), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1071), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1054), .B(n_960), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1061), .B(n_1005), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1074), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1057), .B(n_968), .Y(n_1125) );
NOR2xp67_ASAP7_75t_L g1126 ( .A(n_1068), .B(n_998), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1064), .B(n_1027), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1057), .B(n_1027), .Y(n_1128) );
NAND2xp5_ASAP7_75t_SL g1129 ( .A(n_1092), .B(n_1005), .Y(n_1129) );
AOI21xp5_ASAP7_75t_L g1130 ( .A1(n_1046), .A2(n_948), .B(n_992), .Y(n_1130) );
INVx4_ASAP7_75t_L g1131 ( .A(n_1068), .Y(n_1131) );
NOR2xp33_ASAP7_75t_R g1132 ( .A(n_1088), .B(n_1005), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1061), .B(n_984), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1084), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1062), .B(n_984), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1084), .Y(n_1136) );
INVx1_ASAP7_75t_SL g1137 ( .A(n_1092), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1076), .B(n_998), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1087), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1076), .B(n_998), .Y(n_1140) );
NOR2xp33_ASAP7_75t_L g1141 ( .A(n_1097), .B(n_988), .Y(n_1141) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_1051), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1062), .B(n_984), .Y(n_1143) );
NAND2x1_ASAP7_75t_L g1144 ( .A(n_1080), .B(n_956), .Y(n_1144) );
INVxp67_ASAP7_75t_L g1145 ( .A(n_1048), .Y(n_1145) );
NOR2x1_ASAP7_75t_L g1146 ( .A(n_1080), .B(n_956), .Y(n_1146) );
AND2x4_ASAP7_75t_L g1147 ( .A(n_1058), .B(n_1039), .Y(n_1147) );
INVx2_ASAP7_75t_SL g1148 ( .A(n_1068), .Y(n_1148) );
NOR2xp33_ASAP7_75t_SL g1149 ( .A(n_1100), .B(n_988), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1060), .B(n_1039), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1087), .Y(n_1151) );
NOR3xp33_ASAP7_75t_L g1152 ( .A(n_1069), .B(n_956), .C(n_977), .Y(n_1152) );
NAND3xp33_ASAP7_75t_L g1153 ( .A(n_1152), .B(n_1059), .C(n_1053), .Y(n_1153) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1114), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1105), .B(n_1066), .Y(n_1155) );
INVx2_ASAP7_75t_SL g1156 ( .A(n_1131), .Y(n_1156) );
BUFx3_ASAP7_75t_L g1157 ( .A(n_1131), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1104), .B(n_1083), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1121), .Y(n_1159) );
AOI221xp5_ASAP7_75t_SL g1160 ( .A1(n_1145), .A2(n_1055), .B1(n_1075), .B2(n_1048), .C(n_1086), .Y(n_1160) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1118), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1104), .B(n_1090), .Y(n_1162) );
OR2x2_ASAP7_75t_L g1163 ( .A(n_1105), .B(n_1066), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1134), .B(n_1042), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1121), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1124), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1124), .Y(n_1167) );
INVx1_ASAP7_75t_SL g1168 ( .A(n_1137), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1169 ( .A(n_1107), .Y(n_1169) );
AOI211xp5_ASAP7_75t_L g1170 ( .A1(n_1111), .A2(n_1072), .B(n_1091), .C(n_1075), .Y(n_1170) );
INVxp67_ASAP7_75t_L g1171 ( .A(n_1142), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1112), .B(n_1083), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1139), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1112), .B(n_1083), .Y(n_1174) );
AND2x4_ASAP7_75t_L g1175 ( .A(n_1116), .B(n_1094), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1139), .Y(n_1176) );
INVx1_ASAP7_75t_SL g1177 ( .A(n_1123), .Y(n_1177) );
INVxp67_ASAP7_75t_L g1178 ( .A(n_1141), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1151), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1138), .B(n_1090), .Y(n_1180) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1118), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1127), .B(n_1095), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1136), .B(n_1079), .Y(n_1183) );
INVxp67_ASAP7_75t_SL g1184 ( .A(n_1110), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1138), .B(n_1090), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1109), .B(n_1079), .Y(n_1186) );
AND2x4_ASAP7_75t_SL g1187 ( .A(n_1131), .B(n_1100), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1109), .B(n_1089), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1140), .B(n_1047), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1151), .Y(n_1190) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1115), .B(n_1082), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1140), .B(n_1047), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1115), .Y(n_1193) );
BUFx3_ASAP7_75t_L g1194 ( .A(n_1106), .Y(n_1194) );
HB1xp67_ASAP7_75t_L g1195 ( .A(n_1127), .Y(n_1195) );
AOI21xp33_ASAP7_75t_L g1196 ( .A1(n_1153), .A2(n_1044), .B(n_1056), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1189), .B(n_1113), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1155), .Y(n_1198) );
NAND2x1_ASAP7_75t_L g1199 ( .A(n_1156), .B(n_1106), .Y(n_1199) );
AOI21xp5_ASAP7_75t_L g1200 ( .A1(n_1187), .A2(n_1129), .B(n_1184), .Y(n_1200) );
INVx1_ASAP7_75t_SL g1201 ( .A(n_1168), .Y(n_1201) );
NAND2xp5_ASAP7_75t_SL g1202 ( .A(n_1157), .B(n_1132), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1155), .Y(n_1203) );
AOI21xp5_ASAP7_75t_L g1204 ( .A1(n_1187), .A2(n_1149), .B(n_1065), .Y(n_1204) );
INVx1_ASAP7_75t_SL g1205 ( .A(n_1168), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1158), .B(n_1119), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1163), .Y(n_1207) );
OAI322xp33_ASAP7_75t_L g1208 ( .A1(n_1171), .A2(n_1116), .A3(n_1120), .B1(n_1073), .B2(n_1143), .C1(n_1135), .C2(n_1133), .Y(n_1208) );
NOR4xp75_ASAP7_75t_L g1209 ( .A(n_1156), .B(n_1096), .C(n_1148), .D(n_1108), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1169), .B(n_1120), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1163), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1173), .Y(n_1212) );
AOI21xp33_ASAP7_75t_SL g1213 ( .A1(n_1153), .A2(n_1085), .B(n_1108), .Y(n_1213) );
INVxp67_ASAP7_75t_L g1214 ( .A(n_1194), .Y(n_1214) );
AOI22xp5_ASAP7_75t_L g1215 ( .A1(n_1160), .A2(n_1128), .B1(n_1125), .B2(n_1119), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1173), .Y(n_1216) );
AOI22xp5_ASAP7_75t_L g1217 ( .A1(n_1160), .A2(n_1128), .B1(n_1125), .B2(n_1122), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1176), .Y(n_1218) );
AOI22xp5_ASAP7_75t_L g1219 ( .A1(n_1170), .A2(n_1122), .B1(n_1147), .B2(n_1043), .Y(n_1219) );
AOI21xp33_ASAP7_75t_L g1220 ( .A1(n_1178), .A2(n_1081), .B(n_1073), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1189), .B(n_1113), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1193), .B(n_1150), .Y(n_1222) );
INVx2_ASAP7_75t_SL g1223 ( .A(n_1157), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1176), .Y(n_1224) );
NAND2xp5_ASAP7_75t_SL g1225 ( .A(n_1200), .B(n_1157), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1198), .B(n_1179), .Y(n_1226) );
OR2x2_ASAP7_75t_L g1227 ( .A(n_1203), .B(n_1195), .Y(n_1227) );
OAI21xp33_ASAP7_75t_L g1228 ( .A1(n_1219), .A2(n_1177), .B(n_1158), .Y(n_1228) );
AO22x2_ASAP7_75t_L g1229 ( .A1(n_1201), .A2(n_1190), .B1(n_1179), .B2(n_1193), .Y(n_1229) );
OAI21xp33_ASAP7_75t_L g1230 ( .A1(n_1213), .A2(n_1162), .B(n_1185), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1212), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1216), .Y(n_1232) );
INVx1_ASAP7_75t_SL g1233 ( .A(n_1223), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1197), .B(n_1162), .Y(n_1234) );
OAI21xp5_ASAP7_75t_L g1235 ( .A1(n_1204), .A2(n_1045), .B(n_1146), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1218), .Y(n_1236) );
NOR3xp33_ASAP7_75t_L g1237 ( .A(n_1196), .B(n_1190), .C(n_1103), .Y(n_1237) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1199), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1224), .Y(n_1239) );
AOI221xp5_ASAP7_75t_L g1240 ( .A1(n_1208), .A2(n_1085), .B1(n_1191), .B2(n_1188), .C(n_1164), .Y(n_1240) );
AOI22xp5_ASAP7_75t_L g1241 ( .A1(n_1215), .A2(n_1175), .B1(n_1183), .B2(n_1186), .Y(n_1241) );
AOI221xp5_ASAP7_75t_L g1242 ( .A1(n_1220), .A2(n_1192), .B1(n_1172), .B2(n_1174), .C(n_1175), .Y(n_1242) );
CKINVDCx14_ASAP7_75t_R g1243 ( .A(n_1197), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1221), .B(n_1192), .Y(n_1244) );
AOI221xp5_ASAP7_75t_L g1245 ( .A1(n_1240), .A2(n_1211), .B1(n_1207), .B2(n_1210), .C(n_1205), .Y(n_1245) );
AOI22xp33_ASAP7_75t_SL g1246 ( .A1(n_1243), .A2(n_1223), .B1(n_1187), .B2(n_1194), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1229), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1237), .B(n_1217), .Y(n_1248) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_1242), .A2(n_1222), .B1(n_1214), .B2(n_1221), .C(n_1206), .Y(n_1249) );
OAI21xp33_ASAP7_75t_L g1250 ( .A1(n_1230), .A2(n_1185), .B(n_1180), .Y(n_1250) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_1228), .A2(n_1175), .B1(n_1172), .B2(n_1174), .C(n_1166), .Y(n_1251) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1229), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1226), .Y(n_1253) );
O2A1O1Ixp33_ASAP7_75t_SL g1254 ( .A1(n_1225), .A2(n_1202), .B(n_1209), .C(n_1144), .Y(n_1254) );
AOI221xp5_ASAP7_75t_L g1255 ( .A1(n_1241), .A2(n_1159), .B1(n_1165), .B2(n_1166), .C(n_1167), .Y(n_1255) );
OAI21xp5_ASAP7_75t_L g1256 ( .A1(n_1235), .A2(n_1202), .B(n_1146), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1233), .B(n_1180), .Y(n_1257) );
NOR3xp33_ASAP7_75t_L g1258 ( .A(n_1245), .B(n_1235), .C(n_1238), .Y(n_1258) );
AOI21xp5_ASAP7_75t_L g1259 ( .A1(n_1254), .A2(n_1256), .B(n_1246), .Y(n_1259) );
AOI222xp33_ASAP7_75t_L g1260 ( .A1(n_1249), .A2(n_1233), .B1(n_1226), .B2(n_1236), .C1(n_1239), .C2(n_1231), .Y(n_1260) );
NOR3xp33_ASAP7_75t_L g1261 ( .A(n_1247), .B(n_1232), .C(n_1227), .Y(n_1261) );
NAND3xp33_ASAP7_75t_L g1262 ( .A(n_1252), .B(n_1117), .C(n_1167), .Y(n_1262) );
OAI211xp5_ASAP7_75t_SL g1263 ( .A1(n_1248), .A2(n_1102), .B(n_1078), .C(n_1093), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1253), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1255), .B(n_1244), .Y(n_1265) );
OAI21xp5_ASAP7_75t_L g1266 ( .A1(n_1259), .A2(n_1251), .B(n_1250), .Y(n_1266) );
NAND4xp75_ASAP7_75t_SL g1267 ( .A(n_1258), .B(n_1257), .C(n_1126), .D(n_1234), .Y(n_1267) );
OAI21xp5_ASAP7_75t_SL g1268 ( .A1(n_1260), .A2(n_1263), .B(n_1261), .Y(n_1268) );
NOR2xp33_ASAP7_75t_SL g1269 ( .A(n_1262), .B(n_1100), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_1265), .B(n_1264), .Y(n_1270) );
NOR3xp33_ASAP7_75t_L g1271 ( .A(n_1268), .B(n_1266), .C(n_1270), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1269), .B(n_1182), .Y(n_1272) );
NOR2x1_ASAP7_75t_L g1273 ( .A(n_1267), .B(n_1144), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1272), .Y(n_1274) );
XNOR2x1_ASAP7_75t_L g1275 ( .A(n_1273), .B(n_1052), .Y(n_1275) );
OAI22xp5_ASAP7_75t_L g1276 ( .A1(n_1271), .A2(n_1095), .B1(n_1147), .B2(n_1070), .Y(n_1276) );
AND2x4_ASAP7_75t_L g1277 ( .A(n_1274), .B(n_1147), .Y(n_1277) );
OAI22xp5_ASAP7_75t_SL g1278 ( .A1(n_1276), .A2(n_1275), .B1(n_988), .B2(n_1110), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1277), .Y(n_1279) );
OAI22x1_ASAP7_75t_SL g1280 ( .A1(n_1278), .A2(n_988), .B1(n_1077), .B2(n_956), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1279), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_1280), .A2(n_1181), .B1(n_1161), .B2(n_1154), .Y(n_1282) );
OAI21xp5_ASAP7_75t_SL g1283 ( .A1(n_1281), .A2(n_977), .B(n_969), .Y(n_1283) );
AOI21xp5_ASAP7_75t_L g1284 ( .A1(n_1283), .A2(n_1282), .B(n_1130), .Y(n_1284) );
endmodule