module fake_jpeg_30200_n_50 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_50);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_50;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g21 ( 
.A(n_6),
.B(n_17),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_21),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_37),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_5),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_35),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_1),
.B(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_4),
.B(n_10),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_32),
.C(n_8),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_45),
.C(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_38),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_39),
.C(n_46),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_11),
.C(n_12),
.Y(n_50)
);


endmodule