module fake_jpeg_11409_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_1),
.Y(n_6)
);

BUFx5_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx2_ASAP7_75t_SL g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_1),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx9p33_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_6),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_18),
.Y(n_19)
);

AO22x1_ASAP7_75t_L g16 ( 
.A1(n_8),
.A2(n_0),
.B1(n_3),
.B2(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_6),
.B1(n_16),
.B2(n_12),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_11),
.C(n_9),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_25),
.B(n_22),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_30),
.C(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

OAI221xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_9),
.B1(n_18),
.B2(n_16),
.C(n_10),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_17),
.C(n_7),
.Y(n_39)
);

AOI221xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_37),
.B1(n_17),
.B2(n_13),
.C(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);


endmodule