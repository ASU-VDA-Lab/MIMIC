module fake_netlist_6_2211_n_553 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_553);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_553;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_235;
wire n_536;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_516;
wire n_525;
wire n_491;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_456;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_546;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_162;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_27),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_51),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_4),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NOR2xp67_ASAP7_75t_L g165 ( 
.A(n_72),
.B(n_115),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_26),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_69),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_60),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_24),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_71),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_58),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_67),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_2),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_25),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_31),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_77),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_29),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_62),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_57),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_23),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_17),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_113),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_22),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_18),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_49),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_13),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_134),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_36),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_142),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_2),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_130),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_116),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_56),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_52),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_9),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_89),
.Y(n_217)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_110),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_150),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_127),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_149),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_59),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_92),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_10),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_75),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_11),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_133),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_139),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_74),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_147),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_99),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_98),
.Y(n_234)
);

BUFx8_ASAP7_75t_SL g235 ( 
.A(n_45),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_117),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_66),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_37),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_81),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_85),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_163),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_172),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_4),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

AND2x4_ASAP7_75t_L g251 ( 
.A(n_190),
.B(n_5),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_5),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_6),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_161),
.B(n_6),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_172),
.Y(n_258)
);

NOR2x1_ASAP7_75t_L g259 ( 
.A(n_165),
.B(n_12),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_182),
.B(n_7),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_192),
.B(n_7),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_159),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_172),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_201),
.B(n_8),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_160),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_208),
.B(n_8),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_164),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_172),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_166),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_9),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_197),
.B(n_14),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_167),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_10),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_197),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_11),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_15),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_217),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_186),
.B(n_189),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_253),
.A2(n_226),
.B1(n_176),
.B2(n_185),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_226),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_250),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_242),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_264),
.B1(n_260),
.B2(n_274),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_260),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_249),
.B(n_191),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_254),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_252),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_191),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

INVx4_ASAP7_75t_SL g295 ( 
.A(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_251),
.B(n_224),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_218),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_264),
.A2(n_274),
.B1(n_278),
.B2(n_265),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

AO22x2_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_224),
.B1(n_186),
.B2(n_189),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_259),
.B(n_241),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

AND3x2_ASAP7_75t_L g309 ( 
.A(n_256),
.B(n_240),
.C(n_239),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_243),
.B(n_168),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_169),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_248),
.B(n_276),
.C(n_271),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_245),
.B(n_170),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_245),
.B(n_173),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_174),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_175),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_171),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_L g319 ( 
.A1(n_246),
.A2(n_162),
.B1(n_187),
.B2(n_238),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_247),
.B(n_177),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_272),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_282),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_183),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_257),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_258),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_263),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_298),
.B(n_268),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_284),
.Y(n_329)
);

AND2x6_ASAP7_75t_SL g330 ( 
.A(n_311),
.B(n_246),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_195),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_196),
.B1(n_219),
.B2(n_200),
.Y(n_332)
);

AOI22x1_ASAP7_75t_L g333 ( 
.A1(n_304),
.A2(n_211),
.B1(n_180),
.B2(n_234),
.Y(n_333)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_310),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_203),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_286),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_319),
.B(n_206),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_281),
.B(n_228),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_306),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_300),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_178),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_285),
.A2(n_244),
.B1(n_213),
.B2(n_209),
.Y(n_348)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_SL g350 ( 
.A1(n_317),
.A2(n_214),
.B(n_184),
.C(n_231),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_283),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_305),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_312),
.B(n_229),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_232),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_287),
.B(n_181),
.Y(n_356)
);

AND2x6_ASAP7_75t_SL g357 ( 
.A(n_287),
.B(n_188),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_284),
.B(n_193),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_314),
.B(n_272),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_315),
.B(n_316),
.Y(n_360)
);

NOR2x2_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_194),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_321),
.B(n_217),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_320),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g366 ( 
.A(n_321),
.B(n_272),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_315),
.B(n_198),
.Y(n_367)
);

NAND3xp33_ASAP7_75t_SL g368 ( 
.A(n_332),
.B(n_339),
.C(n_337),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_329),
.B(n_316),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_322),
.B(n_321),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_313),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_348),
.A2(n_356),
.B1(n_365),
.B2(n_353),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_344),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_326),
.A2(n_327),
.B(n_325),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_324),
.B(n_321),
.Y(n_377)
);

AOI21x1_ASAP7_75t_L g378 ( 
.A1(n_359),
.A2(n_220),
.B(n_202),
.Y(n_378)
);

BUFx12f_ASAP7_75t_L g379 ( 
.A(n_357),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_358),
.A2(n_221),
.B1(n_204),
.B2(n_205),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_367),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_295),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_342),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_295),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

O2A1O1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_331),
.A2(n_230),
.B(n_222),
.C(n_215),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_347),
.Y(n_388)
);

OAI22x1_ASAP7_75t_L g389 ( 
.A1(n_333),
.A2(n_199),
.B1(n_307),
.B2(n_309),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_295),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_323),
.B(n_16),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_340),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_392)
);

AOI21x1_ASAP7_75t_L g393 ( 
.A1(n_354),
.A2(n_364),
.B(n_363),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_335),
.A2(n_156),
.B1(n_30),
.B2(n_32),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_346),
.B(n_28),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_334),
.B(n_33),
.Y(n_396)
);

OR2x6_ASAP7_75t_L g397 ( 
.A(n_346),
.B(n_34),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_328),
.B(n_35),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_362),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_336),
.B(n_38),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_338),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_366),
.A2(n_39),
.B(n_40),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

AO22x1_ASAP7_75t_L g406 ( 
.A1(n_361),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_406)
);

BUFx4f_ASAP7_75t_L g407 ( 
.A(n_351),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_SL g408 ( 
.A(n_345),
.B(n_48),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_350),
.A2(n_345),
.B(n_349),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_375),
.A2(n_345),
.B(n_349),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_383),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_349),
.Y(n_412)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_393),
.A2(n_153),
.B(n_53),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_405),
.Y(n_414)
);

AO31x2_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_50),
.A3(n_54),
.B(n_55),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_381),
.A2(n_63),
.B(n_64),
.Y(n_416)
);

OR2x6_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_70),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_382),
.A2(n_152),
.B(n_78),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

O2A1O1Ixp5_ASAP7_75t_L g420 ( 
.A1(n_371),
.A2(n_378),
.B(n_391),
.C(n_377),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_372),
.A2(n_73),
.B1(n_79),
.B2(n_80),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_374),
.Y(n_422)
);

NAND2x1_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_82),
.Y(n_423)
);

AO31x2_ASAP7_75t_L g424 ( 
.A1(n_380),
.A2(n_389),
.A3(n_394),
.B(n_401),
.Y(n_424)
);

A2O1A1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_372),
.A2(n_400),
.B(n_396),
.C(n_387),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_385),
.B(n_83),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_368),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_88),
.B(n_90),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_394),
.B(n_91),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_386),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_392),
.A2(n_93),
.B(n_95),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_409),
.A2(n_96),
.B(n_97),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_386),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_403),
.Y(n_436)
);

AO31x2_ASAP7_75t_L g437 ( 
.A1(n_404),
.A2(n_100),
.A3(n_102),
.B(n_103),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

O2A1O1Ixp33_ASAP7_75t_L g439 ( 
.A1(n_395),
.A2(n_107),
.B(n_109),
.C(n_112),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_384),
.A2(n_114),
.B(n_119),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_411),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_425),
.A2(n_407),
.B1(n_390),
.B2(n_397),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_438),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_412),
.B(n_407),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_406),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_422),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_397),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_430),
.A2(n_417),
.B1(n_421),
.B2(n_426),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_414),
.Y(n_450)
);

O2A1O1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_430),
.A2(n_370),
.B(n_376),
.C(n_373),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_413),
.A2(n_408),
.B(n_121),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_414),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_420),
.A2(n_120),
.B(n_122),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_421),
.A2(n_379),
.B1(n_129),
.B2(n_136),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_151),
.Y(n_456)
);

BUFx12f_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

AOI221xp5_ASAP7_75t_L g458 ( 
.A1(n_432),
.A2(n_123),
.B1(n_137),
.B2(n_138),
.C(n_141),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_433),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_410),
.A2(n_143),
.B(n_145),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_417),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_441),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_431),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

AO21x2_ASAP7_75t_L g465 ( 
.A1(n_454),
.A2(n_410),
.B(n_432),
.Y(n_465)
);

OAI221xp5_ASAP7_75t_SL g466 ( 
.A1(n_455),
.A2(n_427),
.B1(n_439),
.B2(n_416),
.C(n_440),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_447),
.Y(n_467)
);

AO21x2_ASAP7_75t_L g468 ( 
.A1(n_459),
.A2(n_416),
.B(n_440),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

OA21x2_ASAP7_75t_L g470 ( 
.A1(n_459),
.A2(n_418),
.B(n_436),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_460),
.A2(n_435),
.B(n_424),
.Y(n_471)
);

AOI221xp5_ASAP7_75t_L g472 ( 
.A1(n_449),
.A2(n_458),
.B1(n_443),
.B2(n_451),
.C(n_461),
.Y(n_472)
);

NAND2x1_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_429),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_462),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_444),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_445),
.B(n_415),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_457),
.Y(n_477)
);

OA21x2_ASAP7_75t_L g478 ( 
.A1(n_452),
.A2(n_415),
.B(n_437),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_444),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_453),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_481),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_464),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_481),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_448),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_472),
.A2(n_457),
.B1(n_448),
.B2(n_456),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_462),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_480),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_463),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_480),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_475),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_476),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_469),
.B(n_446),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_479),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_444),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_456),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_423),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_483),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_493),
.B(n_471),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_482),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g504 ( 
.A(n_493),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_482),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_492),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_484),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_484),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_471),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_415),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_471),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_437),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_478),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_488),
.B(n_437),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_491),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_485),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_465),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_499),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_515),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_498),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_501),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_503),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_498),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_503),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_508),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_511),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_521),
.B(n_510),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_504),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_524),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_529),
.B(n_520),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_527),
.A2(n_487),
.B(n_517),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_528),
.Y(n_532)
);

AOI221xp5_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_526),
.B1(n_517),
.B2(n_466),
.C(n_477),
.Y(n_533)
);

OAI211xp5_ASAP7_75t_SL g534 ( 
.A1(n_530),
.A2(n_509),
.B(n_518),
.C(n_496),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_L g535 ( 
.A1(n_532),
.A2(n_520),
.B1(n_509),
.B2(n_502),
.Y(n_535)
);

OA211x2_ASAP7_75t_L g536 ( 
.A1(n_533),
.A2(n_473),
.B(n_477),
.C(n_504),
.Y(n_536)
);

AOI211x1_ASAP7_75t_SL g537 ( 
.A1(n_534),
.A2(n_525),
.B(n_522),
.C(n_508),
.Y(n_537)
);

NOR4xp75_ASAP7_75t_L g538 ( 
.A(n_535),
.B(n_489),
.C(n_514),
.D(n_494),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_536),
.A2(n_498),
.B1(n_491),
.B2(n_500),
.Y(n_539)
);

NAND4xp25_ASAP7_75t_L g540 ( 
.A(n_537),
.B(n_507),
.C(n_505),
.D(n_525),
.Y(n_540)
);

AOI211xp5_ASAP7_75t_L g541 ( 
.A1(n_538),
.A2(n_522),
.B(n_516),
.C(n_452),
.Y(n_541)
);

OAI221xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_429),
.B1(n_478),
.B2(n_485),
.C(n_495),
.Y(n_542)
);

NOR3xp33_ASAP7_75t_L g543 ( 
.A(n_540),
.B(n_495),
.C(n_499),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_542),
.B(n_539),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_543),
.Y(n_545)
);

AO21x2_ASAP7_75t_L g546 ( 
.A1(n_543),
.A2(n_468),
.B(n_465),
.Y(n_546)
);

XNOR2x1_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_146),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_545),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_547),
.A2(n_545),
.B1(n_548),
.B2(n_546),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_465),
.B(n_468),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_550),
.A2(n_470),
.B(n_478),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_148),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_552),
.A2(n_478),
.B1(n_468),
.B2(n_470),
.Y(n_553)
);


endmodule