module fake_jpeg_16925_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_21),
.Y(n_44)
);

HAxp5_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_23),
.CON(n_66),
.SN(n_66)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_50),
.B(n_54),
.Y(n_103)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_32),
.B1(n_21),
.B2(n_34),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_53),
.B1(n_57),
.B2(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_32),
.B1(n_21),
.B2(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_16),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_62),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_28),
.B1(n_26),
.B2(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_23),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_64),
.Y(n_79)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_40),
.B(n_42),
.C(n_25),
.Y(n_101)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_38),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_76),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_56),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_78),
.Y(n_123)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_82),
.B(n_96),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_30),
.B(n_18),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_35),
.B1(n_38),
.B2(n_37),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_92),
.B1(n_97),
.B2(n_31),
.Y(n_107)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_87),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_18),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_98),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_27),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_94),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_29),
.B1(n_38),
.B2(n_17),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_64),
.Y(n_96)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_40),
.B1(n_42),
.B2(n_31),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_22),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_104),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_46),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_102),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_25),
.B(n_20),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_60),
.B(n_22),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

AOI22x1_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_25),
.B1(n_31),
.B2(n_17),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_128),
.B(n_94),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_107),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_104),
.A2(n_42),
.B1(n_31),
.B2(n_20),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_111),
.B1(n_127),
.B2(n_81),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_120),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_81),
.B(n_71),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_71),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_73),
.A2(n_20),
.B1(n_25),
.B2(n_27),
.Y(n_127)
);

NAND2x1_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_27),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_142),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_137),
.A2(n_152),
.B(n_112),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_100),
.B1(n_91),
.B2(n_86),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_138),
.A2(n_149),
.B1(n_150),
.B2(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_75),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_82),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_72),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_147),
.B(n_157),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_79),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_106),
.A2(n_84),
.B1(n_76),
.B2(n_95),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_106),
.A2(n_97),
.B1(n_93),
.B2(n_101),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_164),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_97),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_130),
.B(n_19),
.Y(n_193)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_129),
.B1(n_115),
.B2(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_103),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_158),
.B(n_162),
.Y(n_173)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_88),
.C(n_78),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_153),
.C(n_137),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_77),
.B1(n_8),
.B2(n_14),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_132),
.B1(n_116),
.B2(n_5),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_6),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_117),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_124),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_174),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_185),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_111),
.B1(n_114),
.B2(n_121),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_145),
.B1(n_142),
.B2(n_151),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_192),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_144),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_183),
.C(n_190),
.Y(n_204)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_114),
.B(n_113),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_181),
.B(n_196),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_130),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_184),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_116),
.A3(n_132),
.B1(n_109),
.B2(n_126),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_124),
.C(n_126),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_194),
.B(n_197),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_19),
.B(n_120),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_223),
.B1(n_188),
.B2(n_182),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_170),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_209),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_152),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_206),
.C(n_204),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_150),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_139),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_211),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_220),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_139),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_149),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_120),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_195),
.A2(n_118),
.B1(n_88),
.B2(n_19),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_19),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_224),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_187),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_232),
.C(n_234),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_232),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_187),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_193),
.B(n_194),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_233),
.A2(n_241),
.B(n_217),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_172),
.C(n_190),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_242),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_207),
.B1(n_203),
.B2(n_212),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_180),
.C(n_175),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_243),
.C(n_244),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_166),
.B(n_185),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_180),
.C(n_166),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_196),
.C(n_173),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_174),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.C(n_0),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_88),
.C(n_19),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_212),
.C(n_199),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_255),
.B(n_244),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_201),
.B1(n_211),
.B2(n_221),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_253),
.B1(n_264),
.B2(n_262),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_256),
.C(n_230),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

AOI221xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_202),
.B1(n_213),
.B2(n_223),
.C(n_210),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_214),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_263),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_246),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_217),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_260),
.B(n_225),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_229),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_261),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_236),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_250),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_252),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_261),
.B(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_273),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_0),
.Y(n_289)
);

XNOR2x2_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_248),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_258),
.B(n_249),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_272),
.C(n_278),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_234),
.Y(n_278)
);

BUFx4f_ASAP7_75t_SL g280 ( 
.A(n_277),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_280),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_285),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_284),
.A2(n_7),
.B1(n_11),
.B2(n_3),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_264),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_258),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_287),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_249),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_290),
.C(n_5),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_276),
.C(n_274),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_270),
.B1(n_275),
.B2(n_3),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_296),
.A2(n_10),
.B1(n_13),
.B2(n_4),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_298),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_13),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_280),
.C(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_295),
.C(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_289),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_306),
.A3(n_7),
.B1(n_11),
.B2(n_13),
.C1(n_1),
.C2(n_0),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_296),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_284),
.B1(n_10),
.B2(n_4),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_297),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_309),
.A2(n_310),
.B1(n_305),
.B2(n_303),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_311),
.B(n_302),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_314),
.Y(n_315)
);


endmodule