module fake_netlist_1_798_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
NAND2xp5_ASAP7_75t_L g4 ( .A(n_2), .B(n_1), .Y(n_4) );
NAND2xp5_ASAP7_75t_SL g5 ( .A(n_1), .B(n_0), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
OAI22xp5_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_3), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_7), .B(n_5), .Y(n_9) );
OAI22xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_8), .B(n_2), .Y(n_11) );
OAI21xp33_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_8), .B(n_1), .Y(n_12) );
OAI211xp5_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_0), .B(n_2), .C(n_10), .Y(n_13) );
NOR2x1p5_ASAP7_75t_L g14 ( .A(n_13), .B(n_0), .Y(n_14) );
OR2x2_ASAP7_75t_L g15 ( .A(n_12), .B(n_2), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_14), .B(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_16), .Y(n_18) );
endmodule