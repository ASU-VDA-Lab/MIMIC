module fake_jpeg_8904_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_37),
.Y(n_46)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_27),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_22),
.B1(n_19),
.B2(n_17),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_48),
.B1(n_60),
.B2(n_27),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_22),
.B1(n_24),
.B2(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_17),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_22),
.B1(n_19),
.B2(n_31),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_89),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_27),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_80),
.C(n_37),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_41),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_40),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_24),
.B1(n_16),
.B2(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_40),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_67),
.Y(n_112)
);

NOR2x1_ASAP7_75t_R g91 ( 
.A(n_62),
.B(n_24),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_24),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_39),
.B1(n_57),
.B2(n_53),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_106),
.B1(n_111),
.B2(n_69),
.Y(n_133)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_102),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_80),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_98),
.B(n_100),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_68),
.Y(n_120)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_51),
.B1(n_45),
.B2(n_38),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_109),
.B1(n_26),
.B2(n_69),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_39),
.B1(n_51),
.B2(n_45),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_107),
.Y(n_121)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_108),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_37),
.B1(n_38),
.B2(n_16),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_65),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_71),
.C(n_69),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_68),
.A2(n_16),
.B1(n_31),
.B2(n_32),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_20),
.B(n_21),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_81),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_20),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_26),
.B1(n_33),
.B2(n_30),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_135),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_126),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_143),
.C(n_84),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_97),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_80),
.B(n_76),
.C(n_30),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_76),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_131),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_76),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_136),
.B(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_80),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_139),
.B1(n_94),
.B2(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_71),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_139),
.B(n_142),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_79),
.C(n_90),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_0),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_146),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_174),
.B1(n_177),
.B2(n_144),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_147),
.A2(n_94),
.B1(n_114),
.B2(n_93),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_152),
.B1(n_163),
.B2(n_170),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_111),
.B1(n_103),
.B2(n_77),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_154),
.C(n_162),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_118),
.C(n_109),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_155),
.B(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2x1_ASAP7_75t_R g161 ( 
.A(n_126),
.B(n_32),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g203 ( 
.A1(n_161),
.A2(n_28),
.B1(n_25),
.B2(n_18),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_108),
.B1(n_102),
.B2(n_107),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_85),
.Y(n_164)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_168),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_85),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_84),
.B1(n_75),
.B2(n_70),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_99),
.C(n_70),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_173),
.C(n_120),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_32),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_128),
.A2(n_33),
.B1(n_99),
.B2(n_13),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_137),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_32),
.B1(n_28),
.B2(n_25),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_176),
.A2(n_25),
.B1(n_18),
.B2(n_32),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_28),
.B1(n_25),
.B2(n_18),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_138),
.B1(n_129),
.B2(n_133),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_149),
.B1(n_156),
.B2(n_152),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_197),
.C(n_200),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_129),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_191),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_160),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_193),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_20),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

AOI22x1_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_130),
.B1(n_145),
.B2(n_120),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_176),
.B1(n_28),
.B2(n_25),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_130),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_158),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_199),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_145),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_172),
.C(n_156),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_150),
.Y(n_202)
);

HB1xp67_ASAP7_75t_SL g227 ( 
.A(n_202),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_165),
.B(n_157),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_154),
.C(n_173),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_207),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_157),
.C(n_151),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_214),
.C(n_224),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_218),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_220),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_28),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_21),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_11),
.B(n_15),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_203),
.B1(n_183),
.B2(n_189),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_179),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_18),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_180),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_20),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_189),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_200),
.C(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_239),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_237),
.A2(n_0),
.B(n_1),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_178),
.C(n_183),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_198),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_187),
.B1(n_178),
.B2(n_199),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_212),
.B1(n_215),
.B2(n_211),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_209),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_244),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_9),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_0),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_217),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_21),
.C(n_20),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_208),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_252),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_219),
.B1(n_227),
.B2(n_220),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_258),
.B1(n_236),
.B2(n_229),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_215),
.Y(n_255)
);

OAI321xp33_ASAP7_75t_L g257 ( 
.A1(n_241),
.A2(n_215),
.A3(n_242),
.B1(n_244),
.B2(n_233),
.C(n_230),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_4),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_207),
.B1(n_205),
.B2(n_224),
.Y(n_258)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_2),
.B(n_3),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_240),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_262),
.A2(n_265),
.B(n_236),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_20),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_229),
.C(n_235),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_20),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_266),
.B(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_231),
.B(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_231),
.C(n_248),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_271),
.B(n_5),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_278),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_9),
.C(n_11),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_259),
.B(n_253),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_275),
.A2(n_252),
.B(n_261),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_4),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_12),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_286),
.B(n_274),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_276),
.Y(n_297)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_287),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g286 ( 
.A(n_271),
.B(n_6),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_279),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_280),
.A2(n_277),
.B1(n_273),
.B2(n_267),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_294),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_284),
.B(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_296),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_266),
.B(n_278),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_297),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_287),
.A2(n_272),
.B(n_274),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_14),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_299),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_12),
.C(n_13),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_303),
.B(n_14),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_299),
.B(n_15),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_308),
.B(n_304),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_307),
.C(n_305),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_14),
.B(n_21),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_311),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_21),
.B(n_301),
.Y(n_313)
);


endmodule