module fake_jpeg_20733_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

HAxp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_26),
.CON(n_39),
.SN(n_39)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_16),
.B1(n_23),
.B2(n_32),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_19),
.Y(n_50)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_19),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_19),
.B(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_32),
.B1(n_27),
.B2(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_55),
.B1(n_36),
.B2(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_32),
.B1(n_23),
.B2(n_25),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_36),
.B1(n_34),
.B2(n_41),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_63),
.Y(n_88)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_64),
.B(n_69),
.Y(n_101)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_65),
.A2(n_40),
.B1(n_37),
.B2(n_33),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_53),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_72),
.B1(n_77),
.B2(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_17),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_79),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_36),
.B1(n_38),
.B2(n_24),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_73),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_29),
.B(n_24),
.C(n_26),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_22),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_19),
.Y(n_100)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_38),
.B1(n_37),
.B2(n_42),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_40),
.B(n_35),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_40),
.C(n_35),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_78),
.Y(n_83)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_51),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_92),
.C(n_90),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_55),
.B1(n_54),
.B2(n_52),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_71),
.B1(n_63),
.B2(n_61),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_102),
.B1(n_105),
.B2(n_67),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_90),
.B(n_82),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_79),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_76),
.B1(n_57),
.B2(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_110),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_115),
.B1(n_119),
.B2(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_62),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_59),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_120),
.Y(n_131)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_65),
.B1(n_33),
.B2(n_40),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_89),
.B1(n_98),
.B2(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_19),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_97),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_66),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_26),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_101),
.C(n_93),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_83),
.B1(n_90),
.B2(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_104),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_138),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_132),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_94),
.B(n_97),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_139),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_144),
.B1(n_145),
.B2(n_3),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_26),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_31),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_146),
.A2(n_125),
.B1(n_119),
.B2(n_117),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_155),
.B1(n_158),
.B2(n_133),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_108),
.B(n_113),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_144),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_133),
.A2(n_120),
.B1(n_106),
.B2(n_114),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_107),
.B1(n_113),
.B2(n_118),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_130),
.A2(n_126),
.B1(n_112),
.B2(n_25),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_126),
.B1(n_112),
.B2(n_25),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_160),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_30),
.A3(n_10),
.B1(n_11),
.B2(n_15),
.C1(n_13),
.C2(n_12),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_168),
.Y(n_181)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_135),
.B(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_167),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_127),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_157),
.C(n_147),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_169),
.B1(n_172),
.B2(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_161),
.B(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_136),
.B1(n_145),
.B2(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_142),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_129),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_156),
.C(n_157),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_175),
.B(n_178),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_180),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_149),
.C(n_154),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_164),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_179),
.B(n_169),
.CI(n_166),
.CON(n_182),
.SN(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_158),
.C(n_28),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_182),
.B(n_184),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_181),
.B(n_172),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_4),
.B(n_5),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_5),
.C(n_6),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_4),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_9),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_192),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_SL g190 ( 
.A1(n_183),
.A2(n_175),
.B(n_7),
.C(n_8),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_188),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_6),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_193),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_195),
.B(n_197),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_185),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_194),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_199),
.B(n_196),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.C(n_190),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_9),
.Y(n_204)
);


endmodule