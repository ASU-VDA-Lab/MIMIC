module real_jpeg_29217_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g62 ( 
.A(n_0),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_22),
.B1(n_25),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_4),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_4),
.A2(n_40),
.B1(n_60),
.B2(n_61),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_42),
.B1(n_44),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_76)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_9),
.A2(n_22),
.B1(n_25),
.B2(n_29),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_9),
.A2(n_29),
.B1(n_42),
.B2(n_44),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_9),
.A2(n_29),
.B1(n_60),
.B2(n_61),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_10),
.A2(n_22),
.B1(n_25),
.B2(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_22),
.B1(n_25),
.B2(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_11),
.A2(n_32),
.B1(n_42),
.B2(n_44),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g123 ( 
.A1(n_11),
.A2(n_22),
.B(n_24),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_11),
.A2(n_32),
.B1(n_60),
.B2(n_61),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_11),
.B(n_21),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_11),
.A2(n_42),
.B(n_164),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_11),
.A2(n_57),
.B(n_61),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_11),
.B(n_41),
.Y(n_187)
);

XNOR2x2_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_111),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_109),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_92),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_15),
.B(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_73),
.B1(n_74),
.B2(n_91),
.Y(n_15)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_65),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_35),
.B2(n_36),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_18),
.A2(n_19),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_18),
.A2(n_19),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_18),
.B(n_223),
.C(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_19),
.B(n_108),
.C(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_26),
.B(n_30),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_33),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_21),
.A2(n_31),
.B1(n_33),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

INVx5_ASAP7_75t_SL g25 ( 
.A(n_22),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_22),
.A2(n_32),
.B(n_43),
.C(n_163),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_23),
.A2(n_28),
.B(n_32),
.C(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_31),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_32),
.A2(n_42),
.B(n_58),
.C(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_32),
.B(n_102),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_32),
.B(n_59),
.Y(n_199)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_51),
.B2(n_52),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B(n_45),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_41),
.B(n_48),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_44),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_46),
.A2(n_70),
.B(n_72),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_50),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_63),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_54),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_59),
.B1(n_63),
.B2(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_55),
.A2(n_59),
.B1(n_86),
.B2(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_67),
.B(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_60),
.B(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_66),
.B(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_68),
.A2(n_105),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_68),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_68),
.B(n_151),
.C(n_154),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_68),
.A2(n_119),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_71),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_82),
.B(n_87),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_87),
.B1(n_88),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_75),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_75),
.A2(n_83),
.B1(n_95),
.B2(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_79),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_78),
.B(n_143),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_102),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_83),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_85),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.C(n_97),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_93),
.B(n_96),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_97),
.A2(n_98),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.C(n_107),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_99),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_100),
.A2(n_103),
.B1(n_178),
.B2(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_100),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_102),
.B(n_141),
.Y(n_140)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_103),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_103),
.A2(n_178),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_103),
.B(n_124),
.C(n_188),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_103),
.B(n_169),
.C(n_177),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_105),
.B(n_119),
.C(n_120),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_118),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_108),
.B1(n_130),
.B2(n_131),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_136),
.C(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_107),
.A2(n_108),
.B1(n_135),
.B2(n_136),
.Y(n_206)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_243),
.B(n_248),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_231),
.B(n_242),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_156),
.B(n_215),
.C(n_230),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_144),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_115),
.B(n_144),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_127),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_116),
.B(n_128),
.C(n_134),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_124),
.A2(n_149),
.B1(n_186),
.B2(n_189),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_124),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_124),
.B(n_199),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_141),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_135),
.A2(n_136),
.B1(n_183),
.B2(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_135),
.B(n_140),
.Y(n_223)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_150),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_145),
.B(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_148),
.B(n_150),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_154),
.B1(n_155),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_151),
.B(n_196),
.Y(n_195)
);

INVx5_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_214),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_209),
.B(n_213),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_179),
.B(n_208),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_168),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_167),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_172),
.B(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_176),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_203),
.B(n_207),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_190),
.B(n_202),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_185),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_183),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_186),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_194),
.B(n_201),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_198),
.B(n_200),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_205),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_217),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_228),
.B2(n_229),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_222),
.C(n_229),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_228),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_232),
.B(n_233),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_241),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_239),
.C(n_241),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_245),
.Y(n_248)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);


endmodule