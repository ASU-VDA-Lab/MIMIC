module fake_jpeg_15670_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_14),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_18),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_63),
.B1(n_30),
.B2(n_22),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_62),
.B1(n_22),
.B2(n_64),
.Y(n_100)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_59),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_30),
.B1(n_34),
.B2(n_20),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_20),
.B1(n_27),
.B2(n_18),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_34),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_31),
.B(n_20),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_20),
.B(n_28),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_28),
.C(n_42),
.Y(n_102)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_79),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_78),
.A2(n_104),
.B1(n_72),
.B2(n_68),
.Y(n_114)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_90),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_17),
.B1(n_29),
.B2(n_16),
.Y(n_119)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_47),
.B1(n_36),
.B2(n_45),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_98),
.B1(n_105),
.B2(n_59),
.Y(n_110)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_21),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_19),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_69),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_97),
.Y(n_134)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_99),
.B(n_106),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_72),
.B1(n_44),
.B2(n_38),
.Y(n_118)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_46),
.C(n_44),
.Y(n_121)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_46),
.B1(n_44),
.B2(n_38),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_110),
.A2(n_129),
.B1(n_131),
.B2(n_133),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_54),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_121),
.C(n_37),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_21),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_115),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_88),
.B1(n_104),
.B2(n_87),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_125),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_87),
.B1(n_93),
.B2(n_33),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_93),
.B1(n_1),
.B2(n_2),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_86),
.B(n_99),
.C(n_84),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_73),
.B1(n_51),
.B2(n_17),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_81),
.B(n_17),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_73),
.B1(n_29),
.B2(n_17),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_75),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_85),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_82),
.A2(n_73),
.B1(n_29),
.B2(n_11),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_28),
.B(n_26),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_103),
.B(n_97),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_95),
.B1(n_101),
.B2(n_88),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_150),
.B1(n_163),
.B2(n_133),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_103),
.B(n_83),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_138),
.A2(n_142),
.B(n_126),
.Y(n_200)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_144),
.B(n_146),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_75),
.B(n_96),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_0),
.B(n_1),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_105),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_162),
.C(n_120),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_0),
.B(n_1),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_79),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_85),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_153),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_28),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_74),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_117),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_37),
.B(n_28),
.C(n_88),
.D(n_89),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_157),
.A2(n_118),
.B1(n_109),
.B2(n_131),
.Y(n_191)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_57),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_57),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_168),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_121),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_177),
.A2(n_180),
.B(n_200),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_136),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_136),
.B1(n_161),
.B2(n_153),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_182),
.B(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_143),
.B(n_113),
.Y(n_183)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_192),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_119),
.B1(n_120),
.B2(n_109),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_191),
.B1(n_163),
.B2(n_154),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_193),
.C(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_124),
.C(n_126),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_143),
.B(n_108),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_198),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_158),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_124),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_109),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_129),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_33),
.Y(n_227)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_144),
.A2(n_33),
.B1(n_32),
.B2(n_29),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_203),
.A2(n_164),
.B1(n_112),
.B2(n_33),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_145),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_204),
.B(n_207),
.C(n_211),
.Y(n_258)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_146),
.B1(n_147),
.B2(n_136),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_205),
.A2(n_216),
.B1(n_224),
.B2(n_228),
.Y(n_249)
);

AOI222xp33_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_147),
.B1(n_141),
.B2(n_137),
.C1(n_138),
.C2(n_136),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_225),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_142),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_172),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_226),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_196),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_220),
.Y(n_237)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_230),
.B1(n_203),
.B2(n_195),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_137),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_166),
.B(n_155),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_176),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_32),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_156),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_172),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_173),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_169),
.A2(n_0),
.B(n_3),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_232),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_180),
.B1(n_192),
.B2(n_188),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_233),
.A2(n_240),
.B1(n_245),
.B2(n_224),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_225),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_234),
.B(n_250),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_200),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_243),
.C(n_211),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_174),
.B1(n_170),
.B2(n_194),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_186),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_174),
.B1(n_171),
.B2(n_190),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_182),
.Y(n_246)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVxp67_ASAP7_75t_SL g251 ( 
.A(n_228),
.Y(n_251)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_208),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_252),
.A2(n_197),
.B1(n_178),
.B2(n_173),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_202),
.B1(n_185),
.B2(n_5),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_254),
.A2(n_210),
.B1(n_212),
.B2(n_178),
.Y(n_260)
);

FAx1_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_169),
.CI(n_179),
.CON(n_255),
.SN(n_255)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_32),
.B(n_26),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_175),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_187),
.B(n_183),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_255),
.A2(n_212),
.B1(n_229),
.B2(n_227),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_259),
.A2(n_272),
.B1(n_273),
.B2(n_240),
.Y(n_292)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_217),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_265),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_220),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_267),
.C(n_270),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_222),
.C(n_187),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_275),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_222),
.C(n_215),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_171),
.C(n_230),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_278),
.C(n_237),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_232),
.B1(n_191),
.B2(n_169),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_32),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_277),
.B(n_233),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_26),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_282),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_252),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_288),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_241),
.B1(n_257),
.B2(n_244),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_238),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_293),
.C(n_262),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_276),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_264),
.B(n_236),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_295),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_275),
.A2(n_245),
.B1(n_242),
.B2(n_235),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_272),
.B1(n_278),
.B2(n_5),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_9),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_277),
.B(n_259),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_297),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_308),
.Y(n_314)
);

AO221x1_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_273),
.B1(n_274),
.B2(n_282),
.C(n_292),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_SL g312 ( 
.A(n_300),
.B(n_3),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_283),
.C(n_291),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_304),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_289),
.A2(n_270),
.B(n_261),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_303),
.A2(n_10),
.B(n_4),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_285),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_265),
.C(n_271),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_306),
.B(n_307),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_293),
.C(n_266),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_287),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_280),
.B1(n_287),
.B2(n_11),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_316),
.B1(n_7),
.B2(n_8),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_3),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_7),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_263),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_320),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_13),
.B(n_12),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_319),
.B(n_6),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_10),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_324),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_301),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_328),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_330),
.B(n_8),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_8),
.B(n_26),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_314),
.C(n_322),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_321),
.A2(n_317),
.B(n_311),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_335),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_327),
.B(n_323),
.Y(n_337)
);

AOI21x1_ASAP7_75t_L g340 ( 
.A1(n_337),
.A2(n_339),
.B(n_332),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_331),
.C(n_338),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_334),
.Y(n_343)
);


endmodule