module fake_netlist_6_141_n_1682 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1682);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1682;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_27),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_35),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_55),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_45),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_39),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_6),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_7),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_117),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_66),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_28),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_85),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_8),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_8),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_51),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_49),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_65),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_97),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_132),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_131),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_114),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_27),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_53),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_51),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_21),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_14),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_48),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_115),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_90),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_84),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_58),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_3),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_83),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_49),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_39),
.Y(n_195)
);

BUFx8_ASAP7_75t_SL g196 ( 
.A(n_69),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_33),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_40),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_59),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_22),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_63),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_57),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_36),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_60),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_111),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_1),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_48),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_44),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_18),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_74),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_88),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_144),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_41),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_4),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_40),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_77),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_4),
.Y(n_220)
);

BUFx2_ASAP7_75t_R g221 ( 
.A(n_44),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_37),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_50),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_21),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_46),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_61),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_105),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_36),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_116),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_86),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_53),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_104),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_9),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_62),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_56),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_46),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_148),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_50),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_14),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_98),
.Y(n_240)
);

BUFx8_ASAP7_75t_SL g241 ( 
.A(n_68),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_118),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_25),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_139),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_23),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_93),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_121),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_141),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_102),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_120),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_143),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_42),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_79),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_2),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_107),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_38),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_28),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_15),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_20),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_133),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_12),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_64),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_6),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_138),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_47),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_81),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_41),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_9),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_0),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_71),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_95),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_78),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_137),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_11),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_0),
.Y(n_275)
);

INVx4_ASAP7_75t_R g276 ( 
.A(n_147),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_25),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_31),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_20),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_24),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_29),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_112),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_37),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_123),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_130),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_32),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_29),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_101),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_43),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_1),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_72),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_204),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_204),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_204),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_172),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_198),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_196),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_204),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_235),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_241),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_202),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_169),
.B(n_3),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_204),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_191),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_153),
.Y(n_306)
);

BUFx6f_ASAP7_75t_SL g307 ( 
.A(n_232),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_222),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_169),
.B(n_5),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_178),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_222),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_198),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_178),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_252),
.B(n_5),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_155),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_156),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_252),
.B(n_7),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_160),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_252),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_184),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_222),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_161),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_184),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_179),
.B(n_10),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_165),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_222),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_222),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_250),
.B(n_12),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_251),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_250),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_167),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_158),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_174),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_175),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_250),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_183),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_158),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_258),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_180),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_258),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_185),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_188),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_190),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_228),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_193),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_154),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_200),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_192),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_192),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_194),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_194),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_205),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_151),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_228),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_232),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_225),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_195),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_201),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_293),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_180),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_320),
.B(n_151),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_294),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_294),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_305),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_334),
.B(n_173),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_305),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_305),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_349),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_295),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_359),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_299),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_358),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_299),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_320),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_304),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_304),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_308),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_340),
.B(n_323),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_311),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_327),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_330),
.Y(n_399)
);

BUFx8_ASAP7_75t_L g400 ( 
.A(n_307),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_SL g401 ( 
.A(n_312),
.B(n_281),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_331),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_331),
.B(n_173),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_332),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_333),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_342),
.Y(n_413)
);

AND2x2_ASAP7_75t_SL g414 ( 
.A(n_303),
.B(n_189),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_328),
.B(n_176),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_343),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_345),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_328),
.B(n_176),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_320),
.B(n_256),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_344),
.B(n_256),
.Y(n_422)
);

BUFx8_ASAP7_75t_L g423 ( 
.A(n_307),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_314),
.B(n_242),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_351),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_353),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_360),
.B(n_353),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_360),
.B(n_189),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_354),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_297),
.B(n_201),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_369),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_310),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_388),
.B(n_306),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_384),
.B(n_315),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_384),
.B(n_316),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_380),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_429),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_388),
.B(n_318),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_322),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_384),
.B(n_325),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_429),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_371),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_364),
.Y(n_455)
);

AND2x2_ASAP7_75t_SL g456 ( 
.A(n_414),
.B(n_309),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_422),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_364),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

INVx8_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_414),
.B(n_341),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_367),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_367),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_414),
.B(n_346),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_380),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_368),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_371),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_368),
.Y(n_470)
);

OAI21xp33_ASAP7_75t_SL g471 ( 
.A1(n_426),
.A2(n_317),
.B(n_314),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

INVx6_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_385),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_369),
.B(n_310),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_368),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_369),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_366),
.B(n_191),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_370),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_370),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_422),
.B(n_350),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_384),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_371),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_372),
.B(n_357),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_365),
.B(n_360),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_370),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_372),
.B(n_300),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_371),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_376),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_366),
.B(n_242),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_366),
.B(n_317),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_366),
.B(n_152),
.Y(n_498)
);

AND2x2_ASAP7_75t_SL g499 ( 
.A(n_415),
.B(n_248),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_371),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_376),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_415),
.B(n_203),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_421),
.B(n_365),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_386),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_376),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_387),
.Y(n_506)
);

XNOR2x2_ASAP7_75t_L g507 ( 
.A(n_432),
.B(n_324),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_378),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_419),
.B(n_246),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_421),
.B(n_354),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_378),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_378),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_421),
.B(n_152),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_365),
.B(n_335),
.Y(n_514)
);

INVx6_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_389),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_387),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_387),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_426),
.B(n_338),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_377),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_377),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_377),
.Y(n_522)
);

AO22x2_ASAP7_75t_L g523 ( 
.A1(n_432),
.A2(n_238),
.B1(n_243),
.B2(n_257),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_389),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_387),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_419),
.B(n_162),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_430),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_400),
.B(n_339),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_389),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_390),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_390),
.Y(n_531)
);

BUFx4f_ASAP7_75t_L g532 ( 
.A(n_430),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_395),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_390),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_373),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_373),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_395),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_395),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_373),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_SL g540 ( 
.A1(n_432),
.A2(n_210),
.B(n_206),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_430),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_379),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_397),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_397),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_391),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_391),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_373),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_379),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_381),
.B(n_292),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_379),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_400),
.B(n_347),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_373),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_397),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_411),
.B(n_355),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_399),
.Y(n_557)
);

BUFx8_ASAP7_75t_SL g558 ( 
.A(n_401),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_394),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_430),
.A2(n_307),
.B1(n_211),
.B2(n_261),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_430),
.A2(n_220),
.B1(n_206),
.B2(n_211),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_394),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_399),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_373),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_373),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_373),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_394),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_430),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_411),
.B(n_348),
.Y(n_569)
);

AO21x2_ASAP7_75t_L g570 ( 
.A1(n_403),
.A2(n_186),
.B(n_162),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_403),
.B(n_361),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_425),
.B(n_186),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_399),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_373),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_400),
.B(n_352),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_399),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_446),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_443),
.B(n_296),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_571),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_436),
.B(n_430),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_449),
.B(n_182),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_443),
.B(n_302),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_448),
.B(n_456),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_527),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_460),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_446),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_456),
.B(n_430),
.Y(n_587)
);

INVxp33_ASAP7_75t_L g588 ( 
.A(n_542),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_456),
.B(n_430),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_550),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_433),
.B(n_221),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_521),
.B(n_400),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_497),
.B(n_430),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_446),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_L g595 ( 
.A(n_479),
.B(n_191),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_460),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_497),
.B(n_381),
.Y(n_597)
);

OR2x2_ASAP7_75t_SL g598 ( 
.A(n_475),
.B(n_324),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_497),
.B(n_381),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_497),
.B(n_428),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_499),
.B(n_428),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_499),
.B(n_428),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_527),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_499),
.A2(n_248),
.B1(n_262),
.B2(n_253),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_451),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_503),
.B(n_423),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_451),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_571),
.B(n_163),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_463),
.A2(n_329),
.B1(n_262),
.B2(n_187),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_527),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_464),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_541),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_451),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_503),
.B(n_428),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_453),
.B(n_428),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_464),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_466),
.B(n_423),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_465),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_520),
.B(n_423),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_453),
.B(n_428),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_498),
.A2(n_453),
.B1(n_457),
.B2(n_513),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_488),
.B(n_219),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_458),
.B(n_298),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_SL g624 ( 
.A(n_540),
.B(n_150),
.C(n_149),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_457),
.B(n_502),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_509),
.B(n_428),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_452),
.B(n_301),
.Y(n_627)
);

NAND2x1p5_ASAP7_75t_L g628 ( 
.A(n_568),
.B(n_187),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_434),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_498),
.B(n_428),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_498),
.B(n_374),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_445),
.B(n_374),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_510),
.B(n_197),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_510),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_465),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_445),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_L g637 ( 
.A1(n_435),
.A2(n_247),
.B1(n_234),
.B2(n_240),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_513),
.B(n_197),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_455),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_468),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_519),
.A2(n_244),
.B1(n_273),
.B2(n_271),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_541),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_513),
.B(n_212),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_455),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_568),
.B(n_423),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_514),
.B(n_159),
.C(n_157),
.Y(n_646)
);

NOR2xp67_ASAP7_75t_L g647 ( 
.A(n_569),
.B(n_411),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_459),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_556),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_468),
.Y(n_650)
);

BUFx12f_ASAP7_75t_SL g651 ( 
.A(n_513),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_526),
.A2(n_247),
.B1(n_283),
.B2(n_272),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_532),
.B(n_423),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_470),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_551),
.B(n_374),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_496),
.B(n_374),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_550),
.B(n_355),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_491),
.B(n_410),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_493),
.B(n_410),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_556),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_470),
.B(n_410),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_477),
.B(n_410),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_477),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_532),
.B(n_423),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_482),
.B(n_483),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_478),
.B(n_356),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_482),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_483),
.B(n_410),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_492),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_532),
.B(n_191),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_461),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_541),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_492),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_526),
.A2(n_264),
.B1(n_212),
.B2(n_230),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_L g675 ( 
.A(n_484),
.B(n_166),
.C(n_164),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_471),
.A2(n_213),
.B1(n_207),
.B2(n_215),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_532),
.B(n_191),
.Y(n_677)
);

AOI22x1_ASAP7_75t_L g678 ( 
.A1(n_526),
.A2(n_523),
.B1(n_501),
.B2(n_505),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_495),
.B(n_425),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_435),
.B(n_475),
.C(n_522),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_501),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_522),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_461),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_508),
.B(n_425),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_508),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_471),
.B(n_168),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_511),
.B(n_427),
.Y(n_687)
);

NOR2x2_ASAP7_75t_L g688 ( 
.A(n_507),
.B(n_254),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_552),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_512),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_552),
.B(n_356),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_526),
.B(n_382),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_516),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_523),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_570),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_523),
.B(n_362),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_516),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_524),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_438),
.B(n_170),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_524),
.B(n_529),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_439),
.B(n_171),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_529),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_523),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_530),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_530),
.B(n_531),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_531),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_534),
.B(n_427),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_534),
.B(n_431),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_545),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_450),
.A2(n_272),
.B1(n_230),
.B2(n_234),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_545),
.B(n_431),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_528),
.A2(n_286),
.B1(n_227),
.B2(n_229),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_547),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_547),
.B(n_548),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_479),
.B(n_264),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_553),
.A2(n_226),
.B1(n_249),
.B2(n_255),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_476),
.B(n_382),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_548),
.B(n_431),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_515),
.A2(n_289),
.B1(n_260),
.B2(n_266),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_473),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_559),
.B(n_562),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_570),
.A2(n_412),
.B1(n_431),
.B2(n_220),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_559),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_562),
.A2(n_287),
.B(n_231),
.C(n_238),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_567),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_567),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_476),
.B(n_396),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_441),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_476),
.B(n_485),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_575),
.A2(n_285),
.B1(n_270),
.B2(n_268),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_485),
.B(n_572),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_570),
.A2(n_412),
.B1(n_217),
.B2(n_261),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_485),
.B(n_396),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_444),
.B(n_396),
.Y(n_734)
);

INVx11_ASAP7_75t_L g735 ( 
.A(n_588),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_579),
.B(n_558),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_634),
.B(n_362),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_725),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_583),
.B(n_444),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_725),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_577),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_593),
.A2(n_494),
.B(n_444),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_622),
.B(n_444),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_622),
.B(n_494),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_L g745 ( 
.A1(n_587),
.A2(n_560),
.B(n_447),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_581),
.B(n_507),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_720),
.B(n_440),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_625),
.B(n_581),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_720),
.A2(n_671),
.B(n_729),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_589),
.A2(n_447),
.B(n_441),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_L g751 ( 
.A(n_680),
.B(n_181),
.C(n_177),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_610),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_720),
.A2(n_461),
.B(n_442),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_671),
.A2(n_461),
.B(n_442),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_610),
.B(n_440),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_586),
.Y(n_756)
);

AO21x1_ASAP7_75t_L g757 ( 
.A1(n_617),
.A2(n_243),
.B(n_231),
.Y(n_757)
);

AO21x1_ASAP7_75t_L g758 ( 
.A1(n_617),
.A2(n_609),
.B(n_602),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_585),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_666),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_594),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_699),
.B(n_494),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_699),
.B(n_494),
.Y(n_763)
);

BUFx2_ASAP7_75t_SL g764 ( 
.A(n_682),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_701),
.B(n_536),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_608),
.B(n_277),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_671),
.A2(n_461),
.B(n_442),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_621),
.A2(n_515),
.B1(n_473),
.B2(n_572),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_608),
.B(n_282),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_701),
.B(n_536),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_634),
.B(n_647),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_604),
.A2(n_515),
.B1(n_473),
.B2(n_572),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_649),
.B(n_536),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_610),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_671),
.A2(n_442),
.B(n_437),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_691),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_660),
.B(n_539),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_L g778 ( 
.A(n_689),
.B(n_539),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_610),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_607),
.B(n_539),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_613),
.B(n_539),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_596),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_657),
.B(n_590),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_612),
.B(n_440),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_601),
.A2(n_447),
.B(n_441),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_614),
.A2(n_474),
.B(n_462),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_578),
.B(n_363),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_588),
.B(n_473),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_729),
.A2(n_454),
.B(n_437),
.Y(n_789)
);

NOR2x1_ASAP7_75t_R g790 ( 
.A(n_582),
.B(n_199),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_612),
.B(n_440),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_694),
.A2(n_572),
.B(n_481),
.C(n_486),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_703),
.A2(n_572),
.B(n_481),
.C(n_486),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_584),
.A2(n_454),
.B(n_437),
.Y(n_794)
);

INVx11_ASAP7_75t_L g795 ( 
.A(n_624),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_673),
.B(n_549),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_627),
.B(n_209),
.C(n_208),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_612),
.B(n_440),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_681),
.B(n_549),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_686),
.A2(n_554),
.B(n_565),
.C(n_564),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_584),
.Y(n_801)
);

OAI21xp33_ASAP7_75t_L g802 ( 
.A1(n_686),
.A2(n_730),
.B(n_627),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_611),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_605),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_584),
.A2(n_535),
.B(n_500),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_605),
.A2(n_642),
.B1(n_672),
.B2(n_603),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_693),
.B(n_554),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_611),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_612),
.B(n_440),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_623),
.B(n_454),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_642),
.A2(n_561),
.B1(n_554),
.B2(n_565),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_695),
.A2(n_576),
.B(n_506),
.Y(n_812)
);

AOI21x1_ASAP7_75t_L g813 ( 
.A1(n_717),
.A2(n_480),
.B(n_467),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_603),
.A2(n_487),
.B(n_535),
.Y(n_814)
);

NOR2xp67_ASAP7_75t_L g815 ( 
.A(n_712),
.B(n_564),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_702),
.B(n_564),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_603),
.A2(n_487),
.B(n_535),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_704),
.B(n_564),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_683),
.A2(n_487),
.B(n_535),
.Y(n_819)
);

NAND2x1_ASAP7_75t_L g820 ( 
.A(n_683),
.B(n_565),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_616),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_706),
.B(n_565),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_731),
.B(n_683),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_709),
.B(n_487),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_623),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_713),
.B(n_500),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_618),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_723),
.B(n_500),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_695),
.A2(n_576),
.B(n_474),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_659),
.B(n_500),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_638),
.A2(n_576),
.B(n_573),
.C(n_563),
.Y(n_831)
);

INVx11_ASAP7_75t_L g832 ( 
.A(n_592),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_638),
.B(n_566),
.Y(n_833)
);

NOR2x2_ASAP7_75t_L g834 ( 
.A(n_688),
.B(n_214),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_672),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_618),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_633),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_731),
.B(n_469),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_692),
.B(n_566),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_638),
.B(n_566),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_635),
.Y(n_841)
);

BUFx4f_ASAP7_75t_L g842 ( 
.A(n_696),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_643),
.B(n_479),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_717),
.A2(n_472),
.B(n_467),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_643),
.B(n_479),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_643),
.B(n_479),
.Y(n_846)
);

AO21x1_ASAP7_75t_L g847 ( 
.A1(n_606),
.A2(n_257),
.B(n_259),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_628),
.Y(n_848)
);

AOI21x1_ASAP7_75t_L g849 ( 
.A1(n_580),
.A2(n_472),
.B(n_525),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_635),
.B(n_479),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_640),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_600),
.A2(n_462),
.B(n_573),
.Y(n_852)
);

AO21x1_ASAP7_75t_L g853 ( 
.A1(n_606),
.A2(n_710),
.B(n_677),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_628),
.B(n_469),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_633),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_650),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_633),
.B(n_363),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_650),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_654),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_597),
.A2(n_469),
.B(n_574),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_688),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_724),
.A2(n_287),
.B(n_259),
.C(n_290),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_599),
.A2(n_469),
.B(n_574),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_631),
.A2(n_474),
.B(n_573),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_656),
.A2(n_469),
.B(n_574),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_663),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_663),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_667),
.B(n_462),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_667),
.B(n_537),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_637),
.A2(n_700),
.B(n_705),
.C(n_714),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_669),
.B(n_537),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_669),
.B(n_489),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_676),
.A2(n_490),
.B(n_563),
.C(n_557),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_655),
.A2(n_574),
.B(n_382),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_651),
.B(n_216),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_665),
.A2(n_290),
.B(n_408),
.C(n_409),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_658),
.A2(n_490),
.B(n_557),
.C(n_555),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_685),
.B(n_690),
.Y(n_878)
);

AOI21xp33_ASAP7_75t_L g879 ( 
.A1(n_641),
.A2(n_233),
.B(n_218),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_651),
.B(n_223),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_724),
.A2(n_416),
.B(n_413),
.C(n_418),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_615),
.A2(n_574),
.B(n_382),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_685),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_690),
.Y(n_884)
);

OAI21xp33_ASAP7_75t_L g885 ( 
.A1(n_652),
.A2(n_236),
.B(n_224),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_626),
.A2(n_557),
.B(n_555),
.C(n_546),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_697),
.B(n_489),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_697),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_630),
.A2(n_555),
.B(n_546),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_629),
.A2(n_546),
.B(n_544),
.C(n_543),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_698),
.B(n_489),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_620),
.A2(n_382),
.B(n_543),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_698),
.B(n_504),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_727),
.A2(n_733),
.B(n_692),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_721),
.A2(n_382),
.B(n_543),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_661),
.A2(n_544),
.B(n_538),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_632),
.A2(n_382),
.B(n_538),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_726),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_598),
.B(n_239),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_726),
.B(n_544),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_678),
.B(n_504),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_670),
.A2(n_533),
.B(n_518),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_662),
.A2(n_533),
.B(n_518),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_670),
.A2(n_533),
.B(n_518),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_645),
.B(n_504),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_636),
.Y(n_906)
);

NOR2x1_ASAP7_75t_L g907 ( 
.A(n_645),
.B(n_398),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_639),
.B(n_506),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_L g909 ( 
.A(n_646),
.B(n_245),
.C(n_275),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_677),
.A2(n_517),
.B(n_506),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_842),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_801),
.A2(n_772),
.B(n_768),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_748),
.B(n_801),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_813),
.A2(n_687),
.B(n_707),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_783),
.B(n_591),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_825),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_SL g917 ( 
.A(n_746),
.B(n_899),
.C(n_769),
.Y(n_917)
);

CKINVDCx16_ASAP7_75t_R g918 ( 
.A(n_764),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_760),
.B(n_675),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_894),
.A2(n_800),
.B(n_739),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_759),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_766),
.B(n_716),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_SL g923 ( 
.A(n_746),
.B(n_619),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_810),
.B(n_644),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_787),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_749),
.A2(n_753),
.B(n_830),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_833),
.A2(n_653),
.B(n_664),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_766),
.B(n_648),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_883),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_840),
.A2(n_747),
.B(n_762),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_827),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_776),
.B(n_760),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_747),
.A2(n_765),
.B(n_763),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_836),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_SL g935 ( 
.A(n_899),
.B(n_269),
.C(n_265),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_810),
.A2(n_664),
.B1(n_653),
.B2(n_674),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_879),
.A2(n_668),
.B(n_719),
.C(n_679),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_743),
.B(n_684),
.Y(n_938)
);

NOR2x1_ASAP7_75t_SL g939 ( 
.A(n_752),
.B(n_728),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_835),
.A2(n_732),
.B1(n_718),
.B2(n_708),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_735),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_883),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_770),
.A2(n_595),
.B(n_734),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_744),
.B(n_711),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_819),
.A2(n_595),
.B(n_715),
.Y(n_945)
);

BUFx8_ASAP7_75t_L g946 ( 
.A(n_737),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_835),
.B(n_866),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_857),
.B(n_722),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_883),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_771),
.B(n_214),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_782),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_779),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_788),
.B(n_214),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_L g954 ( 
.A1(n_797),
.A2(n_291),
.B(n_263),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_788),
.B(n_237),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_795),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_867),
.B(n_517),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_888),
.B(n_517),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_803),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_797),
.A2(n_715),
.B(n_424),
.C(n_418),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_848),
.B(n_237),
.Y(n_961)
);

AO32x1_ASAP7_75t_L g962 ( 
.A1(n_898),
.A2(n_406),
.A3(n_398),
.B1(n_404),
.B2(n_405),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_906),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_808),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_878),
.B(n_398),
.Y(n_965)
);

NOR2x1_ASAP7_75t_R g966 ( 
.A(n_737),
.B(n_267),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_806),
.A2(n_284),
.B1(n_288),
.B2(n_280),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_L g968 ( 
.A1(n_853),
.A2(n_418),
.B(n_413),
.C(n_416),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_906),
.B(n_413),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_821),
.B(n_405),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_823),
.A2(n_279),
.B1(n_278),
.B2(n_416),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_861),
.B(n_237),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_848),
.B(n_232),
.Y(n_973)
);

BUFx12f_ASAP7_75t_L g974 ( 
.A(n_857),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_841),
.B(n_405),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_851),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_870),
.A2(n_424),
.B(n_417),
.C(n_404),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_804),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_804),
.B(n_232),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_SL g980 ( 
.A1(n_854),
.A2(n_404),
.B(n_406),
.C(n_409),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_837),
.B(n_424),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_856),
.B(n_409),
.Y(n_982)
);

NAND3xp33_ASAP7_75t_L g983 ( 
.A(n_751),
.B(n_408),
.C(n_407),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_854),
.A2(n_375),
.B(n_276),
.Y(n_984)
);

AO32x2_ASAP7_75t_L g985 ( 
.A1(n_855),
.A2(n_13),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_792),
.A2(n_417),
.B(n_408),
.C(n_407),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_823),
.A2(n_375),
.B(n_393),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_793),
.A2(n_875),
.B(n_880),
.C(n_738),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_848),
.B(n_417),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_858),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_754),
.A2(n_375),
.B(n_393),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_751),
.A2(n_407),
.B(n_417),
.C(n_393),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_740),
.B(n_412),
.Y(n_993)
);

NAND2x1_ASAP7_75t_SL g994 ( 
.A(n_779),
.B(n_392),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_736),
.B(n_741),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_862),
.A2(n_392),
.B(n_393),
.C(n_402),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_859),
.B(n_393),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_862),
.A2(n_392),
.B(n_393),
.C(n_402),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_875),
.A2(n_392),
.B(n_375),
.C(n_402),
.Y(n_999)
);

NAND2x1p5_ASAP7_75t_L g1000 ( 
.A(n_774),
.B(n_392),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_883),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_884),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_884),
.B(n_392),
.Y(n_1003)
);

O2A1O1Ixp5_ASAP7_75t_L g1004 ( 
.A1(n_757),
.A2(n_402),
.B(n_73),
.C(n_146),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_756),
.Y(n_1005)
);

O2A1O1Ixp5_ASAP7_75t_L g1006 ( 
.A1(n_847),
.A2(n_67),
.B(n_145),
.C(n_134),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_SL g1007 ( 
.A1(n_838),
.A2(n_16),
.B(n_17),
.Y(n_1007)
);

AOI22x1_ASAP7_75t_L g1008 ( 
.A1(n_905),
.A2(n_412),
.B1(n_383),
.B2(n_70),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_767),
.A2(n_383),
.B(n_412),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_736),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_884),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_761),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_790),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_794),
.A2(n_383),
.B(n_412),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_805),
.A2(n_383),
.B(n_412),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_774),
.B(n_412),
.Y(n_1016)
);

CKINVDCx11_ASAP7_75t_R g1017 ( 
.A(n_834),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_814),
.A2(n_383),
.B(n_54),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_773),
.B(n_383),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_844),
.A2(n_76),
.B(n_128),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_909),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_838),
.A2(n_383),
.B1(n_126),
.B2(n_125),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_778),
.B(n_19),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_742),
.A2(n_849),
.B(n_892),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_817),
.A2(n_383),
.B(n_124),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_832),
.B(n_19),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_789),
.A2(n_119),
.B(n_113),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_905),
.A2(n_109),
.B1(n_106),
.B2(n_100),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_815),
.B(n_99),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_881),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_777),
.B(n_824),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_826),
.B(n_26),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_881),
.A2(n_26),
.B(n_30),
.C(n_31),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_745),
.A2(n_30),
.B(n_33),
.C(n_34),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_828),
.B(n_94),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_755),
.B(n_91),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_908),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_775),
.A2(n_92),
.B(n_89),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_872),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_755),
.B(n_784),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_868),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_869),
.B(n_34),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_885),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_843),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_839),
.A2(n_35),
.B1(n_38),
.B2(n_42),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_871),
.B(n_43),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_845),
.B(n_45),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_913),
.B(n_1037),
.Y(n_1048)
);

AOI221x1_ASAP7_75t_L g1049 ( 
.A1(n_1034),
.A2(n_886),
.B1(n_873),
.B2(n_831),
.C(n_829),
.Y(n_1049)
);

AO31x2_ASAP7_75t_L g1050 ( 
.A1(n_936),
.A2(n_890),
.A3(n_877),
.B(n_895),
.Y(n_1050)
);

AO21x1_ASAP7_75t_L g1051 ( 
.A1(n_922),
.A2(n_901),
.B(n_876),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_929),
.Y(n_1052)
);

AND2x6_ASAP7_75t_L g1053 ( 
.A(n_1036),
.B(n_907),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_918),
.Y(n_1054)
);

CKINVDCx6p67_ASAP7_75t_R g1055 ( 
.A(n_974),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_913),
.B(n_891),
.Y(n_1056)
);

CKINVDCx11_ASAP7_75t_R g1057 ( 
.A(n_1017),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_917),
.A2(n_923),
.B(n_928),
.C(n_988),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_915),
.B(n_780),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_948),
.B(n_781),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1039),
.B(n_893),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_912),
.A2(n_901),
.B(n_904),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_SL g1063 ( 
.A(n_916),
.B(n_846),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_941),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_SL g1065 ( 
.A1(n_1029),
.A2(n_798),
.B(n_809),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_969),
.B(n_796),
.Y(n_1066)
);

AO31x2_ASAP7_75t_L g1067 ( 
.A1(n_977),
.A2(n_933),
.A3(n_986),
.B(n_926),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_920),
.A2(n_812),
.B(n_791),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_924),
.A2(n_839),
.B1(n_811),
.B2(n_807),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1005),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_995),
.B(n_822),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1012),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_963),
.B(n_816),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_911),
.B(n_818),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_931),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1044),
.B(n_799),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_930),
.A2(n_874),
.B(n_900),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_938),
.A2(n_750),
.B(n_865),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_938),
.A2(n_785),
.B(n_863),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_944),
.A2(n_860),
.B(n_786),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_934),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_1043),
.A2(n_850),
.B1(n_868),
.B2(n_900),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_944),
.A2(n_852),
.B(n_864),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1031),
.A2(n_943),
.B(n_937),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1024),
.A2(n_910),
.B(n_902),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_919),
.B(n_887),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_981),
.B(n_887),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_929),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_914),
.A2(n_882),
.B(n_897),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_942),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_SL g1091 ( 
.A1(n_1030),
.A2(n_1033),
.B(n_939),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_978),
.B(n_889),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_946),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1009),
.A2(n_903),
.B(n_896),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1031),
.A2(n_820),
.B1(n_47),
.B2(n_52),
.Y(n_1095)
);

AO31x2_ASAP7_75t_L g1096 ( 
.A1(n_940),
.A2(n_52),
.A3(n_984),
.B(n_999),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_965),
.B(n_947),
.Y(n_1097)
);

AOI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1035),
.A2(n_1032),
.B(n_1046),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_1018),
.A2(n_1025),
.A3(n_945),
.B(n_1042),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_SL g1100 ( 
.A(n_956),
.B(n_1026),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_1013),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1046),
.A2(n_965),
.B(n_1019),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_972),
.B(n_1021),
.Y(n_1103)
);

BUFx10_ASAP7_75t_L g1104 ( 
.A(n_979),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_942),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_947),
.B(n_1041),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_954),
.A2(n_1029),
.B(n_960),
.C(n_1007),
.Y(n_1107)
);

OR2x6_ASAP7_75t_L g1108 ( 
.A(n_949),
.B(n_1001),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1019),
.A2(n_1027),
.B(n_968),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_SL g1110 ( 
.A(n_935),
.B(n_1010),
.C(n_950),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1038),
.A2(n_955),
.B(n_953),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_SL g1112 ( 
.A(n_966),
.B(n_1045),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1014),
.A2(n_1015),
.B(n_1016),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_970),
.A2(n_982),
.B(n_975),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1020),
.A2(n_991),
.B(n_1016),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1004),
.A2(n_992),
.B(n_983),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1028),
.A2(n_1036),
.B1(n_967),
.B2(n_1022),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_SL g1118 ( 
.A1(n_973),
.A2(n_961),
.B(n_989),
.C(n_1003),
.Y(n_1118)
);

AOI21x1_ASAP7_75t_L g1119 ( 
.A1(n_970),
.A2(n_982),
.B(n_975),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_962),
.A2(n_958),
.A3(n_957),
.B(n_1003),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_921),
.B(n_964),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_932),
.A2(n_971),
.B(n_1006),
.C(n_1023),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_976),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_987),
.A2(n_957),
.B(n_958),
.Y(n_1124)
);

BUFx2_ASAP7_75t_R g1125 ( 
.A(n_952),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_951),
.B(n_959),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_SL g1127 ( 
.A(n_1047),
.B(n_990),
.C(n_996),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_952),
.B(n_1011),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1008),
.A2(n_997),
.B(n_998),
.Y(n_1129)
);

NOR2x1_ASAP7_75t_SL g1130 ( 
.A(n_949),
.B(n_1001),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_997),
.A2(n_1040),
.B(n_980),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1002),
.B(n_1040),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_949),
.A2(n_1001),
.B1(n_993),
.B2(n_1000),
.Y(n_1133)
);

AOI221x1_ASAP7_75t_L g1134 ( 
.A1(n_985),
.A2(n_802),
.B1(n_746),
.B2(n_1034),
.C(n_922),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_994),
.A2(n_985),
.B(n_1000),
.C(n_962),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_962),
.A2(n_758),
.A3(n_853),
.B(n_936),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_985),
.A2(n_720),
.B(n_671),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_922),
.A2(n_746),
.B1(n_769),
.B2(n_766),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1024),
.A2(n_742),
.B(n_849),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_916),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_927),
.A2(n_720),
.B(n_671),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1024),
.A2(n_742),
.B(n_849),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_927),
.A2(n_720),
.B(n_671),
.Y(n_1143)
);

NAND3xp33_ASAP7_75t_L g1144 ( 
.A(n_922),
.B(n_769),
.C(n_766),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_916),
.Y(n_1145)
);

AO21x2_ASAP7_75t_L g1146 ( 
.A1(n_920),
.A2(n_912),
.B(n_926),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_918),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_927),
.A2(n_720),
.B(n_671),
.Y(n_1148)
);

BUFx10_ASAP7_75t_L g1149 ( 
.A(n_916),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_913),
.B(n_583),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_941),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1005),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_922),
.A2(n_746),
.B(n_769),
.C(n_766),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_927),
.A2(n_720),
.B(n_671),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_922),
.A2(n_766),
.B1(n_769),
.B2(n_746),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1024),
.A2(n_742),
.B(n_849),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_927),
.A2(n_720),
.B(n_671),
.Y(n_1157)
);

AOI21x1_ASAP7_75t_L g1158 ( 
.A1(n_927),
.A2(n_930),
.B(n_933),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_SL g1159 ( 
.A(n_922),
.B(n_769),
.C(n_766),
.Y(n_1159)
);

AO31x2_ASAP7_75t_L g1160 ( 
.A1(n_936),
.A2(n_758),
.A3(n_853),
.B(n_757),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_922),
.A2(n_746),
.B(n_769),
.C(n_766),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1005),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_L g1163 ( 
.A1(n_927),
.A2(n_930),
.B(n_933),
.Y(n_1163)
);

BUFx8_ASAP7_75t_L g1164 ( 
.A(n_1013),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_916),
.B(n_925),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_927),
.A2(n_720),
.B(n_671),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1024),
.A2(n_742),
.B(n_849),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_928),
.B(n_748),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_L g1169 ( 
.A(n_922),
.B(n_769),
.C(n_766),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_936),
.A2(n_758),
.A3(n_853),
.B(n_757),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_927),
.A2(n_720),
.B(n_671),
.Y(n_1171)
);

OAI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_922),
.A2(n_769),
.B(n_766),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_SL g1173 ( 
.A(n_922),
.B(n_769),
.C(n_766),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_941),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_941),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_922),
.B(n_746),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_941),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1070),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1052),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1072),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1140),
.Y(n_1181)
);

INVx6_ASAP7_75t_L g1182 ( 
.A(n_1149),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1084),
.A2(n_1083),
.B(n_1137),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1176),
.A2(n_1159),
.B1(n_1173),
.B2(n_1138),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1172),
.A2(n_1144),
.B1(n_1169),
.B2(n_1155),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1144),
.A2(n_1169),
.B1(n_1112),
.B2(n_1103),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1112),
.A2(n_1117),
.B1(n_1110),
.B2(n_1100),
.Y(n_1187)
);

BUFx8_ASAP7_75t_SL g1188 ( 
.A(n_1064),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1152),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_SL g1190 ( 
.A1(n_1153),
.A2(n_1161),
.B1(n_1095),
.B2(n_1100),
.Y(n_1190)
);

BUFx8_ASAP7_75t_L g1191 ( 
.A(n_1093),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1162),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1168),
.A2(n_1048),
.B1(n_1071),
.B2(n_1150),
.Y(n_1193)
);

CKINVDCx11_ASAP7_75t_R g1194 ( 
.A(n_1057),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1048),
.B(n_1059),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_SL g1196 ( 
.A1(n_1095),
.A2(n_1053),
.B1(n_1104),
.B2(n_1134),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1145),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1149),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1051),
.A2(n_1086),
.B1(n_1053),
.B2(n_1150),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_SL g1200 ( 
.A1(n_1053),
.A2(n_1104),
.B1(n_1091),
.B2(n_1092),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1075),
.Y(n_1201)
);

CKINVDCx11_ASAP7_75t_R g1202 ( 
.A(n_1055),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1060),
.B(n_1058),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1053),
.A2(n_1074),
.B1(n_1127),
.B2(n_1132),
.Y(n_1204)
);

OAI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1073),
.A2(n_1097),
.B1(n_1066),
.B2(n_1081),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1052),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1147),
.A2(n_1165),
.B1(n_1063),
.B2(n_1146),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1146),
.A2(n_1076),
.B1(n_1116),
.B2(n_1082),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_SL g1209 ( 
.A1(n_1069),
.A2(n_1068),
.B1(n_1097),
.B2(n_1116),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1069),
.A2(n_1056),
.B1(n_1164),
.B2(n_1123),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1108),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1121),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1126),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1151),
.Y(n_1214)
);

BUFx2_ASAP7_75t_SL g1215 ( 
.A(n_1174),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1101),
.A2(n_1107),
.B1(n_1118),
.B2(n_1164),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1106),
.B(n_1061),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1126),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1056),
.A2(n_1106),
.B1(n_1087),
.B2(n_1111),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1175),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_1177),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1062),
.A2(n_1131),
.B1(n_1078),
.B2(n_1080),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1125),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1088),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1049),
.A2(n_1119),
.B1(n_1114),
.B2(n_1128),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1079),
.A2(n_1133),
.B1(n_1109),
.B2(n_1090),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1105),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1124),
.A2(n_1094),
.B1(n_1113),
.B2(n_1129),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1139),
.A2(n_1142),
.B1(n_1156),
.B2(n_1167),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1130),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1096),
.Y(n_1231)
);

BUFx4f_ASAP7_75t_SL g1232 ( 
.A(n_1065),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1122),
.Y(n_1233)
);

INVx4_ASAP7_75t_SL g1234 ( 
.A(n_1096),
.Y(n_1234)
);

OAI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1102),
.A2(n_1098),
.B1(n_1158),
.B2(n_1163),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1096),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_1141),
.Y(n_1237)
);

CKINVDCx6p67_ASAP7_75t_R g1238 ( 
.A(n_1135),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1115),
.A2(n_1143),
.B1(n_1166),
.B2(n_1157),
.Y(n_1239)
);

CKINVDCx6p67_ASAP7_75t_R g1240 ( 
.A(n_1120),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1077),
.A2(n_1171),
.B1(n_1154),
.B2(n_1148),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1120),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1067),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1089),
.A2(n_1085),
.B1(n_1170),
.B2(n_1160),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1160),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1067),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_1160),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_1170),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1170),
.Y(n_1249)
);

BUFx12f_ASAP7_75t_L g1250 ( 
.A(n_1099),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1099),
.Y(n_1251)
);

BUFx4f_ASAP7_75t_L g1252 ( 
.A(n_1099),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1136),
.A2(n_1176),
.B1(n_1159),
.B2(n_1173),
.Y(n_1253)
);

BUFx8_ASAP7_75t_SL g1254 ( 
.A(n_1050),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1140),
.Y(n_1255)
);

INVx3_ASAP7_75t_SL g1256 ( 
.A(n_1140),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1176),
.A2(n_1138),
.B1(n_1155),
.B2(n_1144),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1176),
.A2(n_1138),
.B1(n_746),
.B2(n_1159),
.Y(n_1258)
);

CKINVDCx11_ASAP7_75t_R g1259 ( 
.A(n_1057),
.Y(n_1259)
);

OAI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1155),
.A2(n_1176),
.B1(n_923),
.B2(n_746),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1165),
.B(n_911),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1054),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1052),
.Y(n_1263)
);

CKINVDCx11_ASAP7_75t_R g1264 ( 
.A(n_1057),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1070),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1176),
.B(n_1103),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1176),
.A2(n_746),
.B1(n_769),
.B2(n_766),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1155),
.A2(n_1176),
.B1(n_923),
.B2(n_746),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1084),
.A2(n_936),
.B(n_1083),
.Y(n_1269)
);

AOI21xp33_ASAP7_75t_L g1270 ( 
.A1(n_1153),
.A2(n_1161),
.B(n_1172),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1176),
.A2(n_1138),
.B1(n_1155),
.B2(n_1144),
.Y(n_1271)
);

OAI21xp33_ASAP7_75t_L g1272 ( 
.A1(n_1176),
.A2(n_1138),
.B(n_1155),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1151),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1151),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1176),
.A2(n_1138),
.B1(n_746),
.B2(n_1159),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1057),
.Y(n_1276)
);

OAI21xp33_ASAP7_75t_L g1277 ( 
.A1(n_1176),
.A2(n_1138),
.B(n_1155),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1176),
.A2(n_746),
.B1(n_923),
.B2(n_1144),
.Y(n_1278)
);

CKINVDCx6p67_ASAP7_75t_R g1279 ( 
.A(n_1064),
.Y(n_1279)
);

INVx11_ASAP7_75t_L g1280 ( 
.A(n_1064),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1070),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1176),
.A2(n_1159),
.B1(n_1173),
.B2(n_1138),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1176),
.A2(n_1155),
.B1(n_1173),
.B2(n_1159),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1176),
.A2(n_1138),
.B1(n_746),
.B2(n_1159),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1149),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1176),
.A2(n_1138),
.B1(n_746),
.B2(n_1159),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1176),
.A2(n_1138),
.B1(n_746),
.B2(n_1159),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1250),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1236),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_1194),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1254),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1249),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1242),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1231),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1180),
.Y(n_1295)
);

INVxp33_ASAP7_75t_L g1296 ( 
.A(n_1262),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1234),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1182),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1182),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_SL g1300 ( 
.A1(n_1260),
.A2(n_1268),
.B(n_1257),
.C(n_1271),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1243),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1251),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1248),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1233),
.B(n_1252),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1178),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1189),
.Y(n_1306)
);

OR2x2_ASAP7_75t_L g1307 ( 
.A(n_1203),
.B(n_1240),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1192),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1182),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1285),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1245),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1211),
.B(n_1201),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1235),
.A2(n_1241),
.B(n_1269),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1187),
.A2(n_1283),
.B1(n_1260),
.B2(n_1268),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1233),
.B(n_1252),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1247),
.Y(n_1316)
);

AO21x1_ASAP7_75t_L g1317 ( 
.A1(n_1270),
.A2(n_1205),
.B(n_1225),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1224),
.Y(n_1318)
);

CKINVDCx10_ASAP7_75t_R g1319 ( 
.A(n_1259),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1285),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1285),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1246),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1265),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_R g1324 ( 
.A(n_1181),
.B(n_1197),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1281),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1227),
.Y(n_1326)
);

AO21x2_ASAP7_75t_L g1327 ( 
.A1(n_1235),
.A2(n_1241),
.B(n_1269),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1195),
.B(n_1266),
.Y(n_1328)
);

CKINVDCx14_ASAP7_75t_R g1329 ( 
.A(n_1264),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1183),
.A2(n_1193),
.B(n_1217),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1272),
.A2(n_1277),
.B1(n_1278),
.B2(n_1284),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1232),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1183),
.A2(n_1229),
.B(n_1228),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1205),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1229),
.A2(n_1228),
.B(n_1239),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1225),
.A2(n_1222),
.B(n_1209),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1212),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1239),
.A2(n_1222),
.B(n_1244),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1237),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1213),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1218),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1232),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1267),
.A2(n_1278),
.B1(n_1287),
.B2(n_1275),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1253),
.B(n_1199),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1238),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1209),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1185),
.A2(n_1219),
.B(n_1226),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1244),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1258),
.A2(n_1286),
.B1(n_1275),
.B2(n_1284),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1219),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1230),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1208),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1196),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1196),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1200),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1200),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1186),
.B(n_1185),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1221),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1216),
.A2(n_1198),
.B(n_1261),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1210),
.B(n_1190),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1210),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1190),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1207),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1204),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1184),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1258),
.B(n_1287),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1282),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1300),
.A2(n_1286),
.B(n_1261),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1343),
.A2(n_1331),
.B1(n_1349),
.B2(n_1345),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1305),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1336),
.A2(n_1223),
.B(n_1215),
.C(n_1273),
.Y(n_1371)
);

AND2x2_ASAP7_75t_SL g1372 ( 
.A(n_1360),
.B(n_1223),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1333),
.A2(n_1179),
.B(n_1263),
.Y(n_1373)
);

NAND2xp33_ASAP7_75t_R g1374 ( 
.A(n_1291),
.B(n_1191),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1311),
.B(n_1214),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1314),
.A2(n_1367),
.B1(n_1365),
.B2(n_1364),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1317),
.A2(n_1179),
.B(n_1263),
.Y(n_1377)
);

NOR2x1_ASAP7_75t_L g1378 ( 
.A(n_1359),
.B(n_1274),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1316),
.B(n_1214),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1305),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1365),
.B(n_1256),
.Y(n_1381)
);

A2O1A1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1347),
.A2(n_1220),
.B(n_1263),
.C(n_1206),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1367),
.A2(n_1279),
.B1(n_1256),
.B2(n_1202),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1328),
.B(n_1255),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1297),
.B(n_1280),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1318),
.B(n_1255),
.Y(n_1386)
);

NAND3xp33_ASAP7_75t_L g1387 ( 
.A(n_1357),
.B(n_1276),
.C(n_1188),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1357),
.B(n_1307),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1364),
.A2(n_1362),
.B1(n_1366),
.B2(n_1345),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1362),
.A2(n_1339),
.B1(n_1361),
.B2(n_1344),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1312),
.B(n_1361),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1359),
.B(n_1304),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1326),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1317),
.A2(n_1346),
.B(n_1352),
.C(n_1363),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1319),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1304),
.B(n_1315),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1324),
.Y(n_1397)
);

INVx4_ASAP7_75t_SL g1398 ( 
.A(n_1288),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1333),
.A2(n_1338),
.B(n_1335),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1346),
.B(n_1356),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_SL g1402 ( 
.A(n_1358),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1306),
.B(n_1308),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1352),
.A2(n_1363),
.B(n_1334),
.C(n_1353),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1306),
.B(n_1308),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1291),
.A2(n_1354),
.B1(n_1353),
.B2(n_1332),
.Y(n_1406)
);

OR2x2_ASAP7_75t_SL g1407 ( 
.A(n_1298),
.B(n_1288),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_SL g1408 ( 
.A1(n_1330),
.A2(n_1326),
.B(n_1334),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1354),
.B(n_1344),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1338),
.A2(n_1350),
.B(n_1332),
.C(n_1342),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1335),
.A2(n_1289),
.B(n_1294),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1337),
.B(n_1295),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1290),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1350),
.B(n_1332),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1342),
.A2(n_1296),
.B1(n_1315),
.B2(n_1304),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1323),
.B(n_1325),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1342),
.A2(n_1315),
.B1(n_1320),
.B2(n_1310),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1299),
.A2(n_1309),
.B1(n_1320),
.B2(n_1321),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1288),
.B(n_1301),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1411),
.B(n_1313),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1370),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1411),
.B(n_1313),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_1386),
.Y(n_1423)
);

NOR3xp33_ASAP7_75t_L g1424 ( 
.A(n_1369),
.B(n_1329),
.C(n_1351),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1380),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1403),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1400),
.B(n_1327),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_1393),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1405),
.Y(n_1429)
);

NAND2x1_ASAP7_75t_L g1430 ( 
.A(n_1392),
.B(n_1396),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1388),
.B(n_1348),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1416),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_1392),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1388),
.B(n_1393),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1400),
.B(n_1327),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1373),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1412),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1408),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1410),
.B(n_1302),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1391),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1394),
.B(n_1348),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1409),
.B(n_1293),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1410),
.B(n_1293),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1368),
.A2(n_1358),
.B1(n_1341),
.B2(n_1340),
.Y(n_1444)
);

AND2x4_ASAP7_75t_SL g1445 ( 
.A(n_1433),
.B(n_1396),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1433),
.B(n_1396),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1424),
.A2(n_1376),
.B1(n_1390),
.B2(n_1389),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1429),
.B(n_1399),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1434),
.B(n_1302),
.Y(n_1449)
);

OAI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1424),
.A2(n_1371),
.B1(n_1382),
.B2(n_1381),
.C(n_1378),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1423),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1428),
.Y(n_1452)
);

OAI321xp33_ASAP7_75t_L g1453 ( 
.A1(n_1441),
.A2(n_1371),
.A3(n_1382),
.B1(n_1406),
.B2(n_1404),
.C(n_1415),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1429),
.B(n_1443),
.Y(n_1454)
);

AOI31xp33_ASAP7_75t_L g1455 ( 
.A1(n_1444),
.A2(n_1374),
.A3(n_1387),
.B(n_1417),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1441),
.A2(n_1409),
.B1(n_1381),
.B2(n_1401),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1434),
.B(n_1303),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1436),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1444),
.A2(n_1377),
.B(n_1372),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1443),
.B(n_1419),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1443),
.B(n_1301),
.Y(n_1461)
);

NAND2x1_ASAP7_75t_L g1462 ( 
.A(n_1433),
.B(n_1288),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1439),
.B(n_1303),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1432),
.B(n_1414),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1425),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1437),
.B(n_1401),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1439),
.B(n_1442),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1430),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1420),
.A2(n_1289),
.B(n_1292),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1425),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1440),
.B(n_1322),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1423),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1421),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1439),
.B(n_1442),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1433),
.B(n_1398),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1473),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1473),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1470),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1454),
.B(n_1427),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1463),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1470),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1454),
.B(n_1427),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1467),
.B(n_1435),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1454),
.B(n_1427),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1465),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1470),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1467),
.B(n_1474),
.Y(n_1487)
);

NOR3xp33_ASAP7_75t_L g1488 ( 
.A(n_1453),
.B(n_1413),
.C(n_1383),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1453),
.B(n_1433),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1463),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1467),
.B(n_1431),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1474),
.B(n_1431),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1474),
.B(n_1452),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1465),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1448),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1452),
.B(n_1437),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1458),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1463),
.B(n_1435),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1461),
.B(n_1420),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1469),
.B(n_1435),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1448),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1461),
.B(n_1420),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1457),
.B(n_1428),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1458),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_L g1505 ( 
.A(n_1462),
.B(n_1438),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1457),
.B(n_1466),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1461),
.B(n_1422),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1448),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1457),
.B(n_1426),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1481),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1506),
.B(n_1466),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1480),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1489),
.B(n_1455),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1480),
.Y(n_1514)
);

INVxp67_ASAP7_75t_SL g1515 ( 
.A(n_1497),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1506),
.B(n_1449),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1490),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1490),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1491),
.B(n_1492),
.Y(n_1519)
);

OAI321xp33_ASAP7_75t_L g1520 ( 
.A1(n_1489),
.A2(n_1447),
.A3(n_1459),
.B1(n_1450),
.B2(n_1456),
.C(n_1438),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1505),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1487),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1476),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1487),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1476),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1477),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1491),
.B(n_1449),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1493),
.B(n_1449),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1492),
.B(n_1456),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1487),
.B(n_1468),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1481),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1497),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1499),
.B(n_1468),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1493),
.B(n_1472),
.Y(n_1534)
);

INVxp67_ASAP7_75t_SL g1535 ( 
.A(n_1497),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1499),
.B(n_1468),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1481),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1477),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1499),
.B(n_1468),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1502),
.B(n_1460),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1503),
.B(n_1472),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1503),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1481),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1509),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1502),
.B(n_1460),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1483),
.B(n_1471),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1502),
.B(n_1460),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1507),
.B(n_1464),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1509),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1496),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1488),
.B(n_1413),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1513),
.B(n_1488),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1522),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1521),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1522),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1540),
.B(n_1505),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1540),
.B(n_1507),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1529),
.B(n_1496),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1511),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1534),
.B(n_1483),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1521),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_1551),
.Y(n_1562)
);

AOI211xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1520),
.A2(n_1455),
.B(n_1450),
.C(n_1475),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1524),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1511),
.B(n_1495),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1524),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1534),
.B(n_1483),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1540),
.B(n_1507),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1545),
.B(n_1479),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1541),
.B(n_1498),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1542),
.B(n_1495),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1545),
.B(n_1547),
.Y(n_1572)
);

NOR3xp33_ASAP7_75t_L g1573 ( 
.A(n_1520),
.B(n_1459),
.C(n_1462),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1521),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1542),
.B(n_1501),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1550),
.B(n_1519),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1541),
.B(n_1395),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1523),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1550),
.B(n_1501),
.Y(n_1579)
);

OAI32xp33_ASAP7_75t_L g1580 ( 
.A1(n_1512),
.A2(n_1447),
.A3(n_1500),
.B1(n_1451),
.B2(n_1374),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1547),
.B(n_1479),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1519),
.B(n_1395),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1544),
.B(n_1508),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1528),
.B(n_1498),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1544),
.B(n_1508),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1523),
.Y(n_1586)
);

AOI322xp5_ASAP7_75t_L g1587 ( 
.A1(n_1552),
.A2(n_1479),
.A3(n_1482),
.B1(n_1484),
.B2(n_1548),
.C1(n_1539),
.C2(n_1536),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1553),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1553),
.Y(n_1589)
);

OAI322xp33_ASAP7_75t_L g1590 ( 
.A1(n_1559),
.A2(n_1518),
.A3(n_1512),
.B1(n_1514),
.B2(n_1517),
.C1(n_1500),
.C2(n_1528),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1573),
.A2(n_1530),
.B1(n_1446),
.B2(n_1536),
.Y(n_1591)
);

OAI322xp33_ASAP7_75t_L g1592 ( 
.A1(n_1558),
.A2(n_1514),
.A3(n_1518),
.B1(n_1517),
.B2(n_1500),
.C1(n_1549),
.C2(n_1546),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1563),
.B(n_1530),
.Y(n_1593)
);

NOR2x1_ASAP7_75t_L g1594 ( 
.A(n_1562),
.B(n_1451),
.Y(n_1594)
);

OAI31xp33_ASAP7_75t_L g1595 ( 
.A1(n_1556),
.A2(n_1533),
.A3(n_1536),
.B(n_1539),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1564),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1577),
.A2(n_1539),
.B(n_1533),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1582),
.B(n_1549),
.Y(n_1598)
);

OAI21xp33_ASAP7_75t_L g1599 ( 
.A1(n_1580),
.A2(n_1516),
.B(n_1527),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1576),
.B(n_1516),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1562),
.B(n_1475),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1560),
.B(n_1527),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1564),
.B(n_1525),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1556),
.A2(n_1372),
.B1(n_1407),
.B2(n_1445),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1555),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1566),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1566),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1572),
.A2(n_1445),
.B(n_1475),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1561),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1586),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1580),
.B(n_1397),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1588),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1594),
.Y(n_1613)
);

CKINVDCx14_ASAP7_75t_R g1614 ( 
.A(n_1611),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1601),
.B(n_1572),
.Y(n_1615)
);

OAI32xp33_ASAP7_75t_L g1616 ( 
.A1(n_1593),
.A2(n_1560),
.A3(n_1567),
.B1(n_1574),
.B2(n_1554),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1591),
.A2(n_1568),
.B(n_1557),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1609),
.B(n_1569),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1610),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1595),
.B(n_1569),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1597),
.B(n_1581),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1602),
.Y(n_1622)
);

OAI211xp5_ASAP7_75t_L g1623 ( 
.A1(n_1599),
.A2(n_1561),
.B(n_1554),
.C(n_1574),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1589),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1596),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1598),
.B(n_1397),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1605),
.B(n_1581),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1600),
.B(n_1567),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1606),
.B(n_1557),
.Y(n_1629)
);

OAI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1604),
.A2(n_1570),
.B1(n_1433),
.B2(n_1578),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1608),
.B(n_1565),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1629),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1627),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1628),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1618),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1624),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1613),
.A2(n_1607),
.B1(n_1590),
.B2(n_1592),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1625),
.Y(n_1638)
);

OAI322xp33_ASAP7_75t_L g1639 ( 
.A1(n_1614),
.A2(n_1603),
.A3(n_1586),
.B1(n_1570),
.B2(n_1584),
.C1(n_1575),
.C2(n_1571),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1614),
.B(n_1604),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1622),
.B(n_1587),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1634),
.B(n_1612),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1640),
.B(n_1615),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1637),
.A2(n_1623),
.B(n_1641),
.Y(n_1644)
);

NOR3x1_ASAP7_75t_L g1645 ( 
.A(n_1635),
.B(n_1617),
.C(n_1619),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1637),
.B(n_1630),
.Y(n_1646)
);

NAND4xp25_ASAP7_75t_L g1647 ( 
.A(n_1633),
.B(n_1626),
.C(n_1631),
.D(n_1616),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1636),
.Y(n_1648)
);

OAI31xp33_ASAP7_75t_L g1649 ( 
.A1(n_1632),
.A2(n_1626),
.A3(n_1630),
.B(n_1620),
.Y(n_1649)
);

OAI211xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1638),
.A2(n_1631),
.B(n_1603),
.C(n_1584),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1642),
.Y(n_1651)
);

AOI222xp33_ASAP7_75t_L g1652 ( 
.A1(n_1646),
.A2(n_1621),
.B1(n_1639),
.B2(n_1535),
.C1(n_1532),
.C2(n_1515),
.Y(n_1652)
);

AOI21xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1644),
.A2(n_1579),
.B(n_1583),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1649),
.A2(n_1585),
.B(n_1532),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_SL g1655 ( 
.A(n_1647),
.B(n_1402),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1652),
.B(n_1655),
.C(n_1643),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1653),
.B(n_1645),
.Y(n_1657)
);

AOI221xp5_ASAP7_75t_L g1658 ( 
.A1(n_1654),
.A2(n_1650),
.B1(n_1648),
.B2(n_1568),
.C(n_1402),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1651),
.B(n_1525),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1655),
.A2(n_1475),
.B1(n_1535),
.B2(n_1515),
.Y(n_1660)
);

NAND4xp25_ASAP7_75t_SL g1661 ( 
.A(n_1652),
.B(n_1531),
.C(n_1543),
.D(n_1510),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1656),
.A2(n_1475),
.B1(n_1526),
.B2(n_1538),
.Y(n_1662)
);

NAND4xp75_ASAP7_75t_L g1663 ( 
.A(n_1657),
.B(n_1531),
.C(n_1543),
.D(n_1537),
.Y(n_1663)
);

NAND4xp75_ASAP7_75t_L g1664 ( 
.A(n_1658),
.B(n_1531),
.C(n_1543),
.D(n_1537),
.Y(n_1664)
);

NOR2xp67_ASAP7_75t_L g1665 ( 
.A(n_1661),
.B(n_1526),
.Y(n_1665)
);

NOR2xp67_ASAP7_75t_L g1666 ( 
.A(n_1660),
.B(n_1659),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1666),
.Y(n_1667)
);

NOR2xp67_ASAP7_75t_L g1668 ( 
.A(n_1662),
.B(n_1665),
.Y(n_1668)
);

NAND3x1_ASAP7_75t_L g1669 ( 
.A(n_1663),
.B(n_1538),
.C(n_1548),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1667),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1670),
.A2(n_1668),
.B1(n_1664),
.B2(n_1669),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1671),
.B(n_1510),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1671),
.A2(n_1537),
.B1(n_1510),
.B2(n_1321),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_R g1674 ( 
.A(n_1672),
.B(n_1384),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1673),
.A2(n_1546),
.B1(n_1478),
.B2(n_1486),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1675),
.A2(n_1478),
.B1(n_1486),
.B2(n_1494),
.Y(n_1676)
);

OR2x6_ASAP7_75t_L g1677 ( 
.A(n_1674),
.B(n_1309),
.Y(n_1677)
);

AOI22x1_ASAP7_75t_L g1678 ( 
.A1(n_1677),
.A2(n_1298),
.B1(n_1375),
.B2(n_1379),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1676),
.B(n_1310),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1298),
.B1(n_1385),
.B2(n_1494),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1680),
.A2(n_1485),
.B1(n_1504),
.B2(n_1298),
.C(n_1486),
.Y(n_1681)
);

AOI211xp5_ASAP7_75t_L g1682 ( 
.A1(n_1681),
.A2(n_1385),
.B(n_1418),
.C(n_1485),
.Y(n_1682)
);


endmodule