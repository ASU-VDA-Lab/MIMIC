module real_jpeg_5656_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_0),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_0),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_0),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_0),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_0),
.B(n_209),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_0),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_0),
.B(n_295),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_1),
.Y(n_214)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_1),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_1),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_1),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_2),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_3),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_4),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_4),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_4),
.B(n_214),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_4),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_4),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_4),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_4),
.B(n_187),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_5),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_5),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_80),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_5),
.B(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_6),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_6),
.Y(n_120)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_7),
.Y(n_486)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_8),
.Y(n_216)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_8),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_8),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_9),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_9),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_39),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_9),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_9),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_9),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_9),
.B(n_404),
.Y(n_403)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_11),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_11),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_11),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_11),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_11),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_11),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_11),
.B(n_398),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_12),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_12),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_13),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_13),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_13),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_13),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_13),
.B(n_77),
.Y(n_132)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_15),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_15),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_15),
.B(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_15),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_15),
.B(n_44),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_15),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_15),
.B(n_387),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_16),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_16),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_16),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_16),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_16),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_16),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_16),
.B(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_16),
.B(n_344),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_17),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_17),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_17),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_17),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_18),
.B(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_18),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_18),
.B(n_56),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_18),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_18),
.B(n_308),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_18),
.B(n_344),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_18),
.B(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_18),
.B(n_395),
.Y(n_394)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_485),
.B(n_487),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_176),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_175),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_138),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_25),
.B(n_138),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_100),
.B2(n_137),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_69),
.C(n_83),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_28),
.B(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_47),
.C(n_54),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_29),
.A2(n_30),
.B1(n_47),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_31),
.B(n_36),
.C(n_43),
.Y(n_114)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_43),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_42),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_42),
.Y(n_377)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_42),
.Y(n_395)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_46),
.Y(n_168)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_46),
.Y(n_322)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_46),
.Y(n_399)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_47),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.C(n_53),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_48),
.B(n_53),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_49),
.B(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_52),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_54),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_62),
.C(n_65),
.Y(n_113)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_59),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_68),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_62),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_104),
.C(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_86),
.C(n_90),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_65),
.A2(n_68),
.B1(n_90),
.B2(n_91),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_67),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_69),
.A2(n_83),
.B1(n_84),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_75),
.C(n_82),
.Y(n_122)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_82),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_77),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_78),
.Y(n_342)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_81),
.Y(n_220)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_93),
.C(n_96),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_85),
.B(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_86),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_89),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_90),
.A2(n_91),
.B1(n_150),
.B2(n_200),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_149),
.C(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_96),
.A2(n_97),
.B1(n_170),
.B2(n_171),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_159),
.C(n_170),
.Y(n_158)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_99),
.Y(n_388)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_115),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.C(n_114),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_102),
.B(n_113),
.CI(n_114),
.CON(n_143),
.SN(n_143)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_105),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_110),
.Y(n_248)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_123),
.B2(n_136),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_134),
.B2(n_135),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_144),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_143),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g492 ( 
.A(n_143),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_144),
.B(n_480),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_156),
.C(n_158),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_145),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_154),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_146),
.B(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_148),
.B(n_154),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_199),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_152),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_153),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_156),
.B(n_158),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_169),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_169),
.Y(n_183)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_183),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_168),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_168),
.Y(n_370)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

AO21x1_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_477),
.B(n_483),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_278),
.B(n_476),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_227),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_179),
.B(n_227),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_221),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_180),
.B(n_222),
.C(n_225),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_201),
.C(n_203),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_181),
.B(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_198),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_182),
.B(n_462),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_184),
.A2(n_185),
.B1(n_198),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_194),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_186),
.B(n_194),
.Y(n_452)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_189),
.B(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_198),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_203),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_215),
.C(n_217),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_204),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_212),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_212),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_214),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_217),
.Y(n_256)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_220),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.C(n_234),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_229),
.B(n_232),
.Y(n_472)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_234),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_254),
.C(n_257),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_236),
.B(n_465),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.C(n_245),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_237),
.A2(n_238),
.B1(n_443),
.B2(n_444),
.Y(n_442)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_240),
.A2(n_241),
.B(n_244),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_240),
.B(n_245),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.C(n_251),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_420)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_251),
.B(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_252),
.B(n_355),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_257),
.Y(n_466)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_269),
.C(n_274),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_259),
.B(n_454),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.C(n_266),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_260),
.B(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_262),
.A2(n_266),
.B1(n_267),
.B2(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_262),
.Y(n_433)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_265),
.Y(n_298)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_269),
.B(n_274),
.Y(n_454)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_470),
.B(n_475),
.Y(n_278)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_457),
.B(n_469),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_439),
.B(n_456),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_413),
.B(n_438),
.Y(n_281)
);

AOI21x1_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_381),
.B(n_412),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_347),
.B(n_380),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_324),
.B(n_346),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_302),
.B(n_323),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_299),
.B(n_301),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_297),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_297),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

INVx3_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_304),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_312),
.B2(n_313),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_315),
.C(n_319),
.Y(n_345)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_310),
.Y(n_335)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_311),
.Y(n_334)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_319),
.B2(n_320),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_318),
.Y(n_356)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_345),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_345),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_336),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_335),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_335),
.C(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_332),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_366),
.C(n_367),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_339),
.Y(n_366)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_343),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_348),
.B(n_350),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_364),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_351),
.B(n_365),
.C(n_368),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_352),
.B(n_354),
.C(n_357),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_360),
.B1(n_361),
.B2(n_363),
.Y(n_357)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_358),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_363),
.Y(n_390)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

MAJx2_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_375),
.C(n_378),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_375),
.B1(n_378),
.B2(n_379),
.Y(n_371)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_372),
.Y(n_378)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_375),
.Y(n_379)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_411),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_411),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_392),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_391),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_384),
.B(n_391),
.C(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_390),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_389),
.Y(n_385)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_390),
.B(n_427),
.C(n_428),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_392),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_400),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_402),
.C(n_409),
.Y(n_416)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_393),
.Y(n_493)
);

FAx1_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_396),
.CI(n_397),
.CON(n_393),
.SN(n_393)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_396),
.C(n_397),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_402),
.B1(n_409),
.B2(n_410),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_408),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_408),
.Y(n_423)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_436),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_436),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_425),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_416),
.B(n_417),
.C(n_425),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_421),
.B2(n_422),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_448),
.C(n_449),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_424),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_429),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_430),
.C(n_435),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_431),
.B1(n_434),
.B2(n_435),
.Y(n_429)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_430),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_431),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_455),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_455),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_446),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_445),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_445),
.C(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_443),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_451),
.C(n_453),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_453),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_467),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_467),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_459),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_464),
.C(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_473),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_479),
.B(n_482),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx8_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx13_ASAP7_75t_L g489 ( 
.A(n_486),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_490),
.Y(n_487)
);

BUFx12f_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);


endmodule