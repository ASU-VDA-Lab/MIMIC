module fake_netlist_1_6993_n_530 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_530);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_530;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_73;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_388;
wire n_139;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g70 ( .A(n_69), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_41), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_16), .Y(n_72) );
CKINVDCx5p33_ASAP7_75t_R g73 ( .A(n_54), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_67), .Y(n_74) );
INVx2_ASAP7_75t_L g75 ( .A(n_10), .Y(n_75) );
CKINVDCx16_ASAP7_75t_R g76 ( .A(n_40), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_4), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_65), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_3), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_14), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_22), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_30), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_26), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_60), .Y(n_84) );
BUFx3_ASAP7_75t_L g85 ( .A(n_42), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_33), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_39), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_53), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_50), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_66), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_48), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_52), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_51), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_29), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_34), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_57), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_47), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_38), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_62), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_59), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_55), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_43), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_1), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_15), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_9), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_49), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_58), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_3), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_44), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_20), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_19), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_10), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_4), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_19), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_61), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_37), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_35), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_15), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_111), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_111), .Y(n_121) );
XOR2xp5_ASAP7_75t_L g122 ( .A(n_105), .B(n_0), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_111), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_83), .B(n_0), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_76), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_76), .B(n_1), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_71), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_93), .B(n_103), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_71), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_107), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_72), .Y(n_135) );
AND2x6_ASAP7_75t_L g136 ( .A(n_107), .B(n_27), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_74), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_107), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_115), .Y(n_140) );
BUFx8_ASAP7_75t_L g141 ( .A(n_117), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_93), .A2(n_2), .B1(n_5), .B2(n_6), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_103), .B(n_2), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_74), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_117), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_78), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_117), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_75), .B(n_5), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_78), .Y(n_149) );
INVx1_ASAP7_75t_SL g150 ( .A(n_90), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_70), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_82), .B(n_6), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_75), .B(n_7), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_82), .B(n_7), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_118), .B(n_31), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_119), .B(n_8), .Y(n_157) );
BUFx8_ASAP7_75t_L g158 ( .A(n_84), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_84), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_86), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_119), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_86), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_89), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_89), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_94), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_148), .A2(n_97), .B1(n_114), .B2(n_113), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_124), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_148), .B(n_72), .Y(n_168) );
INVxp67_ASAP7_75t_L g169 ( .A(n_150), .Y(n_169) );
AO22x2_ASAP7_75t_L g170 ( .A1(n_142), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_141), .Y(n_171) );
NAND3xp33_ASAP7_75t_L g172 ( .A(n_158), .B(n_104), .C(n_114), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_130), .B(n_73), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_130), .B(n_77), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_135), .B(n_77), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_126), .A2(n_79), .B1(n_113), .B2(n_112), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_124), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_153), .B(n_79), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_124), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_128), .B(n_92), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_129), .Y(n_189) );
AND2x6_ASAP7_75t_L g190 ( .A(n_157), .B(n_98), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_129), .Y(n_191) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_156), .B(n_91), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
INVx1_ASAP7_75t_SL g194 ( .A(n_127), .Y(n_194) );
AO22x2_ASAP7_75t_L g195 ( .A1(n_122), .A2(n_101), .B1(n_95), .B2(n_110), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_157), .B(n_80), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_161), .B(n_80), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_129), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_129), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_136), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_128), .B(n_96), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_131), .B(n_99), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_123), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_129), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_159), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_136), .Y(n_207) );
INVx4_ASAP7_75t_SL g208 ( .A(n_156), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_165), .B(n_106), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_127), .Y(n_210) );
INVxp33_ASAP7_75t_L g211 ( .A(n_143), .Y(n_211) );
AO21x2_ASAP7_75t_L g212 ( .A1(n_152), .A2(n_99), .B(n_110), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_132), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_159), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_143), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_162), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_136), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_131), .B(n_102), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_123), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_125), .B(n_97), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_137), .B(n_81), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_132), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_137), .B(n_106), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g225 ( .A1(n_158), .A2(n_104), .B1(n_112), .B2(n_109), .Y(n_225) );
INVxp33_ASAP7_75t_L g226 ( .A(n_122), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_204), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_185), .Y(n_228) );
AND2x6_ASAP7_75t_SL g229 ( .A(n_226), .B(n_154), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_185), .Y(n_230) );
INVxp67_ASAP7_75t_L g231 ( .A(n_169), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_185), .Y(n_232) );
CKINVDCx6p67_ASAP7_75t_R g233 ( .A(n_221), .Y(n_233) );
AND3x1_ASAP7_75t_SL g234 ( .A(n_195), .B(n_165), .C(n_149), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_206), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_214), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_204), .Y(n_237) );
BUFx3_ASAP7_75t_L g238 ( .A(n_171), .Y(n_238) );
INVx5_ASAP7_75t_L g239 ( .A(n_190), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_186), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
BUFx4f_ASAP7_75t_L g242 ( .A(n_190), .Y(n_242) );
AND2x4_ASAP7_75t_SL g243 ( .A(n_221), .B(n_158), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_220), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_171), .B(n_151), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_215), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_217), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_179), .B(n_141), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_174), .B(n_144), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_201), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
BUFx8_ASAP7_75t_L g253 ( .A(n_210), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_190), .Y(n_255) );
BUFx8_ASAP7_75t_SL g256 ( .A(n_216), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_190), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_190), .A2(n_136), .B1(n_141), .B2(n_156), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_187), .B(n_141), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_219), .B(n_146), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_190), .A2(n_136), .B1(n_156), .B2(n_149), .Y(n_261) );
OR2x6_ASAP7_75t_L g262 ( .A(n_221), .B(n_144), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_224), .B(n_146), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_222), .B(n_123), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_209), .B(n_123), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_177), .Y(n_266) );
NAND2x1p5_ASAP7_75t_L g267 ( .A(n_173), .B(n_164), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_209), .B(n_156), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_209), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_221), .Y(n_270) );
BUFx12f_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_198), .B(n_156), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_198), .B(n_156), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_168), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_168), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_194), .B(n_133), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_178), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_183), .A2(n_121), .B1(n_120), .B2(n_145), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_173), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_167), .Y(n_280) );
BUFx4f_ASAP7_75t_L g281 ( .A(n_207), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_225), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_173), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_182), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_188), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_207), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_183), .B(n_88), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_193), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_263), .B(n_211), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
BUFx4f_ASAP7_75t_L g291 ( .A(n_262), .Y(n_291) );
BUFx10_ASAP7_75t_L g292 ( .A(n_243), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_263), .B(n_211), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_269), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_240), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_271), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_269), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_240), .B(n_224), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_271), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_262), .B(n_175), .Y(n_300) );
AOI21x1_ASAP7_75t_L g301 ( .A1(n_268), .A2(n_203), .B(n_202), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_250), .B(n_175), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
INVx3_ASAP7_75t_SL g304 ( .A(n_233), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_262), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_228), .Y(n_306) );
NOR2xp67_ASAP7_75t_L g307 ( .A(n_231), .B(n_180), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_262), .Y(n_308) );
INVx4_ASAP7_75t_L g309 ( .A(n_242), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_270), .B(n_196), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_256), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_239), .B(n_196), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_242), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_244), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_228), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_243), .B(n_195), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_248), .B(n_270), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_253), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_253), .Y(n_319) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_254), .A2(n_197), .B(n_172), .C(n_166), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_238), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_244), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_253), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_272), .A2(n_192), .B(n_196), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_275), .B(n_197), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_241), .Y(n_326) );
INVx4_ASAP7_75t_L g327 ( .A(n_242), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_275), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_233), .A2(n_170), .B1(n_195), .B2(n_192), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_230), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_254), .A2(n_170), .B1(n_202), .B2(n_203), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_282), .A2(n_170), .B1(n_195), .B2(n_212), .Y(n_332) );
INVx5_ASAP7_75t_L g333 ( .A(n_239), .Y(n_333) );
AOI22xp33_ASAP7_75t_SL g334 ( .A1(n_238), .A2(n_207), .B1(n_218), .B2(n_212), .Y(n_334) );
INVxp67_ASAP7_75t_L g335 ( .A(n_276), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_273), .A2(n_218), .B(n_212), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_230), .Y(n_337) );
O2A1O1Ixp33_ASAP7_75t_SL g338 ( .A1(n_259), .A2(n_191), .B(n_223), .C(n_184), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_241), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_244), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_316), .A2(n_288), .B1(n_266), .B2(n_277), .Y(n_341) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_316), .A2(n_234), .B1(n_276), .B2(n_287), .Y(n_342) );
INVx3_ASAP7_75t_SL g343 ( .A(n_292), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_291), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_291), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_304), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_306), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_311), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_300), .A2(n_285), .B1(n_284), .B2(n_277), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_336), .A2(n_267), .B(n_261), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_291), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_335), .B(n_260), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_324), .A2(n_267), .B(n_264), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_306), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_304), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_329), .A2(n_239), .B1(n_235), .B2(n_236), .Y(n_356) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_332), .A2(n_239), .B1(n_235), .B2(n_236), .Y(n_357) );
INVx4_ASAP7_75t_L g358 ( .A(n_292), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_318), .A2(n_239), .B1(n_247), .B2(n_246), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_295), .A2(n_284), .B1(n_232), .B2(n_245), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_292), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_305), .A2(n_258), .B1(n_278), .B2(n_247), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_315), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_330), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_337), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_298), .B(n_289), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_320), .A2(n_232), .B(n_265), .C(n_255), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_298), .B(n_252), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_333), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_293), .B(n_302), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_333), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_308), .B(n_255), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_371), .B(n_293), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_345), .B(n_333), .Y(n_375) );
AOI22xp33_ASAP7_75t_SL g376 ( .A1(n_344), .A2(n_323), .B1(n_319), .B2(n_317), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_349), .A2(n_331), .B1(n_310), .B2(n_320), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g378 ( .A1(n_352), .A2(n_307), .B1(n_296), .B2(n_299), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_341), .A2(n_321), .B1(n_325), .B2(n_334), .Y(n_379) );
INVx11_ASAP7_75t_L g380 ( .A(n_348), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_321), .B1(n_309), .B2(n_313), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_367), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g383 ( .A1(n_344), .A2(n_309), .B1(n_313), .B2(n_327), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_371), .A2(n_290), .B1(n_294), .B2(n_297), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_342), .B(n_164), .C(n_163), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_366), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_343), .B(n_351), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_357), .A2(n_338), .B(n_301), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_356), .A2(n_303), .B1(n_328), .B2(n_340), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_351), .A2(n_257), .B1(n_255), .B2(n_314), .Y(n_391) );
OAI211xp5_ASAP7_75t_SL g392 ( .A1(n_361), .A2(n_133), .B(n_138), .C(n_229), .Y(n_392) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_345), .A2(n_313), .B1(n_327), .B2(n_309), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_347), .A2(n_322), .B1(n_327), .B2(n_257), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_369), .A2(n_252), .B1(n_218), .B2(n_257), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_369), .A2(n_138), .B(n_100), .C(n_338), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_279), .B1(n_283), .B2(n_252), .Y(n_397) );
OAI21xp33_ASAP7_75t_L g398 ( .A1(n_368), .A2(n_145), .B(n_147), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_353), .A2(n_326), .B(n_339), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_386), .Y(n_400) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_392), .B(n_362), .C(n_116), .D(n_108), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_376), .A2(n_354), .B1(n_364), .B2(n_360), .Y(n_402) );
AND2x2_ASAP7_75t_SL g403 ( .A(n_390), .B(n_358), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_387), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_389), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_392), .A2(n_365), .B1(n_363), .B2(n_373), .Y(n_406) );
AOI222xp33_ASAP7_75t_L g407 ( .A1(n_374), .A2(n_343), .B1(n_360), .B2(n_364), .C1(n_346), .C2(n_355), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_376), .A2(n_365), .B1(n_343), .B2(n_358), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_382), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_389), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_388), .B(n_370), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_375), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_379), .A2(n_359), .B1(n_355), .B2(n_346), .Y(n_413) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_384), .A2(n_385), .B1(n_377), .B2(n_396), .C(n_393), .Y(n_414) );
OA21x2_ASAP7_75t_L g415 ( .A1(n_399), .A2(n_350), .B(n_353), .Y(n_415) );
OAI31xp33_ASAP7_75t_SL g416 ( .A1(n_378), .A2(n_373), .A3(n_350), .B(n_139), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_398), .A2(n_160), .B1(n_164), .B2(n_163), .C(n_155), .Y(n_417) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_381), .A2(n_372), .B(n_370), .C(n_160), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_375), .B(n_372), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_393), .B(n_333), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_394), .B(n_160), .C(n_163), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_383), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_391), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_395), .B(n_333), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_376), .B(n_326), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g428 ( .A1(n_376), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_404), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_404), .Y(n_431) );
OAI33xp33_ASAP7_75t_L g432 ( .A1(n_428), .A2(n_200), .A3(n_205), .B1(n_213), .B2(n_223), .B3(n_199), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_409), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_400), .B(n_11), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_405), .A2(n_189), .B(n_199), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_411), .B(n_12), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_415), .Y(n_437) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_407), .A2(n_134), .B(n_155), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_401), .A2(n_134), .B1(n_155), .B2(n_237), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_412), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_423), .B(n_68), .Y(n_441) );
NAND2x1_ASAP7_75t_L g442 ( .A(n_429), .B(n_339), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_408), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_419), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_403), .A2(n_134), .B1(n_227), .B2(n_237), .Y(n_445) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_405), .A2(n_227), .B(n_312), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_426), .B(n_402), .Y(n_447) );
OR2x6_ASAP7_75t_L g448 ( .A(n_427), .B(n_339), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_429), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_403), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_424), .B(n_134), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_410), .B(n_16), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_406), .B(n_17), .Y(n_453) );
NOR2x1_ASAP7_75t_L g454 ( .A(n_413), .B(n_181), .Y(n_454) );
XNOR2xp5_ASAP7_75t_L g455 ( .A(n_420), .B(n_17), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_421), .B(n_64), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_416), .B(n_18), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_425), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_414), .A2(n_218), .B1(n_312), .B2(n_267), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_433), .Y(n_461) );
OAI33xp33_ASAP7_75t_L g462 ( .A1(n_430), .A2(n_431), .A3(n_444), .B1(n_458), .B2(n_443), .B3(n_453), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_436), .B(n_422), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_434), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_434), .Y(n_465) );
NOR2x1p5_ASAP7_75t_L g466 ( .A(n_441), .B(n_181), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_SL g467 ( .A1(n_438), .A2(n_417), .B(n_23), .C(n_24), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_459), .B(n_181), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_440), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_453), .B(n_21), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_452), .Y(n_471) );
AND2x2_ASAP7_75t_SL g472 ( .A(n_441), .B(n_281), .Y(n_472) );
OAI22xp5_ASAP7_75t_SL g473 ( .A1(n_455), .A2(n_25), .B1(n_28), .B2(n_32), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_449), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_457), .B(n_36), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_447), .B(n_45), .Y(n_476) );
INVxp33_ASAP7_75t_SL g477 ( .A(n_454), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_450), .B(n_46), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_451), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_456), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_448), .B(n_56), .Y(n_481) );
OAI31xp33_ASAP7_75t_L g482 ( .A1(n_473), .A2(n_456), .A3(n_439), .B(n_445), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_464), .B(n_448), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_465), .B(n_448), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_479), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_461), .Y(n_486) );
NAND2x1p5_ASAP7_75t_L g487 ( .A(n_466), .B(n_442), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_474), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_471), .B(n_437), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_462), .A2(n_432), .B1(n_460), .B2(n_446), .Y(n_490) );
NAND2x1p5_ASAP7_75t_L g491 ( .A(n_481), .B(n_442), .Y(n_491) );
AOI21xp33_ASAP7_75t_SL g492 ( .A1(n_477), .A2(n_435), .B(n_63), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_469), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_467), .A2(n_281), .B(n_279), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_463), .B(n_280), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_472), .A2(n_281), .B1(n_208), .B2(n_249), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_468), .B(n_208), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_476), .B(n_251), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_486), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_488), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_492), .A2(n_467), .B(n_470), .C(n_475), .Y(n_501) );
NAND4xp25_ASAP7_75t_L g502 ( .A(n_482), .B(n_483), .C(n_484), .D(n_490), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_485), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_495), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_489), .B(n_478), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_491), .A2(n_286), .B1(n_487), .B2(n_490), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_498), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_497), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_497), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_494), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_496), .A2(n_466), .B1(n_438), .B2(n_480), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_493), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_486), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_486), .Y(n_514) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_511), .B(n_502), .C(n_501), .D(n_506), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_512), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_503), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_506), .A2(n_504), .B1(n_510), .B2(n_505), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_515), .A2(n_499), .B1(n_500), .B2(n_514), .C(n_513), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_516), .Y(n_520) );
OAI211xp5_ASAP7_75t_L g521 ( .A1(n_518), .A2(n_507), .B(n_509), .C(n_508), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_517), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_520), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_522), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_523), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_525), .B(n_519), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_526), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_527), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_528), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_529), .A2(n_524), .B(n_521), .Y(n_530) );
endmodule