module fake_jpeg_23695_n_222 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_9),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_35),
.B(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

OR2x4_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_32),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_21),
.Y(n_51)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_60),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_32),
.B1(n_21),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_18),
.B1(n_17),
.B2(n_4),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_51),
.B(n_55),
.Y(n_89)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_31),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_33),
.B1(n_25),
.B2(n_30),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_68),
.B1(n_18),
.B2(n_17),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_23),
.B(n_28),
.C(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_67),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

OR2x2_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_71),
.Y(n_96)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_36),
.A2(n_33),
.B1(n_25),
.B2(n_27),
.Y(n_68)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_45),
.B1(n_40),
.B2(n_38),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_33),
.B1(n_19),
.B2(n_26),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_16),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_90),
.B(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_39),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_8),
.B(n_9),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_36),
.B1(n_41),
.B2(n_22),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_83),
.B1(n_80),
.B2(n_73),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_19),
.B1(n_22),
.B2(n_41),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_92),
.B1(n_99),
.B2(n_70),
.Y(n_108)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_94),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_55),
.B1(n_56),
.B2(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_3),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g121 ( 
.A(n_91),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_18),
.B1(n_17),
.B2(n_4),
.Y(n_92)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_97),
.Y(n_106)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_52),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_3),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_107),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_102),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_91),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_47),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_110),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_12),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_66),
.B1(n_57),
.B2(n_62),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_112),
.B1(n_117),
.B2(n_128),
.Y(n_150)
);

OAI22x1_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_62),
.B1(n_6),
.B2(n_7),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_119),
.B(n_96),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_74),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_123),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_7),
.B(n_8),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_84),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_9),
.B(n_10),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_14),
.Y(n_127)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_84),
.B1(n_96),
.B2(n_101),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_137),
.Y(n_158)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_152),
.B1(n_112),
.B2(n_116),
.C(n_111),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_118),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_99),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_108),
.C(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_141),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_142),
.B(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_85),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_100),
.B(n_86),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_86),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_82),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_97),
.B(n_98),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_160),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_115),
.B1(n_126),
.B2(n_120),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_170),
.C(n_164),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_105),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_165),
.Y(n_174)
);

NOR2x1p5_ASAP7_75t_SL g164 ( 
.A(n_131),
.B(n_117),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_152),
.B(n_132),
.C(n_148),
.D(n_141),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_121),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_104),
.C(n_106),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_142),
.B(n_139),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_169),
.B1(n_171),
.B2(n_168),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_144),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_179),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_178),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_150),
.C(n_132),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_168),
.B1(n_164),
.B2(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_186),
.A2(n_173),
.B1(n_162),
.B2(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_193),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_195),
.B1(n_179),
.B2(n_175),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_155),
.B1(n_162),
.B2(n_152),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_197),
.A2(n_201),
.B(n_195),
.C(n_190),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_135),
.B(n_153),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_200),
.B(n_130),
.Y(n_209)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_170),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_172),
.C(n_188),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.C(n_172),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_140),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_210),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_188),
.C(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_207),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_181),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_167),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_136),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_213),
.A2(n_198),
.B1(n_201),
.B2(n_196),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_212),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_217),
.B(n_110),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_104),
.C(n_136),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_219),
.A3(n_202),
.B1(n_146),
.B2(n_140),
.C1(n_145),
.C2(n_94),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_146),
.C(n_121),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_91),
.Y(n_222)
);


endmodule