module fake_jpeg_20561_n_237 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_114;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_24),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_20),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_25),
.B(n_29),
.Y(n_58)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_28),
.B1(n_21),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_47),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_44),
.C(n_45),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_49),
.C(n_8),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_44),
.C(n_20),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_19),
.B1(n_21),
.B2(n_28),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_26),
.B1(n_32),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_26),
.B1(n_32),
.B2(n_27),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_57),
.B1(n_75),
.B2(n_4),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_18),
.B1(n_16),
.B2(n_3),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_18),
.B1(n_16),
.B2(n_29),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_58),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_59),
.B(n_79),
.Y(n_108)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_30),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_34),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_40),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_34),
.B(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_81),
.B(n_8),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_5),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_5),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_48),
.B(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_6),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_7),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_97),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_70),
.Y(n_119)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_99),
.Y(n_113)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_64),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_59),
.C(n_70),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_119),
.C(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_50),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_124),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_74),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_107),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_123),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_136),
.B(n_134),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_59),
.B(n_9),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_137),
.B(n_11),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_73),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_86),
.B(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_9),
.B(n_10),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_11),
.B(n_107),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_133),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_65),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_67),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_77),
.Y(n_160)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_63),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_95),
.B(n_9),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_85),
.B1(n_90),
.B2(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_148),
.B1(n_157),
.B2(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_130),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_103),
.C(n_12),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_101),
.B1(n_93),
.B2(n_76),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_156),
.Y(n_165)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_162),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_153),
.C(n_159),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_93),
.B1(n_106),
.B2(n_109),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_99),
.B1(n_89),
.B2(n_82),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_119),
.A2(n_98),
.B1(n_82),
.B2(n_89),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_174),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_132),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_112),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_128),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_110),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_181),
.Y(n_183)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_117),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_117),
.B(n_146),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_141),
.C(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_111),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_184),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_180),
.A2(n_162),
.B1(n_145),
.B2(n_156),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_160),
.C(n_148),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_190),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_151),
.B1(n_157),
.B2(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_187),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_163),
.B1(n_110),
.B2(n_142),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_164),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_133),
.C(n_142),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_195),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_174),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_SL g196 ( 
.A(n_175),
.B(n_116),
.C(n_124),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_169),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_172),
.B1(n_179),
.B2(n_170),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_199),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_179),
.B1(n_173),
.B2(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_201),
.A2(n_202),
.B1(n_167),
.B2(n_164),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_137),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_173),
.B1(n_168),
.B2(n_171),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_206),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_204),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_213),
.C(n_139),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_210),
.B(n_212),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_214),
.B(n_113),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_196),
.C(n_125),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_182),
.C(n_185),
.Y(n_213)
);

OAI21x1_ASAP7_75t_SL g214 ( 
.A1(n_200),
.A2(n_191),
.B(n_150),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_208),
.B(n_199),
.C(n_198),
.Y(n_218)
);

AOI221xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_223),
.B1(n_211),
.B2(n_123),
.C(n_118),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_220),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_204),
.B1(n_158),
.B2(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_224),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_154),
.C(n_139),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_215),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_228),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_135),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_229),
.B(n_227),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_114),
.C(n_131),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_223),
.C(n_120),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_120),
.C(n_114),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_231),
.C(n_84),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_61),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);


endmodule