module fake_jpeg_24044_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

AND2x2_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_4),
.Y(n_10)
);

AND2x2_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_7),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_20),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_1),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_22),
.B(n_11),
.C(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_2),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_16),
.B1(n_11),
.B2(n_14),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_10),
.B1(n_23),
.B2(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_11),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_36),
.C(n_38),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_10),
.B1(n_27),
.B2(n_14),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_18),
.C(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_18),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_26),
.C(n_30),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.C(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_33),
.B1(n_40),
.B2(n_39),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_44),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_39),
.C(n_46),
.Y(n_53)
);

XNOR2x2_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_50),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

OAI21x1_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_54),
.B(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_2),
.Y(n_58)
);


endmodule