module fake_jpeg_21426_n_346 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_45),
.Y(n_56)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_16),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_16),
.B1(n_17),
.B2(n_29),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_64),
.A2(n_38),
.B1(n_36),
.B2(n_41),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_50),
.B1(n_17),
.B2(n_29),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_70),
.A2(n_84),
.B1(n_100),
.B2(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_72),
.B(n_75),
.Y(n_124)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_15),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_79),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_80),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_83),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_54),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_49),
.B1(n_46),
.B2(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_15),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_85),
.Y(n_141)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_98),
.B1(n_108),
.B2(n_91),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_89),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_28),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_28),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_94),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_32),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_102),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_17),
.B1(n_46),
.B2(n_59),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_65),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_37),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_38),
.B1(n_36),
.B2(n_42),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_63),
.B(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_107),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_43),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_52),
.A2(n_48),
.B1(n_44),
.B2(n_25),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_68),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_47),
.B1(n_43),
.B2(n_34),
.Y(n_142)
);

BUFx2_ASAP7_75t_SL g110 ( 
.A(n_52),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_40),
.B1(n_37),
.B2(n_25),
.Y(n_127)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_43),
.C(n_40),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_43),
.C(n_111),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_78),
.B1(n_112),
.B2(n_71),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_75),
.A2(n_25),
.B1(n_35),
.B2(n_24),
.Y(n_138)
);

OAI22x1_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_30),
.B1(n_18),
.B2(n_84),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_136),
.B(n_124),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_150),
.B(n_24),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_72),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_148),
.B(n_156),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_73),
.B(n_105),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_131),
.B1(n_119),
.B2(n_115),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_151),
.A2(n_47),
.B(n_92),
.Y(n_203)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_81),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_169),
.Y(n_195)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_83),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_107),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_125),
.B(n_99),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_160),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

OAI22x1_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_87),
.B1(n_80),
.B2(n_143),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_165),
.Y(n_191)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_94),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_136),
.B1(n_102),
.B2(n_145),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_171),
.B1(n_134),
.B2(n_113),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_116),
.C(n_120),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_133),
.C(n_109),
.Y(n_178)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_77),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_184),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_R g177 ( 
.A(n_158),
.B(n_133),
.C(n_126),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_177),
.A2(n_183),
.B(n_207),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_179),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_106),
.C(n_104),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_139),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_18),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_186),
.B(n_47),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_193),
.B1(n_197),
.B2(n_166),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_149),
.A2(n_134),
.B1(n_86),
.B2(n_144),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_190),
.A2(n_192),
.B1(n_206),
.B2(n_152),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_149),
.A2(n_134),
.B1(n_144),
.B2(n_132),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_121),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_198),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_98),
.B1(n_121),
.B2(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_47),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_203),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_174),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_151),
.A2(n_88),
.B1(n_76),
.B2(n_93),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_SL g207 ( 
.A1(n_153),
.A2(n_30),
.B(n_18),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_215),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_181),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_153),
.B(n_164),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_228),
.B(n_234),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_220),
.B1(n_226),
.B2(n_192),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_184),
.A2(n_169),
.B1(n_173),
.B2(n_170),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_161),
.Y(n_221)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_224),
.B(n_227),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_198),
.Y(n_225)
);

AO22x1_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_230),
.B1(n_231),
.B2(n_194),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_157),
.B1(n_165),
.B2(n_172),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_155),
.C(n_30),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_175),
.A2(n_147),
.B(n_135),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_33),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_33),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_186),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_177),
.Y(n_233)
);

INVx13_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_203),
.A2(n_34),
.B(n_74),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_74),
.B(n_22),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_190),
.B(n_180),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_22),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_236),
.B(n_230),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_238),
.A2(n_242),
.B1(n_252),
.B2(n_256),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_195),
.C(n_179),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_248),
.C(n_221),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_260),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_250),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_195),
.C(n_178),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_222),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_213),
.A2(n_204),
.B1(n_182),
.B2(n_22),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_223),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_262),
.B(n_234),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_219),
.A2(n_182),
.B1(n_33),
.B2(n_3),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_209),
.A2(n_33),
.B1(n_2),
.B2(n_3),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_225),
.B1(n_208),
.B2(n_212),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_220),
.B(n_8),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_210),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_224),
.C(n_215),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_232),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_266),
.Y(n_291)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_268),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_251),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_272),
.Y(n_287)
);

AO22x1_ASAP7_75t_SL g270 ( 
.A1(n_240),
.A2(n_216),
.B1(n_209),
.B2(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_217),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_274),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_217),
.B(n_211),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_237),
.B1(n_257),
.B2(n_256),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_235),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_278),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_226),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_208),
.C(n_227),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_283),
.C(n_245),
.Y(n_288)
);

FAx1_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_1),
.CI(n_2),
.CON(n_282),
.SN(n_282)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_254),
.B(n_253),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_239),
.B(n_6),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_268),
.A2(n_237),
.B1(n_239),
.B2(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_247),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_288),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_1),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_293),
.B1(n_280),
.B2(n_270),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_264),
.B(n_257),
.Y(n_290)
);

XOR2x2_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_279),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_249),
.B1(n_244),
.B2(n_258),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_246),
.C(n_252),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_296),
.C(n_301),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_246),
.C(n_9),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_6),
.C(n_13),
.Y(n_301)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_305),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_294),
.Y(n_320)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_308),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_267),
.C(n_281),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_313),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_285),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_270),
.B1(n_282),
.B2(n_283),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_282),
.B1(n_9),
.B2(n_10),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_295),
.A2(n_14),
.B(n_13),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_314),
.A2(n_14),
.B(n_12),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_288),
.Y(n_316)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_316),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_307),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_324),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_303),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_323),
.B1(n_313),
.B2(n_296),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_291),
.C(n_300),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_304),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_329),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_315),
.B(n_306),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_303),
.C(n_300),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_328),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_332),
.B(n_334),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_327),
.B(n_322),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_333),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_326),
.C(n_294),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_337),
.A2(n_335),
.B(n_314),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_339),
.C(n_338),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_311),
.C(n_301),
.Y(n_342)
);

AOI322xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_290),
.A3(n_6),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_2),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_1),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_SL g345 ( 
.A1(n_344),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_4),
.C(n_5),
.Y(n_346)
);


endmodule