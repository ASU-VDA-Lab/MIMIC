module fake_jpeg_26621_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_25),
.Y(n_62)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_56),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_22),
.B1(n_34),
.B2(n_20),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_20),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_62),
.B(n_21),
.C(n_16),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_22),
.B1(n_16),
.B2(n_21),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_41),
.B1(n_36),
.B2(n_32),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_22),
.B1(n_40),
.B2(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_70),
.B1(n_96),
.B2(n_94),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_22),
.B1(n_40),
.B2(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_83),
.B1(n_33),
.B2(n_19),
.Y(n_117)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_62),
.Y(n_100)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_38),
.B1(n_36),
.B2(n_44),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_54),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_21),
.B1(n_26),
.B2(n_30),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_52),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_26),
.B1(n_30),
.B2(n_20),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_25),
.B1(n_19),
.B2(n_33),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_28),
.B1(n_29),
.B2(n_18),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_100),
.B(n_25),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_58),
.B1(n_64),
.B2(n_29),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_102),
.A2(n_117),
.B1(n_32),
.B2(n_18),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_110),
.B1(n_118),
.B2(n_67),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_64),
.B1(n_50),
.B2(n_57),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_50),
.B1(n_37),
.B2(n_54),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_44),
.B1(n_46),
.B2(n_45),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_126),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_121),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_27),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_74),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_149),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_72),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_148),
.B(n_101),
.Y(n_161)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_135),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_147),
.B1(n_24),
.B2(n_29),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_90),
.B1(n_85),
.B2(n_67),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_144),
.B1(n_124),
.B2(n_105),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_139),
.B(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_76),
.B1(n_86),
.B2(n_87),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_87),
.B1(n_89),
.B2(n_78),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_152),
.B1(n_153),
.B2(n_105),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_33),
.B1(n_32),
.B2(n_19),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_SL g148 ( 
.A(n_100),
.B(n_118),
.C(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_73),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_154),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_92),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_80),
.B1(n_46),
.B2(n_45),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_43),
.Y(n_154)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_101),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_159),
.B(n_164),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_161),
.A2(n_162),
.B(n_179),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_98),
.B(n_112),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_112),
.C(n_43),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_189),
.C(n_0),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_37),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_37),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_152),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_168),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_122),
.A3(n_125),
.B1(n_106),
.B2(n_111),
.C1(n_37),
.C2(n_27),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_123),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_172),
.B(n_183),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_28),
.B1(n_14),
.B2(n_13),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_178),
.B1(n_180),
.B2(n_187),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_111),
.B(n_122),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_135),
.B1(n_17),
.B2(n_28),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_133),
.A2(n_123),
.B1(n_125),
.B2(n_44),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_17),
.B(n_1),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_133),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_138),
.B(n_140),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_46),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_191),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_11),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_143),
.B(n_11),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_184),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_135),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_186),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_46),
.B1(n_45),
.B2(n_29),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_45),
.C(n_24),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_15),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_129),
.B(n_28),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_192),
.A2(n_207),
.B1(n_211),
.B2(n_9),
.Y(n_243)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_193),
.B(n_198),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_155),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_210),
.B(n_214),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_217),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_140),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_205),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_128),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_206),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_128),
.B1(n_156),
.B2(n_134),
.Y(n_207)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_218),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_160),
.A2(n_17),
.B(n_135),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_158),
.B(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_179),
.B(n_162),
.C(n_166),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_175),
.A2(n_12),
.B1(n_10),
.B2(n_2),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_169),
.B1(n_10),
.B2(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_158),
.B(n_12),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_187),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_222),
.B(n_164),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_224),
.B(n_234),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_208),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_189),
.C(n_174),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_232),
.C(n_233),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_197),
.B(n_188),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_231),
.B(n_219),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_170),
.C(n_180),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_170),
.C(n_177),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_178),
.B(n_186),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_171),
.CI(n_169),
.CON(n_238),
.SN(n_238)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_208),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_171),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_242),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_211),
.B1(n_219),
.B2(n_208),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_0),
.Y(n_242)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_200),
.B(n_0),
.C(n_1),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_195),
.C(n_202),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_220),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_245),
.B(n_215),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_225),
.A2(n_194),
.B1(n_193),
.B2(n_214),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_249),
.A2(n_269),
.B1(n_241),
.B2(n_247),
.Y(n_271)
);

XOR2x2_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_194),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_250),
.A2(n_254),
.B(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_235),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_258),
.B(n_261),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_226),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_247),
.A2(n_213),
.B(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_203),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_263),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_202),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_268),
.Y(n_276)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_267),
.A2(n_261),
.B1(n_250),
.B2(n_259),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_233),
.C(n_232),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_272),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_249),
.B1(n_260),
.B2(n_257),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_228),
.C(n_230),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_265),
.B(n_224),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_273),
.B(n_258),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_265),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_1),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_266),
.B1(n_251),
.B2(n_259),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_228),
.C(n_234),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_284),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_244),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_248),
.C(n_237),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_242),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_229),
.C(n_199),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_196),
.Y(n_293)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_290),
.A2(n_298),
.B1(n_4),
.B2(n_5),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_253),
.C(n_260),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_293),
.Y(n_310)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_274),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_299),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_278),
.B1(n_282),
.B2(n_276),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_1),
.C(n_2),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_2),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_3),
.B(n_4),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_301),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_277),
.B1(n_274),
.B2(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_309),
.B(n_296),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_307),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_275),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_9),
.C(n_5),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_297),
.C(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_318),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_316),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_295),
.C(n_301),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_4),
.C(n_5),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_306),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_SL g320 ( 
.A(n_307),
.B(n_4),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_321),
.B(n_322),
.Y(n_324)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_305),
.A2(n_6),
.B(n_7),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_312),
.A2(n_6),
.B(n_7),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_313),
.B1(n_303),
.B2(n_302),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_328),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_311),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_304),
.Y(n_331)
);

OAI21x1_ASAP7_75t_SL g330 ( 
.A1(n_327),
.A2(n_317),
.B(n_313),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_330),
.B(n_331),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_326),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_329),
.B(n_327),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_324),
.B1(n_309),
.B2(n_9),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_6),
.B1(n_9),
.B2(n_257),
.Y(n_337)
);


endmodule