module fake_jpeg_21376_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_20),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_46),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_47),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_27),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_26),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_23),
.Y(n_67)
);

OR2x4_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_19),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_32),
.Y(n_72)
);

AOI32xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_22),
.A3(n_33),
.B1(n_39),
.B2(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_61),
.Y(n_94)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_72),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_24),
.B(n_30),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_SL g97 ( 
.A(n_66),
.B(n_67),
.C(n_84),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_74),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_22),
.B1(n_33),
.B2(n_31),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_85),
.B1(n_86),
.B2(n_25),
.Y(n_111)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

OA22x2_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_41),
.B1(n_36),
.B2(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_75),
.B(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_79),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_35),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_43),
.B(n_31),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_22),
.B1(n_17),
.B2(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_36),
.B1(n_25),
.B2(n_32),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_49),
.B1(n_36),
.B2(n_35),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_23),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_23),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_49),
.B1(n_54),
.B2(n_36),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_96),
.B1(n_108),
.B2(n_74),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_3),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_20),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_74),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_25),
.B1(n_18),
.B2(n_2),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_112),
.B(n_113),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_0),
.B(n_1),
.Y(n_112)
);

OR2x4_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_18),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_1),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_2),
.B(n_3),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_62),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_79),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_121),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_75),
.C(n_76),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_139),
.C(n_112),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_106),
.B1(n_110),
.B2(n_96),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_72),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_130),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_98),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_80),
.B1(n_87),
.B2(n_63),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_129),
.B1(n_103),
.B2(n_92),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_60),
.B1(n_70),
.B2(n_61),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_60),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_132),
.B(n_133),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_81),
.B(n_4),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_4),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_4),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_114),
.B(n_100),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_5),
.B(n_6),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_5),
.B(n_8),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_14),
.C(n_6),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_126),
.Y(n_172)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_159),
.B1(n_136),
.B2(n_127),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_160),
.B1(n_139),
.B2(n_131),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_114),
.B(n_113),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_149),
.B(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_151),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_105),
.B(n_92),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_106),
.C(n_97),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_102),
.C(n_97),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_121),
.C(n_124),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_122),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_102),
.B(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_104),
.B1(n_7),
.B2(n_8),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_167),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_169),
.B(n_144),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_127),
.B1(n_128),
.B2(n_125),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_172),
.C(n_175),
.Y(n_179)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_148),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_118),
.C(n_123),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_117),
.C(n_116),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_141),
.C(n_154),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_156),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_182),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_153),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_168),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_171),
.B1(n_169),
.B2(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_153),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_147),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_170),
.C(n_157),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_136),
.B1(n_141),
.B2(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_190),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_146),
.B1(n_154),
.B2(n_159),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_197),
.C(n_198),
.Y(n_202)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_196),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_200),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_185),
.B(n_184),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_161),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_157),
.C(n_145),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_160),
.B(n_147),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_178),
.C(n_164),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_191),
.B(n_180),
.CI(n_182),
.CON(n_204),
.SN(n_204)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_196),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_151),
.C(n_135),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_207),
.B(n_192),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_186),
.C(n_132),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.C(n_201),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_133),
.C(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_212),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_193),
.B(n_195),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_214),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_189),
.C(n_127),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_189),
.B1(n_205),
.B2(n_207),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_206),
.B(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_206),
.B(n_138),
.Y(n_220)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_221),
.A3(n_215),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_5),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_138),
.C(n_104),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_9),
.B(n_10),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_222),
.Y(n_225)
);


endmodule