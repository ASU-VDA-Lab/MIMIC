module real_jpeg_18662_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_0),
.A2(n_129),
.B1(n_134),
.B2(n_135),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_0),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_1),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_1),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_2),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_3),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_33),
.B1(n_95),
.B2(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_3),
.A2(n_33),
.B1(n_244),
.B2(n_269),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_3),
.A2(n_33),
.B1(n_305),
.B2(n_308),
.Y(n_304)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_4),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_5),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_5),
.A2(n_54),
.B1(n_85),
.B2(n_87),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_54),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_5),
.B(n_220),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g279 ( 
.A1(n_5),
.A2(n_280),
.A3(n_283),
.B1(n_286),
.B2(n_290),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_5),
.B(n_101),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_5),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_5),
.B(n_61),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_6),
.Y(n_90)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_6),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_6),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_7),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_7),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_7),
.A2(n_110),
.B1(n_197),
.B2(n_200),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_7),
.A2(n_110),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

BUFx4f_ASAP7_75t_L g150 ( 
.A(n_10),
.Y(n_150)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_10),
.Y(n_181)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_227),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_224),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_188),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_15),
.B(n_188),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_126),
.C(n_165),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_16),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_58),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_17),
.B(n_59),
.C(n_92),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_28),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_19),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_R g170 ( 
.A(n_20),
.B(n_54),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_20)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_21),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_22),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_28),
.B(n_38),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_30),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_32),
.Y(n_159)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_53),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_46),
.B2(n_50),
.Y(n_39)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_40),
.Y(n_211)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_54),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_54),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_54),
.B(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_56),
.A2(n_152),
.B1(n_155),
.B2(n_164),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_91),
.B2(n_92),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_72),
.B(n_84),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_61),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_61),
.B(n_84),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_61),
.B(n_268),
.Y(n_298)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_70),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_65),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_74),
.B1(n_77),
.B2(n_80),
.Y(n_73)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_72),
.B(n_84),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_72),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_72),
.B(n_196),
.Y(n_350)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_76),
.Y(n_203)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_83),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g255 ( 
.A(n_90),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x4_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_108),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_93),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_101),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_94),
.B(n_117),
.Y(n_169)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_101),
.B(n_109),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_101),
.B(n_218),
.Y(n_217)
);

AO22x2_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_117),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_113),
.Y(n_220)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_115),
.A2(n_119),
.B1(n_121),
.B2(n_124),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_117),
.Y(n_356)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_122),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_122),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_124),
.Y(n_240)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_126),
.A2(n_165),
.B1(n_166),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_126),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_151),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_127),
.B(n_151),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_136),
.B(n_139),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_128),
.A2(n_141),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_133),
.Y(n_285)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_138),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_139),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_141),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_141),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_144),
.Y(n_302)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_147),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_183),
.B(n_186),
.Y(n_182)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_171),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_167),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

AND2x4_ASAP7_75t_SL g216 ( 
.A(n_169),
.B(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_182),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_173),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_174),
.Y(n_262)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_177),
.Y(n_289)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_180),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_181),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_182),
.B(n_303),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_205),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_204),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_194),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_195),
.B(n_267),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2x1_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_223),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_215),
.B2(n_216),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_218),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_237),
.A3(n_241),
.B1(n_246),
.B2(n_250),
.Y(n_236)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_274),
.B(n_367),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_271),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_231),
.B(n_271),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.C(n_263),
.Y(n_231)
);

XOR2x1_ASAP7_75t_L g362 ( 
.A(n_232),
.B(n_363),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_235),
.A2(n_263),
.B1(n_264),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_235),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_256),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_236),
.A2(n_256),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_236),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_256),
.Y(n_358)
);

OA21x2_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_261),
.B(n_262),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_259),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_301),
.B(n_303),
.Y(n_300)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI21x1_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_361),
.B(n_366),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_342),
.B(n_360),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_317),
.B(n_341),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_299),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_278),
.B(n_299),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_297),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_297),
.Y(n_339)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_312),
.Y(n_299)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_315),
.C(n_344),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_336),
.B(n_340),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_332),
.B(n_335),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_328),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_334),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_339),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_345),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_357),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_351),
.B2(n_352),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_352),
.C(n_357),
.Y(n_365)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NOR2x1_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_365),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_362),
.B(n_365),
.Y(n_366)
);


endmodule