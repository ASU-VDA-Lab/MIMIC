module real_jpeg_6767_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_1),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_2),
.A2(n_59),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_2),
.A2(n_59),
.B1(n_177),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_2),
.A2(n_59),
.B1(n_120),
.B2(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_3),
.A2(n_81),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_3),
.B(n_142),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_3),
.B(n_196),
.C(n_340),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g343 ( 
.A1(n_3),
.A2(n_344),
.B1(n_345),
.B2(n_347),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_3),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_3),
.B(n_205),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_3),
.A2(n_86),
.B1(n_388),
.B2(n_391),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_69),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_4),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_4),
.A2(n_116),
.B1(n_272),
.B2(n_275),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_4),
.A2(n_116),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_4),
.A2(n_116),
.B1(n_372),
.B2(n_389),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_5),
.A2(n_134),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_5),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_5),
.A2(n_138),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_5),
.A2(n_138),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_5),
.A2(n_138),
.B1(n_186),
.B2(n_378),
.Y(n_377)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_7),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_7),
.Y(n_220)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_7),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_7),
.Y(n_288)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_7),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_10),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_10),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_10),
.A2(n_187),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_10),
.A2(n_187),
.B1(n_226),
.B2(n_229),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_10),
.A2(n_141),
.B1(n_187),
.B2(n_329),
.Y(n_328)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_11),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_11),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_11),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_12),
.A2(n_108),
.B1(n_176),
.B2(n_179),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_12),
.A2(n_108),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_13),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_13),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_14),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_14),
.A2(n_52),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_14),
.A2(n_52),
.B1(n_367),
.B2(n_369),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_14),
.A2(n_52),
.B1(n_422),
.B2(n_427),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_15),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_15),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_15),
.A2(n_98),
.B1(n_150),
.B2(n_153),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_15),
.A2(n_50),
.B1(n_98),
.B2(n_207),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_15),
.A2(n_70),
.B1(n_98),
.B2(n_214),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_456),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_331),
.B(n_450),
.Y(n_17)
);

NAND3xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_279),
.C(n_307),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_255),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_20),
.A2(n_452),
.B(n_453),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_230),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_21),
.B(n_230),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_144),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_22),
.B(n_145),
.C(n_199),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_64),
.C(n_111),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_23),
.B(n_111),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_48),
.B(n_56),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_24),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_24),
.B(n_206),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_24),
.A2(n_205),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_24),
.A2(n_205),
.B1(n_271),
.B2(n_419),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_24),
.A2(n_314),
.B(n_466),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_25),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_25),
.A2(n_203),
.B1(n_245),
.B2(n_253),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_25),
.A2(n_203),
.B1(n_245),
.B2(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_25),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_28),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_28),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_28),
.Y(n_426)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_29),
.Y(n_152)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_29),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_29),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_29),
.Y(n_346)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_29),
.Y(n_349)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_30),
.Y(n_411)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_32),
.Y(n_415)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_33),
.Y(n_180)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_33),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_38),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_39),
.Y(n_130)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_40),
.Y(n_274)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_48),
.Y(n_253)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_50),
.Y(n_207)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_57),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

INVx8_ASAP7_75t_L g407 ( 
.A(n_58),
.Y(n_407)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_63),
.Y(n_249)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_63),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_64),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_85),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_65),
.B(n_85),
.Y(n_258)
);

OAI32xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.A3(n_72),
.B1(n_76),
.B2(n_80),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g276 ( 
.A(n_68),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_71),
.Y(n_242)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_92),
.B1(n_102),
.B2(n_104),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_86),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_86),
.A2(n_104),
.B(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_86),
.A2(n_193),
.B(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_86),
.A2(n_191),
.B(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_86),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_86),
.A2(n_377),
.B1(n_388),
.B2(n_391),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_86),
.A2(n_193),
.B(n_219),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_89),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_91),
.Y(n_382)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_93),
.A2(n_184),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_94),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_95),
.Y(n_390)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_101),
.Y(n_378)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_110),
.Y(n_368)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_110),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_117),
.B1(n_132),
.B2(n_142),
.Y(n_111)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_112),
.Y(n_243)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_117),
.A2(n_301),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_117),
.B(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_118),
.A2(n_133),
.B1(n_143),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_118),
.A2(n_143),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_118),
.A2(n_210),
.B(n_300),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_127),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_119)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_120),
.Y(n_302)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_127),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_136),
.Y(n_329)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_142),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_143),
.B(n_328),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_143),
.A2(n_470),
.B(n_471),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_199),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_181),
.B2(n_182),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_146),
.B(n_182),
.Y(n_293)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_156),
.B1(n_173),
.B2(n_175),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_149),
.A2(n_174),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_156),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_156),
.A2(n_173),
.B1(n_343),
.B2(n_350),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_156),
.A2(n_173),
.B1(n_350),
.B2(n_361),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_156),
.A2(n_173),
.B1(n_361),
.B2(n_421),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_166),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_164),
.Y(n_157)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_158),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_164),
.Y(n_355)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_165),
.Y(n_353)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_165),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_172),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_173),
.B(n_225),
.Y(n_238)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_174),
.B(n_235),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_174),
.B(n_344),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_174),
.A2(n_223),
.B(n_235),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_175),
.Y(n_290)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_189),
.B(n_397),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_217),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_209),
.B2(n_216),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_201),
.B(n_216),
.C(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_204),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_217),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_235),
.B(n_238),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_223),
.A2(n_238),
.B(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_223),
.B(n_224),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_223),
.A2(n_440),
.B(n_441),
.Y(n_439)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_228),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.C(n_254),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_254),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.C(n_244),
.Y(n_233)
);

FAx1_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_239),
.CI(n_244),
.CON(n_257),
.SN(n_257)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_250),
.B(n_344),
.Y(n_412)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_277),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_256),
.B(n_277),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.C(n_259),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_257),
.B(n_448),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_257),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_258),
.B(n_259),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.C(n_269),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_260),
.A2(n_261),
.B1(n_267),
.B2(n_268),
.Y(n_435)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_263),
.B(n_344),
.Y(n_397)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_269),
.B(n_435),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g450 ( 
.A1(n_279),
.A2(n_307),
.B(n_451),
.C(n_454),
.D(n_455),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_306),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_280),
.B(n_306),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_284),
.C(n_305),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_292),
.B1(n_304),
.B2(n_305),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_289),
.B2(n_291),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_286),
.B1(n_326),
.B2(n_330),
.Y(n_325)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_286),
.B(n_289),
.Y(n_324)
);

AOI21xp33_ASAP7_75t_L g474 ( 
.A1(n_286),
.A2(n_324),
.B(n_326),
.Y(n_474)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_298),
.C(n_303),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_298),
.B1(n_299),
.B2(n_303),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_308),
.B(n_309),
.Y(n_455)
);

BUFx24_ASAP7_75t_SL g478 ( 
.A(n_309),
.Y(n_478)
);

FAx1_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.CI(n_323),
.CON(n_309),
.SN(n_309)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_310),
.B(n_311),
.C(n_323),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_319),
.B(n_322),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_319),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_SL g419 ( 
.A1(n_315),
.A2(n_344),
.B(n_412),
.Y(n_419)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_320),
.Y(n_441)
);

FAx1_ASAP7_75t_SL g460 ( 
.A(n_322),
.B(n_461),
.CI(n_474),
.CON(n_460),
.SN(n_460)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_328),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_445),
.B(n_449),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_430),
.B(n_444),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_401),
.B(n_429),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_373),
.B(n_400),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_356),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_336),
.B(n_356),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_342),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_342),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_349),
.Y(n_363)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_365),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_360),
.B2(n_364),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_358),
.B(n_364),
.C(n_365),
.Y(n_402)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_360),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_363),
.B(n_414),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_366),
.Y(n_380)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_384),
.B(n_399),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_383),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_375),
.B(n_383),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_394),
.B(n_398),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_386),
.B(n_387),
.Y(n_398)
);

INVx4_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_403),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_417),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_418),
.C(n_420),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_416),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_416),
.Y(n_438)
);

OAI32xp33_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_408),
.A3(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_421),
.Y(n_440)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_431),
.B(n_432),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_433),
.A2(n_434),
.B1(n_436),
.B2(n_437),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_439),
.C(n_442),
.Y(n_446)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_438),
.A2(n_439),
.B1(n_442),
.B2(n_443),
.Y(n_437)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_438),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_439),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_446),
.B(n_447),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_475),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_460),
.Y(n_476)
);

BUFx24_ASAP7_75t_SL g480 ( 
.A(n_460),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_469),
.B2(n_473),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_464),
.A2(n_465),
.B1(n_467),
.B2(n_468),
.Y(n_463)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_464),
.Y(n_468)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_465),
.Y(n_467)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_469),
.Y(n_473)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);


endmodule