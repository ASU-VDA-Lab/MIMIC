module fake_jpeg_31815_n_410 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_410);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_59),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_61),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_64),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_68),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_0),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_76),
.Y(n_109)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_75),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_1),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_46),
.Y(n_129)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_28),
.B1(n_35),
.B2(n_34),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_94),
.B1(n_31),
.B2(n_39),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_94),
.B(n_46),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_60),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_34),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_128),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_31),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_52),
.B(n_59),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_152),
.Y(n_179)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_30),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_30),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_153),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_97),
.A2(n_53),
.B1(n_47),
.B2(n_55),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_157),
.B1(n_158),
.B2(n_90),
.Y(n_167)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_78),
.B1(n_77),
.B2(n_65),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_164),
.B1(n_107),
.B2(n_90),
.Y(n_183)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx2_ASAP7_75t_R g152 ( 
.A(n_109),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_106),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_162),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_88),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_96),
.A2(n_29),
.B1(n_40),
.B2(n_39),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_100),
.A2(n_72),
.B1(n_71),
.B2(n_80),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_89),
.A2(n_84),
.B1(n_33),
.B2(n_45),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_32),
.CI(n_40),
.CON(n_182),
.SN(n_182)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_35),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_86),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_183),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_104),
.B1(n_88),
.B2(n_113),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_168),
.A2(n_146),
.B1(n_130),
.B2(n_107),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_SL g170 ( 
.A(n_152),
.B(n_99),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_105),
.B(n_38),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_172),
.B(n_182),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_135),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_104),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_190),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_154),
.C(n_139),
.Y(n_177)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_177),
.B(n_158),
.CI(n_164),
.CON(n_204),
.SN(n_204)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_139),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_151),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_156),
.Y(n_202)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_189),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_203),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_208),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_187),
.C(n_177),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

XNOR2x1_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_195),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_130),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_191),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_213),
.Y(n_240)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_183),
.B1(n_167),
.B2(n_168),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_185),
.A2(n_160),
.B1(n_148),
.B2(n_137),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_147),
.B1(n_194),
.B2(n_126),
.Y(n_243)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_38),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_216),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_178),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_187),
.A2(n_176),
.B(n_179),
.C(n_172),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_179),
.A3(n_182),
.B1(n_180),
.B2(n_169),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_224),
.A2(n_226),
.B1(n_231),
.B2(n_232),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_179),
.B1(n_188),
.B2(n_185),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_199),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_171),
.B1(n_182),
.B2(n_169),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_180),
.B1(n_134),
.B2(n_174),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_178),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_241),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_184),
.C(n_133),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_242),
.C(n_245),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_184),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_147),
.C(n_174),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_206),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_204),
.C(n_207),
.Y(n_245)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_263),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_218),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_247),
.B(n_251),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_240),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_249),
.Y(n_297)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_215),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_252),
.B(n_261),
.Y(n_300)
);

XOR2x2_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_204),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_269),
.B(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_224),
.A2(n_208),
.B1(n_202),
.B2(n_211),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_260),
.A2(n_234),
.B1(n_115),
.B2(n_102),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_230),
.B(n_216),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_232),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_198),
.C(n_197),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_225),
.A2(n_213),
.B1(n_214),
.B2(n_209),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_264),
.A2(n_272),
.B1(n_273),
.B2(n_236),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_32),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_226),
.B(n_200),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_268),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_241),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_213),
.C(n_133),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_163),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_199),
.B(n_135),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_262),
.B(n_274),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_210),
.B1(n_132),
.B2(n_161),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_222),
.A2(n_210),
.B1(n_144),
.B2(n_205),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_239),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_279),
.A2(n_280),
.B(n_285),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_282),
.B(n_258),
.Y(n_311)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_235),
.Y(n_284)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_228),
.B(n_221),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_286),
.A2(n_298),
.B(n_269),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_250),
.A2(n_221),
.B1(n_229),
.B2(n_236),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_289),
.A2(n_290),
.B1(n_155),
.B2(n_95),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_234),
.Y(n_291)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_259),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_296),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_299),
.B1(n_272),
.B2(n_273),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_125),
.C(n_155),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_249),
.B(n_1),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_148),
.B(n_163),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_258),
.A2(n_127),
.B1(n_111),
.B2(n_114),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_264),
.Y(n_303)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_263),
.C(n_270),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_307),
.C(n_310),
.Y(n_329)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_288),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_306),
.B(n_2),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_254),
.C(n_253),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_260),
.Y(n_309)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_309),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_254),
.C(n_256),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_321),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_312),
.A2(n_281),
.B(n_284),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_246),
.C(n_114),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_290),
.C(n_298),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_1),
.Y(n_315)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_316),
.A2(n_279),
.B1(n_294),
.B2(n_291),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_317),
.Y(n_335)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_277),
.Y(n_320)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_320),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_286),
.B(n_125),
.Y(n_321)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_322),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_287),
.B1(n_292),
.B2(n_299),
.Y(n_323)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_323),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_340),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_285),
.B(n_280),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_285),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_332),
.B(n_45),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_45),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_4),
.B(n_5),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_293),
.B1(n_283),
.B2(n_278),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_338),
.A2(n_314),
.B1(n_319),
.B2(n_308),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_278),
.Y(n_339)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_339),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_128),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_45),
.Y(n_355)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_5),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_307),
.C(n_304),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_345),
.C(n_348),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_313),
.C(n_318),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_350),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_321),
.C(n_322),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_339),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_357),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_2),
.C(n_4),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_352),
.B(n_6),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_4),
.Y(n_353)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_353),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_341),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_326),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_328),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_331),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_366),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_362),
.B(n_369),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_33),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_348),
.B(n_326),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_344),
.A2(n_327),
.B(n_335),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_370),
.A2(n_344),
.B(n_353),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_325),
.C(n_330),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_6),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_334),
.C(n_338),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_350),
.C(n_351),
.Y(n_375)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

XOR2x2_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_358),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_383),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_379),
.Y(n_384)
);

OAI211xp5_ASAP7_75t_SL g376 ( 
.A1(n_361),
.A2(n_356),
.B(n_346),
.C(n_324),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_376),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_336),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_381),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_8),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_365),
.Y(n_382)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_382),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_378),
.B(n_372),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_392),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_364),
.C(n_367),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_391),
.B(n_374),
.C(n_383),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_377),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_384),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_395),
.Y(n_402)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_386),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_396),
.B(n_399),
.Y(n_403)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_389),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_397),
.B(n_398),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_368),
.C(n_11),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_387),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_394),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_402),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_390),
.C(n_396),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_405),
.Y(n_406)
);

AOI322xp5_ASAP7_75t_L g407 ( 
.A1(n_406),
.A2(n_400),
.A3(n_391),
.B1(n_388),
.B2(n_14),
.C1(n_10),
.C2(n_12),
.Y(n_407)
);

O2A1O1Ixp33_ASAP7_75t_SL g408 ( 
.A1(n_407),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_408),
.Y(n_409)
);

AO21x1_ASAP7_75t_L g410 ( 
.A1(n_409),
.A2(n_11),
.B(n_16),
.Y(n_410)
);


endmodule