module fake_aes_5949_n_31 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_31);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVxp33_ASAP7_75t_SL g13 ( .A(n_1), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_10), .B(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_8), .Y(n_15) );
BUFx8_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
OAI21xp33_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_7), .B(n_11), .Y(n_18) );
OR2x2_ASAP7_75t_L g19 ( .A(n_17), .B(n_0), .Y(n_19) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_19), .Y(n_20) );
INVx2_ASAP7_75t_SL g21 ( .A(n_18), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_21), .B(n_15), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_21), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_14), .B(n_20), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
NOR2xp33_ASAP7_75t_L g26 ( .A(n_24), .B(n_16), .Y(n_26) );
NAND2xp33_ASAP7_75t_R g27 ( .A(n_26), .B(n_0), .Y(n_27) );
AND2x4_ASAP7_75t_L g28 ( .A(n_25), .B(n_1), .Y(n_28) );
AO21x1_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_16), .B(n_17), .Y(n_29) );
XNOR2xp5_ASAP7_75t_L g30 ( .A(n_29), .B(n_27), .Y(n_30) );
AO221x2_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_3), .B1(n_6), .B2(n_9), .C(n_12), .Y(n_31) );
endmodule