module fake_netlist_1_8070_n_951 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_951);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_951;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_838;
wire n_705;
wire n_949;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_383;
wire n_288;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_476;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_939;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_539;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_269;
NOR2xp67_ASAP7_75t_L g266 ( .A(n_41), .B(n_212), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_147), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_169), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_174), .Y(n_269) );
BUFx10_ASAP7_75t_L g270 ( .A(n_132), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_101), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_185), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_84), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_226), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_157), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_210), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_229), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_247), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_151), .Y(n_279) );
CKINVDCx14_ASAP7_75t_R g280 ( .A(n_261), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_227), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_84), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_48), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_253), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_252), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g286 ( .A(n_76), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_138), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_189), .Y(n_288) );
INVxp33_ASAP7_75t_SL g289 ( .A(n_141), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_208), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_188), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_88), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_113), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_73), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_116), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_5), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_57), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_191), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_206), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_86), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_140), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_152), .B(n_173), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_55), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_195), .Y(n_304) );
CKINVDCx16_ASAP7_75t_R g305 ( .A(n_137), .Y(n_305) );
INVxp33_ASAP7_75t_L g306 ( .A(n_43), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_263), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_109), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_211), .Y(n_309) );
INVxp67_ASAP7_75t_SL g310 ( .A(n_213), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_257), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_172), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_130), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_110), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_32), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_255), .Y(n_316) );
CKINVDCx14_ASAP7_75t_R g317 ( .A(n_96), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_190), .Y(n_318) );
INVxp33_ASAP7_75t_SL g319 ( .A(n_1), .Y(n_319) );
CKINVDCx14_ASAP7_75t_R g320 ( .A(n_178), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_161), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_214), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_120), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_68), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_89), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_46), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_217), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_43), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_223), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_79), .B(n_225), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_29), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_102), .Y(n_332) );
CKINVDCx16_ASAP7_75t_R g333 ( .A(n_216), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_184), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_237), .B(n_127), .Y(n_335) );
NOR2xp67_ASAP7_75t_L g336 ( .A(n_24), .B(n_207), .Y(n_336) );
NOR2xp67_ASAP7_75t_L g337 ( .A(n_67), .B(n_131), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_58), .Y(n_338) );
INVxp33_ASAP7_75t_L g339 ( .A(n_61), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_80), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_154), .Y(n_341) );
BUFx2_ASAP7_75t_SL g342 ( .A(n_146), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_103), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_75), .Y(n_344) );
BUFx10_ASAP7_75t_L g345 ( .A(n_11), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_91), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_149), .B(n_41), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_249), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_72), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_52), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_0), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_136), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_42), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_44), .Y(n_354) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_193), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_199), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_181), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_187), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_200), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_95), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_88), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_244), .Y(n_362) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_175), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_20), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_209), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_33), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_17), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_32), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_155), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_127), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_6), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_239), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_144), .Y(n_373) );
NOR2xp67_ASAP7_75t_L g374 ( .A(n_145), .B(n_150), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_107), .Y(n_375) );
INVxp33_ASAP7_75t_L g376 ( .A(n_61), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_201), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_129), .B(n_158), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_115), .Y(n_379) );
INVxp33_ASAP7_75t_SL g380 ( .A(n_108), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_243), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_13), .Y(n_382) );
INVxp67_ASAP7_75t_L g383 ( .A(n_221), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_204), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_83), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_5), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_171), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_79), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_100), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_220), .Y(n_390) );
BUFx5_ASAP7_75t_L g391 ( .A(n_166), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_251), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_265), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_228), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_242), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_148), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_236), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_11), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_51), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_163), .B(n_230), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_231), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_53), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_215), .Y(n_403) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_180), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_260), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_69), .Y(n_406) );
INVxp33_ASAP7_75t_L g407 ( .A(n_49), .Y(n_407) );
BUFx3_ASAP7_75t_L g408 ( .A(n_97), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_16), .Y(n_409) );
INVxp33_ASAP7_75t_SL g410 ( .A(n_50), .Y(n_410) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_183), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_258), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_331), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_341), .B(n_0), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_331), .B(n_2), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_331), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_385), .B(n_2), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_385), .B(n_3), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_317), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_341), .B(n_329), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_315), .B(n_3), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_341), .B(n_408), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_317), .A2(n_7), .B1(n_4), .B2(n_6), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_408), .B(n_4), .Y(n_425) );
CKINVDCx8_ASAP7_75t_R g426 ( .A(n_305), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_282), .Y(n_428) );
INVx6_ASAP7_75t_L g429 ( .A(n_270), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_298), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_350), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_306), .B(n_8), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_338), .B(n_9), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_348), .B(n_10), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_282), .B(n_10), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_306), .B(n_12), .Y(n_437) );
INVx5_ASAP7_75t_L g438 ( .A(n_298), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_339), .B(n_12), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_295), .Y(n_440) );
OR2x6_ASAP7_75t_L g441 ( .A(n_342), .B(n_14), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_295), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_298), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_283), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_297), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_339), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_298), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_268), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_301), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_297), .B(n_15), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_301), .Y(n_451) );
AND2x2_ASAP7_75t_SL g452 ( .A(n_333), .B(n_128), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_430), .Y(n_453) );
BUFx10_ASAP7_75t_L g454 ( .A(n_429), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_446), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_427), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_427), .Y(n_457) );
NAND2xp33_ASAP7_75t_L g458 ( .A(n_419), .B(n_391), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_435), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_423), .B(n_413), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_435), .Y(n_461) );
INVx5_ASAP7_75t_L g462 ( .A(n_413), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_415), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_415), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_415), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_430), .Y(n_466) );
BUFx6f_ASAP7_75t_SL g467 ( .A(n_452), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_417), .Y(n_468) );
INVx6_ASAP7_75t_L g469 ( .A(n_423), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_430), .Y(n_470) );
OR2x6_ASAP7_75t_L g471 ( .A(n_441), .B(n_340), .Y(n_471) );
NAND2xp33_ASAP7_75t_L g472 ( .A(n_419), .B(n_391), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_429), .B(n_376), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_417), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_429), .B(n_291), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_429), .B(n_407), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_420), .B(n_304), .Y(n_477) );
INVx6_ASAP7_75t_L g478 ( .A(n_423), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_444), .B(n_407), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_413), .B(n_283), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_432), .B(n_280), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_431), .A2(n_380), .B1(n_410), .B2(n_319), .Y(n_482) );
INVx4_ASAP7_75t_SL g483 ( .A(n_418), .Y(n_483) );
OR2x6_ASAP7_75t_L g484 ( .A(n_441), .B(n_340), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_426), .B(n_383), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_418), .B(n_354), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_432), .B(n_280), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_418), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_430), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_437), .B(n_286), .Y(n_490) );
BUFx4f_ASAP7_75t_L g491 ( .A(n_425), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_479), .A2(n_455), .B(n_439), .C(n_490), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_464), .A2(n_436), .B1(n_450), .B2(n_441), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_490), .A2(n_433), .B(n_421), .C(n_424), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_491), .B(n_452), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_481), .B(n_434), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_481), .B(n_425), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_487), .B(n_425), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_477), .B(n_426), .Y(n_499) );
INVx3_ASAP7_75t_SL g500 ( .A(n_471), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_469), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_491), .B(n_436), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_487), .B(n_448), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_483), .B(n_436), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_464), .A2(n_450), .B1(n_448), .B2(n_422), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_459), .Y(n_506) );
NAND2x1_ASAP7_75t_L g507 ( .A(n_471), .B(n_450), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_473), .B(n_289), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_476), .B(n_345), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_460), .B(n_416), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_483), .B(n_267), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_465), .A2(n_422), .B1(n_410), .B2(n_319), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_467), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_480), .B(n_281), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_483), .B(n_272), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_482), .B(n_292), .Y(n_516) );
OR2x6_ASAP7_75t_L g517 ( .A(n_484), .B(n_414), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_478), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_459), .Y(n_519) );
INVx8_ASAP7_75t_L g520 ( .A(n_484), .Y(n_520) );
NOR2xp67_ASAP7_75t_L g521 ( .A(n_485), .B(n_440), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_468), .A2(n_299), .B1(n_311), .B2(n_285), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_456), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_462), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_467), .A2(n_334), .B1(n_393), .B2(n_313), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_475), .B(n_281), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_478), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_486), .B(n_287), .Y(n_528) );
INVx4_ASAP7_75t_L g529 ( .A(n_454), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_486), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_474), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_474), .A2(n_393), .B1(n_334), .B2(n_371), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_463), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_488), .B(n_287), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_488), .A2(n_371), .B1(n_375), .B2(n_367), .Y(n_535) );
NAND2x1p5_ASAP7_75t_L g536 ( .A(n_463), .B(n_294), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_463), .B(n_428), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_457), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_458), .B(n_289), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_457), .A2(n_445), .B1(n_442), .B2(n_296), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_462), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_461), .B(n_373), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_466), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_466), .B(n_276), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_453), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_470), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_472), .B(n_320), .Y(n_547) );
INVx4_ASAP7_75t_L g548 ( .A(n_453), .Y(n_548) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_511), .A2(n_400), .B(n_330), .C(n_278), .Y(n_549) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_520), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_495), .A2(n_343), .B1(n_382), .B2(n_293), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_504), .A2(n_312), .B(n_310), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_529), .B(n_274), .Y(n_553) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_520), .Y(n_554) );
NOR2xp33_ASAP7_75t_R g555 ( .A(n_513), .B(n_293), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_504), .A2(n_404), .B(n_355), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_497), .A2(n_411), .B(n_279), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_523), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_492), .A2(n_303), .B(n_314), .C(n_308), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_498), .A2(n_284), .B(n_277), .Y(n_560) );
INVx4_ASAP7_75t_L g561 ( .A(n_500), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_502), .A2(n_290), .B(n_288), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_537), .Y(n_563) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_500), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_523), .Y(n_565) );
NOR2xp33_ASAP7_75t_SL g566 ( .A(n_522), .B(n_343), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_493), .A2(n_382), .B1(n_375), .B2(n_379), .Y(n_567) );
AOI21x1_ASAP7_75t_L g568 ( .A1(n_511), .A2(n_489), .B(n_470), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_508), .B(n_271), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_499), .B(n_273), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_530), .A2(n_323), .B(n_325), .C(n_324), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_508), .B(n_300), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_547), .A2(n_321), .B(n_309), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_538), .Y(n_574) );
O2A1O1Ixp5_ASAP7_75t_L g575 ( .A1(n_507), .A2(n_335), .B(n_269), .C(n_316), .Y(n_575) );
O2A1O1Ixp33_ASAP7_75t_L g576 ( .A1(n_495), .A2(n_328), .B(n_332), .C(n_326), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_501), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_533), .A2(n_357), .B(n_356), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_534), .A2(n_365), .B(n_359), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_536), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_503), .B(n_344), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_516), .B(n_349), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_509), .B(n_351), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_535), .B(n_389), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g585 ( .A1(n_510), .A2(n_353), .B(n_366), .C(n_360), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_539), .A2(n_370), .B(n_386), .C(n_368), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_521), .B(n_307), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_514), .A2(n_384), .B(n_381), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_512), .B(n_388), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_505), .A2(n_347), .B1(n_402), .B2(n_398), .Y(n_590) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_506), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_542), .A2(n_394), .B(n_392), .Y(n_592) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_506), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g594 ( .A1(n_528), .A2(n_409), .B(n_361), .C(n_364), .Y(n_594) );
INVx4_ASAP7_75t_L g595 ( .A(n_501), .Y(n_595) );
INVx2_ASAP7_75t_SL g596 ( .A(n_517), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g597 ( .A1(n_519), .A2(n_336), .B(n_337), .C(n_266), .Y(n_597) );
BUFx2_ASAP7_75t_L g598 ( .A(n_532), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_526), .B(n_354), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_525), .A2(n_361), .B1(n_399), .B2(n_364), .Y(n_600) );
AO21x1_ASAP7_75t_L g601 ( .A1(n_544), .A2(n_397), .B(n_396), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_540), .A2(n_406), .B(n_399), .C(n_405), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_540), .B(n_406), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_519), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_515), .A2(n_412), .B(n_401), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_518), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_515), .A2(n_316), .B(n_275), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_544), .A2(n_318), .B(n_275), .Y(n_608) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_527), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_543), .A2(n_322), .B(n_318), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_541), .A2(n_322), .B(n_369), .C(n_327), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_L g612 ( .A1(n_524), .A2(n_377), .B(n_395), .C(n_387), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_548), .B(n_372), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_548), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_546), .A2(n_377), .B(n_395), .C(n_387), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_546), .Y(n_616) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_545), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_L g618 ( .A1(n_494), .A2(n_302), .B(n_378), .C(n_374), .Y(n_618) );
BUFx2_ASAP7_75t_L g619 ( .A(n_500), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_493), .A2(n_346), .B1(n_358), .B2(n_352), .Y(n_620) );
OR2x6_ASAP7_75t_L g621 ( .A(n_520), .B(n_346), .Y(n_621) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_531), .A2(n_346), .B(n_362), .C(n_301), .Y(n_622) );
OR2x6_ASAP7_75t_L g623 ( .A(n_520), .B(n_346), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_496), .B(n_390), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_537), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_499), .B(n_403), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_504), .A2(n_453), .B(n_438), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_563), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_573), .A2(n_616), .B(n_604), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_558), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_564), .B(n_391), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_575), .A2(n_438), .B(n_391), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_565), .Y(n_633) );
INVx5_ASAP7_75t_L g634 ( .A(n_621), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_621), .A2(n_363), .B1(n_438), .B2(n_443), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_574), .A2(n_453), .B(n_363), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_623), .A2(n_447), .B1(n_449), .B2(n_443), .Y(n_637) );
NOR2x1_ASAP7_75t_SL g638 ( .A(n_623), .B(n_443), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_567), .B(n_551), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_562), .A2(n_451), .B(n_449), .Y(n_640) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_617), .Y(n_641) );
O2A1O1Ixp5_ASAP7_75t_L g642 ( .A1(n_601), .A2(n_451), .B(n_133), .C(n_134), .Y(n_642) );
AO32x2_ASAP7_75t_L g643 ( .A1(n_590), .A2(n_451), .A3(n_21), .B1(n_18), .B2(n_19), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_625), .Y(n_644) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_568), .A2(n_139), .B(n_135), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_582), .B(n_22), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_564), .Y(n_647) );
OAI21x1_ASAP7_75t_L g648 ( .A1(n_627), .A2(n_143), .B(n_142), .Y(n_648) );
AO31x2_ASAP7_75t_L g649 ( .A1(n_597), .A2(n_26), .A3(n_23), .B(n_25), .Y(n_649) );
AO31x2_ASAP7_75t_L g650 ( .A1(n_610), .A2(n_28), .A3(n_25), .B(n_27), .Y(n_650) );
INVx5_ASAP7_75t_L g651 ( .A(n_550), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_596), .B(n_28), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_570), .B(n_30), .Y(n_653) );
AO32x2_ASAP7_75t_L g654 ( .A1(n_600), .A2(n_30), .A3(n_31), .B1(n_33), .B2(n_34), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_619), .B(n_31), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_580), .A2(n_37), .B1(n_35), .B2(n_36), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_571), .A2(n_589), .B1(n_584), .B2(n_586), .C(n_585), .Y(n_657) );
INVx8_ASAP7_75t_L g658 ( .A(n_554), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_576), .A2(n_40), .B(n_38), .C(n_39), .Y(n_659) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_554), .Y(n_660) );
BUFx4f_ASAP7_75t_L g661 ( .A(n_554), .Y(n_661) );
INVx3_ASAP7_75t_L g662 ( .A(n_561), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_560), .A2(n_557), .B(n_588), .Y(n_663) );
BUFx3_ASAP7_75t_L g664 ( .A(n_609), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_583), .B(n_39), .Y(n_665) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_591), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_594), .A2(n_611), .B(n_579), .C(n_592), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_591), .Y(n_668) );
AO31x2_ASAP7_75t_L g669 ( .A1(n_607), .A2(n_47), .A3(n_45), .B(n_46), .Y(n_669) );
AO21x1_ASAP7_75t_L g670 ( .A1(n_615), .A2(n_156), .B(n_153), .Y(n_670) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_591), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_599), .A2(n_160), .B(n_159), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_624), .A2(n_164), .B(n_162), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_549), .A2(n_167), .B(n_165), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_569), .A2(n_170), .B(n_168), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_626), .A2(n_603), .B1(n_581), .B2(n_572), .Y(n_676) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_593), .Y(n_677) );
AO31x2_ASAP7_75t_L g678 ( .A1(n_608), .A2(n_54), .A3(n_56), .B(n_59), .Y(n_678) );
O2A1O1Ixp5_ASAP7_75t_L g679 ( .A1(n_587), .A2(n_177), .B(n_264), .C(n_262), .Y(n_679) );
AO32x2_ASAP7_75t_L g680 ( .A1(n_620), .A2(n_60), .A3(n_62), .B1(n_63), .B2(n_64), .Y(n_680) );
AO31x2_ASAP7_75t_L g681 ( .A1(n_606), .A2(n_64), .A3(n_65), .B(n_66), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_578), .A2(n_179), .B(n_176), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_552), .B(n_68), .Y(n_683) );
AO31x2_ASAP7_75t_L g684 ( .A1(n_605), .A2(n_70), .A3(n_71), .B(n_72), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_614), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_556), .B(n_74), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_602), .Y(n_687) );
AO31x2_ASAP7_75t_L g688 ( .A1(n_613), .A2(n_74), .A3(n_75), .B(n_77), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_577), .B(n_77), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_609), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_577), .Y(n_691) );
AO32x2_ASAP7_75t_L g692 ( .A1(n_595), .A2(n_78), .A3(n_80), .B1(n_81), .B2(n_82), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_553), .Y(n_693) );
AO31x2_ASAP7_75t_L g694 ( .A1(n_612), .A2(n_85), .A3(n_86), .B(n_87), .Y(n_694) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_559), .A2(n_87), .B(n_89), .C(n_90), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_573), .A2(n_196), .B(n_259), .Y(n_696) );
AO21x1_ASAP7_75t_L g697 ( .A1(n_618), .A2(n_197), .B(n_256), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_555), .Y(n_698) );
AO31x2_ASAP7_75t_L g699 ( .A1(n_612), .A2(n_92), .A3(n_93), .B(n_94), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_573), .A2(n_198), .B(n_254), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_573), .A2(n_194), .B(n_250), .Y(n_701) );
AO32x2_ASAP7_75t_L g702 ( .A1(n_590), .A2(n_98), .A3(n_99), .B1(n_100), .B2(n_101), .Y(n_702) );
AO21x1_ASAP7_75t_L g703 ( .A1(n_618), .A2(n_205), .B(n_248), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_566), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_676), .A2(n_218), .B(n_246), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g706 ( .A1(n_687), .A2(n_111), .B(n_112), .Y(n_706) );
AO31x2_ASAP7_75t_L g707 ( .A1(n_670), .A2(n_114), .A3(n_115), .B(n_116), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_639), .B(n_117), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_630), .Y(n_709) );
AO21x2_ASAP7_75t_L g710 ( .A1(n_632), .A2(n_224), .B(n_245), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_667), .A2(n_222), .B(n_241), .Y(n_711) );
AO21x2_ASAP7_75t_L g712 ( .A1(n_697), .A2(n_219), .B(n_240), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_642), .A2(n_118), .B(n_119), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_636), .A2(n_640), .B(n_674), .Y(n_714) );
AO31x2_ASAP7_75t_L g715 ( .A1(n_703), .A2(n_121), .A3(n_122), .B(n_123), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_633), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_628), .B(n_121), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_658), .Y(n_718) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_634), .Y(n_719) );
AO31x2_ASAP7_75t_L g720 ( .A1(n_659), .A2(n_124), .A3(n_125), .B(n_126), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g721 ( .A1(n_683), .A2(n_182), .B(n_186), .Y(n_721) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_641), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_644), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_655), .B(n_192), .Y(n_724) );
BUFx6f_ASAP7_75t_L g725 ( .A(n_641), .Y(n_725) );
OAI21x1_ASAP7_75t_L g726 ( .A1(n_648), .A2(n_202), .B(n_203), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_702), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_685), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_702), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_665), .B(n_232), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_698), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_652), .A2(n_233), .B1(n_234), .B2(n_235), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_702), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_693), .B(n_238), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_643), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_686), .B(n_695), .Y(n_736) );
OR2x2_ASAP7_75t_L g737 ( .A(n_662), .B(n_647), .Y(n_737) );
AND2x4_ASAP7_75t_L g738 ( .A(n_660), .B(n_664), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_673), .A2(n_675), .B(n_672), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_666), .B(n_671), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_679), .A2(n_700), .B(n_696), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_643), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_643), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_681), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_701), .A2(n_689), .B(n_682), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_691), .B(n_668), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_704), .B(n_656), .Y(n_747) );
BUFx3_ASAP7_75t_L g748 ( .A(n_690), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_681), .Y(n_749) );
NOR2xp67_ASAP7_75t_L g750 ( .A(n_635), .B(n_631), .Y(n_750) );
AND2x4_ASAP7_75t_L g751 ( .A(n_638), .B(n_671), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_684), .Y(n_752) );
INVx2_ASAP7_75t_SL g753 ( .A(n_666), .Y(n_753) );
AND2x4_ASAP7_75t_L g754 ( .A(n_666), .B(n_677), .Y(n_754) );
BUFx2_ASAP7_75t_L g755 ( .A(n_677), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_637), .A2(n_699), .B(n_694), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_684), .Y(n_757) );
BUFx8_ASAP7_75t_L g758 ( .A(n_692), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_654), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_654), .A2(n_680), .B1(n_692), .B2(n_649), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_654), .A2(n_680), .B1(n_692), .B2(n_649), .Y(n_761) );
INVx2_ASAP7_75t_SL g762 ( .A(n_694), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_669), .A2(n_678), .B(n_650), .Y(n_763) );
NOR2xp67_ASAP7_75t_L g764 ( .A(n_688), .B(n_678), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_688), .B(n_598), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_657), .B(n_687), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_L g767 ( .A1(n_653), .A2(n_646), .B(n_663), .C(n_667), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_657), .B(n_687), .Y(n_768) );
OAI21xp5_ASAP7_75t_L g769 ( .A1(n_687), .A2(n_676), .B(n_629), .Y(n_769) );
INVx3_ASAP7_75t_L g770 ( .A(n_651), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_661), .Y(n_771) );
AO31x2_ASAP7_75t_L g772 ( .A1(n_670), .A2(n_697), .A3(n_703), .B(n_622), .Y(n_772) );
OA21x2_ASAP7_75t_L g773 ( .A1(n_632), .A2(n_642), .B(n_645), .Y(n_773) );
AO31x2_ASAP7_75t_L g774 ( .A1(n_670), .A2(n_697), .A3(n_703), .B(n_622), .Y(n_774) );
AND2x4_ASAP7_75t_L g775 ( .A(n_651), .B(n_550), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_657), .B(n_687), .Y(n_776) );
INVx2_ASAP7_75t_SL g777 ( .A(n_661), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_657), .B(n_687), .Y(n_778) );
OA21x2_ASAP7_75t_L g779 ( .A1(n_632), .A2(n_642), .B(n_645), .Y(n_779) );
NAND2x1p5_ASAP7_75t_L g780 ( .A(n_651), .B(n_634), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_765), .B(n_708), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_709), .B(n_716), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_751), .B(n_754), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_766), .B(n_768), .Y(n_784) );
AO21x2_ASAP7_75t_L g785 ( .A1(n_764), .A2(n_756), .B(n_769), .Y(n_785) );
BUFx2_ASAP7_75t_L g786 ( .A(n_758), .Y(n_786) );
AND2x4_ASAP7_75t_L g787 ( .A(n_722), .B(n_725), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_723), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_744), .Y(n_789) );
OA21x2_ASAP7_75t_L g790 ( .A1(n_752), .A2(n_757), .B(n_749), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_722), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_725), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_725), .Y(n_793) );
OA21x2_ASAP7_75t_L g794 ( .A1(n_760), .A2(n_761), .B(n_742), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_717), .Y(n_795) );
INVx4_ASAP7_75t_L g796 ( .A(n_780), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_766), .B(n_768), .Y(n_797) );
OA21x2_ASAP7_75t_L g798 ( .A1(n_735), .A2(n_743), .B(n_767), .Y(n_798) );
AND2x4_ASAP7_75t_L g799 ( .A(n_753), .B(n_775), .Y(n_799) );
OA21x2_ASAP7_75t_L g800 ( .A1(n_727), .A2(n_733), .B(n_729), .Y(n_800) );
AO21x2_ASAP7_75t_L g801 ( .A1(n_713), .A2(n_745), .B(n_714), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_776), .B(n_778), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_759), .B(n_746), .Y(n_803) );
INVx3_ASAP7_75t_L g804 ( .A(n_775), .Y(n_804) );
BUFx2_ASAP7_75t_L g805 ( .A(n_758), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_728), .B(n_706), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_720), .B(n_724), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_747), .B(n_762), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_720), .B(n_736), .Y(n_809) );
BUFx4f_ASAP7_75t_SL g810 ( .A(n_731), .Y(n_810) );
AND2x4_ASAP7_75t_L g811 ( .A(n_770), .B(n_755), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_737), .Y(n_812) );
AND2x4_ASAP7_75t_L g813 ( .A(n_738), .B(n_748), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_720), .B(n_736), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_719), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_739), .A2(n_741), .B(n_711), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_738), .B(n_715), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_771), .B(n_718), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_730), .B(n_734), .Y(n_819) );
OR2x6_ASAP7_75t_L g820 ( .A(n_740), .B(n_721), .Y(n_820) );
BUFx3_ASAP7_75t_L g821 ( .A(n_777), .Y(n_821) );
BUFx2_ASAP7_75t_L g822 ( .A(n_710), .Y(n_822) );
OR2x6_ASAP7_75t_L g823 ( .A(n_730), .B(n_705), .Y(n_823) );
AND2x4_ASAP7_75t_L g824 ( .A(n_710), .B(n_726), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_707), .B(n_732), .Y(n_825) );
AND2x4_ASAP7_75t_L g826 ( .A(n_750), .B(n_712), .Y(n_826) );
AND2x4_ASAP7_75t_L g827 ( .A(n_772), .B(n_774), .Y(n_827) );
OR2x6_ASAP7_75t_L g828 ( .A(n_773), .B(n_779), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_774), .B(n_779), .Y(n_829) );
AO21x2_ASAP7_75t_L g830 ( .A1(n_763), .A2(n_764), .B(n_756), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_709), .B(n_716), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_789), .Y(n_832) );
AND2x4_ASAP7_75t_L g833 ( .A(n_786), .B(n_805), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_789), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_809), .B(n_814), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_800), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_800), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_781), .B(n_808), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_809), .B(n_814), .Y(n_839) );
INVx5_ASAP7_75t_L g840 ( .A(n_796), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_794), .B(n_797), .Y(n_841) );
AO21x2_ASAP7_75t_L g842 ( .A1(n_816), .A2(n_829), .B(n_825), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_790), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_790), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_790), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_784), .B(n_802), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_794), .B(n_817), .Y(n_847) );
INVx2_ASAP7_75t_SL g848 ( .A(n_813), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_798), .B(n_807), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_803), .B(n_784), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_798), .B(n_807), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_798), .B(n_782), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_782), .B(n_831), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_810), .B(n_818), .Y(n_854) );
AND2x2_ASAP7_75t_SL g855 ( .A(n_824), .B(n_826), .Y(n_855) );
INVx3_ASAP7_75t_L g856 ( .A(n_787), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_788), .Y(n_857) );
INVx3_ASAP7_75t_L g858 ( .A(n_820), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_812), .B(n_795), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_827), .B(n_806), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_835), .B(n_827), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_832), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_853), .B(n_815), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_835), .B(n_785), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_854), .B(n_821), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_834), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_839), .B(n_860), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_839), .B(n_785), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_860), .B(n_785), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_847), .B(n_830), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_847), .B(n_830), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_841), .B(n_830), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_841), .B(n_801), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_849), .B(n_801), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_846), .B(n_811), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_849), .B(n_822), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_851), .B(n_822), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_852), .B(n_828), .Y(n_878) );
OR2x2_ASAP7_75t_L g879 ( .A(n_838), .B(n_828), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_852), .B(n_828), .Y(n_880) );
INVx4_ASAP7_75t_L g881 ( .A(n_840), .Y(n_881) );
OR2x2_ASAP7_75t_L g882 ( .A(n_850), .B(n_819), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_859), .B(n_783), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_843), .Y(n_884) );
BUFx3_ASAP7_75t_L g885 ( .A(n_840), .Y(n_885) );
OR2x2_ASAP7_75t_L g886 ( .A(n_867), .B(n_833), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_867), .B(n_855), .Y(n_887) );
AND2x2_ASAP7_75t_L g888 ( .A(n_864), .B(n_855), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_864), .B(n_858), .Y(n_889) );
NAND2x1_ASAP7_75t_L g890 ( .A(n_881), .B(n_833), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_868), .B(n_858), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_884), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_868), .B(n_858), .Y(n_893) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_865), .B(n_833), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_870), .B(n_836), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_870), .B(n_837), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_862), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_882), .B(n_857), .Y(n_898) );
INVx3_ASAP7_75t_L g899 ( .A(n_881), .Y(n_899) );
OR2x2_ASAP7_75t_L g900 ( .A(n_873), .B(n_879), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_873), .B(n_842), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_871), .B(n_842), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_866), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_871), .B(n_842), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_872), .B(n_844), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_872), .B(n_844), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_874), .B(n_845), .Y(n_907) );
INVx1_ASAP7_75t_SL g908 ( .A(n_885), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_898), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_907), .B(n_874), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_902), .B(n_869), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_902), .B(n_869), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_907), .B(n_863), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_895), .B(n_861), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_897), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_904), .B(n_878), .Y(n_916) );
NOR2x1_ASAP7_75t_L g917 ( .A(n_890), .B(n_885), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_896), .B(n_876), .Y(n_918) );
OR2x2_ASAP7_75t_L g919 ( .A(n_901), .B(n_876), .Y(n_919) );
OR2x2_ASAP7_75t_L g920 ( .A(n_901), .B(n_877), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_904), .B(n_878), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_903), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_896), .B(n_880), .Y(n_923) );
INVx3_ASAP7_75t_L g924 ( .A(n_899), .Y(n_924) );
INVx1_ASAP7_75t_SL g925 ( .A(n_886), .Y(n_925) );
OR2x2_ASAP7_75t_L g926 ( .A(n_900), .B(n_877), .Y(n_926) );
INVx1_ASAP7_75t_SL g927 ( .A(n_925), .Y(n_927) );
OR2x2_ASAP7_75t_L g928 ( .A(n_919), .B(n_900), .Y(n_928) );
AOI32xp33_ASAP7_75t_L g929 ( .A1(n_917), .A2(n_887), .A3(n_888), .B1(n_894), .B2(n_908), .Y(n_929) );
OR2x2_ASAP7_75t_L g930 ( .A(n_919), .B(n_905), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_911), .B(n_905), .Y(n_931) );
OR2x2_ASAP7_75t_L g932 ( .A(n_920), .B(n_906), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_915), .Y(n_933) );
AOI322xp5_ASAP7_75t_L g934 ( .A1(n_911), .A2(n_912), .A3(n_910), .B1(n_918), .B2(n_916), .C1(n_921), .C2(n_913), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_929), .A2(n_924), .B1(n_926), .B2(n_914), .Y(n_935) );
HB1xp67_ASAP7_75t_L g936 ( .A(n_927), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_928), .Y(n_937) );
OAI211xp5_ASAP7_75t_SL g938 ( .A1(n_934), .A2(n_909), .B(n_875), .C(n_922), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_936), .B(n_923), .Y(n_939) );
AOI221xp5_ASAP7_75t_L g940 ( .A1(n_938), .A2(n_933), .B1(n_931), .B2(n_932), .C(n_930), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g941 ( .A1(n_935), .A2(n_889), .B1(n_891), .B2(n_893), .C(n_883), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_937), .Y(n_942) );
NAND4xp25_ASAP7_75t_SL g943 ( .A(n_941), .B(n_940), .C(n_939), .D(n_942), .Y(n_943) );
NOR3xp33_ASAP7_75t_L g944 ( .A(n_943), .B(n_804), .C(n_848), .Y(n_944) );
NOR3xp33_ASAP7_75t_L g945 ( .A(n_944), .B(n_799), .C(n_856), .Y(n_945) );
INVx4_ASAP7_75t_L g946 ( .A(n_945), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_946), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_947), .A2(n_799), .B(n_823), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_948), .B(n_892), .Y(n_949) );
OR2x6_ASAP7_75t_L g950 ( .A(n_949), .B(n_791), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g951 ( .A1(n_950), .A2(n_792), .B(n_793), .Y(n_951) );
endmodule