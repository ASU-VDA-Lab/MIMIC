module fake_jpeg_1532_n_590 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_590);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_590;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_4),
.B(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_12),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_16),
.B(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

AND2x4_ASAP7_75t_SL g60 ( 
.A(n_33),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_60),
.B(n_75),
.Y(n_129)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_63),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_67),
.B(n_83),
.Y(n_162)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_70),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_51),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_72),
.B(n_104),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_74),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g201 ( 
.A(n_77),
.Y(n_201)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_84),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_85),
.Y(n_203)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_92),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_88),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_90),
.Y(n_213)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_93),
.Y(n_163)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_32),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_98),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_97),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_23),
.B(n_17),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_107),
.Y(n_143)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g198 ( 
.A(n_103),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_51),
.B(n_17),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_28),
.B(n_16),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_23),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_117),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_29),
.B(n_14),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_113),
.B(n_37),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_123),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_45),
.B(n_15),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_43),
.Y(n_137)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_29),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_27),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_31),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_31),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_137),
.B(n_176),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_75),
.B(n_50),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_139),
.B(n_153),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_50),
.B1(n_43),
.B2(n_68),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_147),
.B(n_42),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_148),
.B(n_158),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_30),
.Y(n_153)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_64),
.A2(n_30),
.B1(n_27),
.B2(n_24),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_166),
.A2(n_174),
.B1(n_36),
.B2(n_53),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_169),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_60),
.B(n_24),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_170),
.A2(n_175),
.B(n_181),
.C(n_193),
.Y(n_266)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_171),
.B(n_7),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_65),
.A2(n_26),
.B1(n_37),
.B2(n_15),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_1),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_59),
.B(n_1),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_66),
.Y(n_178)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_69),
.Y(n_179)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_119),
.B(n_63),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_103),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_199),
.Y(n_214)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_185),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_85),
.B(n_1),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_105),
.B(n_2),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_195),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_93),
.B(n_3),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_106),
.B(n_3),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_202),
.Y(n_248)
);

BUFx16f_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

CKINVDCx6p67_ASAP7_75t_R g249 ( 
.A(n_200),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_109),
.B(n_86),
.Y(n_202)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_110),
.B(n_26),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_77),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_112),
.B(n_5),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_210),
.B(n_7),
.Y(n_261)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_215),
.Y(n_292)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_216),
.Y(n_302)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_218),
.Y(n_300)
);

OA22x2_ASAP7_75t_L g219 ( 
.A1(n_170),
.A2(n_89),
.B1(n_116),
.B2(n_115),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_219),
.B(n_226),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_129),
.A2(n_102),
.B1(n_26),
.B2(n_77),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_220),
.A2(n_269),
.B1(n_273),
.B2(n_287),
.Y(n_289)
);

CKINVDCx9p33_ASAP7_75t_R g221 ( 
.A(n_191),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_221),
.Y(n_297)
);

CKINVDCx12_ASAP7_75t_R g222 ( 
.A(n_209),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_222),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_223),
.Y(n_321)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_225),
.Y(n_343)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_227),
.Y(n_326)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_136),
.Y(n_228)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_228),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_128),
.Y(n_235)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_235),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_151),
.B(n_5),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_236),
.B(n_241),
.Y(n_291)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_171),
.A2(n_19),
.B1(n_53),
.B2(n_36),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_239),
.A2(n_256),
.B1(n_282),
.B2(n_283),
.Y(n_290)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_130),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_240),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_151),
.B(n_5),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_150),
.Y(n_244)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_244),
.Y(n_306)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_245),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_129),
.B(n_6),
.C(n_7),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_246),
.B(n_255),
.Y(n_305)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_163),
.Y(n_250)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_252),
.Y(n_296)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_133),
.Y(n_253)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_152),
.B(n_7),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_181),
.A2(n_36),
.B1(n_53),
.B2(n_19),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_257),
.A2(n_258),
.B1(n_277),
.B2(n_239),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_196),
.A2(n_42),
.B1(n_48),
.B2(n_91),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_164),
.Y(n_259)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_261),
.B(n_262),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_143),
.B(n_10),
.Y(n_262)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_140),
.Y(n_263)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_155),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_265),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_191),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_271),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_140),
.Y(n_268)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_268),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_193),
.A2(n_42),
.B1(n_48),
.B2(n_13),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_270),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_143),
.B(n_10),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_210),
.A2(n_42),
.B1(n_48),
.B2(n_12),
.Y(n_273)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_211),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_274),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_142),
.B(n_12),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_278),
.Y(n_325)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_142),
.A2(n_13),
.B1(n_48),
.B2(n_197),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_138),
.B(n_13),
.C(n_152),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_126),
.Y(n_279)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_192),
.Y(n_280)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_186),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_281),
.Y(n_331)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_145),
.Y(n_283)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_149),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_189),
.Y(n_295)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_161),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_286),
.A2(n_126),
.B1(n_203),
.B2(n_212),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_195),
.A2(n_175),
.B1(n_167),
.B2(n_213),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

AND2x2_ASAP7_75t_SL g299 ( 
.A(n_248),
.B(n_135),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_299),
.B(n_312),
.Y(n_367)
);

OAI22x1_ASAP7_75t_L g310 ( 
.A1(n_214),
.A2(n_202),
.B1(n_169),
.B2(n_138),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_310),
.A2(n_318),
.B1(n_249),
.B2(n_228),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_256),
.A2(n_196),
.B(n_203),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_313),
.A2(n_230),
.B(n_245),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_198),
.B1(n_146),
.B2(n_189),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_316),
.A2(n_335),
.B1(n_258),
.B2(n_263),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_237),
.B(n_266),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_332),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_259),
.A2(n_212),
.B1(n_144),
.B2(n_141),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_269),
.A2(n_198),
.B1(n_159),
.B2(n_162),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_320),
.B(n_327),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_233),
.A2(n_167),
.B1(n_204),
.B2(n_213),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_233),
.B(n_127),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_264),
.A2(n_177),
.B1(n_149),
.B2(n_172),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_242),
.B(n_172),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_338),
.B(n_295),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_231),
.A2(n_132),
.B1(n_177),
.B2(n_190),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_339),
.A2(n_268),
.B1(n_223),
.B2(n_247),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_220),
.A2(n_190),
.B1(n_183),
.B2(n_188),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_341),
.A2(n_290),
.B(n_335),
.Y(n_376)
);

INVx13_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_345),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_243),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_347),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_173),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_313),
.A2(n_219),
.B1(n_217),
.B2(n_260),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_350),
.A2(n_366),
.B1(n_370),
.B2(n_374),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_317),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_351),
.B(n_353),
.Y(n_392)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_296),
.B(n_227),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_355),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_319),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_357),
.C(n_331),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_337),
.B(n_311),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_219),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_365),
.C(n_385),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_328),
.B(n_227),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_361),
.Y(n_402)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_293),
.Y(n_360)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_360),
.Y(n_420)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_326),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_362),
.A2(n_341),
.B1(n_327),
.B2(n_322),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_244),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_363),
.B(n_364),
.Y(n_413)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_299),
.B(n_224),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_244),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_371),
.Y(n_417)
);

INVx13_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_369),
.Y(n_416)
);

INVx13_ASAP7_75t_L g370 ( 
.A(n_302),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_336),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_373),
.A2(n_376),
.B(n_381),
.Y(n_391)
);

INVx13_ASAP7_75t_L g374 ( 
.A(n_302),
.Y(n_374)
);

AND2x6_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_249),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_375),
.B(n_378),
.Y(n_394)
);

AND2x2_ASAP7_75t_SL g377 ( 
.A(n_332),
.B(n_229),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_288),
.C(n_308),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_246),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_380),
.Y(n_400)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_301),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_301),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_383),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_289),
.A2(n_238),
.B1(n_284),
.B2(n_253),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_289),
.A2(n_235),
.B1(n_232),
.B2(n_251),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_333),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_304),
.B(n_285),
.C(n_249),
.Y(n_385)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_386),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_373),
.A2(n_304),
.B(n_303),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_387),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_388),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_367),
.A2(n_320),
.B1(n_305),
.B2(n_310),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_396),
.A2(n_409),
.B1(n_421),
.B2(n_372),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_348),
.B(n_303),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_398),
.B(n_384),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_399),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_348),
.A2(n_288),
.B(n_308),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_408),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_342),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_407),
.C(n_415),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_410),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_367),
.B(n_342),
.C(n_309),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_367),
.A2(n_333),
.B1(n_330),
.B2(n_336),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_356),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_330),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_346),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_344),
.A2(n_297),
.B(n_307),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_412),
.A2(n_387),
.B(n_391),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_358),
.B(n_298),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_346),
.A2(n_314),
.B1(n_322),
.B2(n_315),
.Y(n_421)
);

INVx13_ASAP7_75t_L g423 ( 
.A(n_416),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_423),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_389),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_425),
.B(n_345),
.Y(n_482)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_392),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_416),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_431),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_357),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_428),
.B(n_438),
.Y(n_455)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_429),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_394),
.A2(n_383),
.B1(n_376),
.B2(n_372),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_430),
.A2(n_445),
.B1(n_447),
.B2(n_436),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_411),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_355),
.Y(n_432)
);

OAI21xp33_ASAP7_75t_L g466 ( 
.A1(n_432),
.A2(n_434),
.B(n_435),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_393),
.B(n_354),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_380),
.Y(n_435)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_382),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_377),
.Y(n_439)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_404),
.A2(n_394),
.B1(n_409),
.B2(n_396),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_440),
.A2(n_419),
.B1(n_418),
.B2(n_399),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_389),
.B(n_385),
.C(n_377),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_403),
.C(n_415),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_377),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_442),
.B(n_443),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_400),
.B(n_379),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_352),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_444),
.B(n_420),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_404),
.A2(n_372),
.B1(n_375),
.B2(n_362),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_447),
.B(n_420),
.Y(n_481)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_448),
.Y(n_464)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_450),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_371),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_452),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_400),
.B(n_360),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_453),
.A2(n_449),
.B(n_391),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_454),
.A2(n_462),
.B(n_468),
.Y(n_496)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_459),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_460),
.A2(n_461),
.B1(n_446),
.B2(n_433),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_388),
.B1(n_408),
.B2(n_407),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_453),
.A2(n_412),
.B(n_344),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_440),
.A2(n_402),
.B(n_417),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_438),
.Y(n_469)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_469),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_431),
.B(n_452),
.Y(n_472)
);

NOR2x1_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_442),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_473),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_424),
.B(n_417),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_474),
.B(n_478),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_422),
.C(n_441),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_443),
.B(n_398),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_477),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_437),
.B(n_413),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_434),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_479),
.A2(n_433),
.B1(n_439),
.B2(n_445),
.Y(n_484)
);

AO22x1_ASAP7_75t_SL g480 ( 
.A1(n_437),
.A2(n_366),
.B1(n_399),
.B2(n_421),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_437),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_481),
.B(n_425),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_482),
.B(n_422),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_483),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_484),
.A2(n_485),
.B1(n_492),
.B2(n_488),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_479),
.A2(n_465),
.B1(n_460),
.B2(n_461),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_485),
.A2(n_490),
.B1(n_492),
.B2(n_493),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_486),
.B(n_487),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_454),
.A2(n_446),
.B(n_432),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_497),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_498),
.C(n_503),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_465),
.A2(n_433),
.B1(n_427),
.B2(n_435),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_468),
.A2(n_451),
.B1(n_444),
.B2(n_448),
.Y(n_493)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

FAx1_ASAP7_75t_SL g497 ( 
.A(n_476),
.B(n_450),
.CI(n_429),
.CON(n_497),
.SN(n_497)
);

MAJIxp5_ASAP7_75t_SL g498 ( 
.A(n_481),
.B(n_423),
.C(n_374),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_298),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_499),
.B(n_505),
.Y(n_518)
);

AO21x1_ASAP7_75t_L g501 ( 
.A1(n_470),
.A2(n_423),
.B(n_395),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_501),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_470),
.C(n_477),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_456),
.B(n_345),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_315),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_506),
.B(n_480),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_455),
.B(n_361),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_507),
.B(n_463),
.Y(n_520)
);

XNOR2x1_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_523),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_500),
.A2(n_457),
.B1(n_469),
.B2(n_472),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_513),
.A2(n_495),
.B1(n_503),
.B2(n_506),
.Y(n_528)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_501),
.Y(n_515)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_515),
.Y(n_533)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_494),
.Y(n_516)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_516),
.Y(n_536)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_504),
.Y(n_517)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_517),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_484),
.A2(n_457),
.B1(n_462),
.B2(n_480),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_520),
.Y(n_529)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_502),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_526),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_487),
.B(n_471),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_524),
.B(n_486),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_505),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_491),
.A2(n_480),
.B1(n_471),
.B2(n_467),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_527),
.B(n_464),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_528),
.A2(n_532),
.B1(n_534),
.B2(n_535),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_499),
.C(n_489),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_530),
.B(n_521),
.C(n_518),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_511),
.A2(n_496),
.B(n_483),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_511),
.A2(n_467),
.B1(n_463),
.B2(n_458),
.Y(n_534)
);

AOI221xp5_ASAP7_75t_L g535 ( 
.A1(n_516),
.A2(n_497),
.B1(n_496),
.B2(n_498),
.C(n_458),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_510),
.A2(n_497),
.B1(n_464),
.B2(n_463),
.Y(n_537)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_537),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_539),
.B(n_521),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_541),
.B(n_515),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_509),
.B(n_390),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_542),
.B(n_543),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_517),
.B(n_395),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_544),
.B(n_546),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_545),
.B(n_551),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_533),
.A2(n_514),
.B1(n_525),
.B2(n_527),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_508),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_547),
.A2(n_549),
.B(n_543),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_536),
.B(n_512),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_540),
.B(n_390),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_550),
.B(n_554),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_540),
.B(n_518),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_529),
.A2(n_519),
.B1(n_524),
.B2(n_523),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_555),
.B(n_556),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_529),
.A2(n_386),
.B1(n_364),
.B2(n_314),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_553),
.B(n_531),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_557),
.B(n_548),
.C(n_545),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_552),
.A2(n_532),
.B(n_541),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_562),
.Y(n_568)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_561),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_544),
.A2(n_530),
.B(n_531),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_551),
.A2(n_539),
.B(n_537),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_563),
.A2(n_364),
.B1(n_386),
.B2(n_326),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_548),
.B(n_538),
.C(n_307),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_565),
.B(n_566),
.Y(n_574)
);

XOR2x2_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_374),
.Y(n_566)
);

NOR3xp33_ASAP7_75t_L g569 ( 
.A(n_558),
.B(n_544),
.C(n_546),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_569),
.B(n_570),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_564),
.B(n_343),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_571),
.B(n_572),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_334),
.C(n_292),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_565),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_576),
.B(n_577),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_573),
.B(n_560),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_568),
.B(n_557),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_579),
.A2(n_569),
.B(n_574),
.Y(n_581)
);

OAI321xp33_ASAP7_75t_L g585 ( 
.A1(n_581),
.A2(n_582),
.A3(n_369),
.B1(n_370),
.B2(n_334),
.C(n_340),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_580),
.A2(n_560),
.B(n_566),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_583),
.A2(n_578),
.B1(n_306),
.B2(n_340),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_584),
.A2(n_585),
.B1(n_306),
.B2(n_369),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_586),
.A2(n_370),
.B1(n_343),
.B2(n_292),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_587),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_588),
.B(n_216),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_589),
.B(n_228),
.Y(n_590)
);


endmodule