module fake_jpeg_16927_n_112 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_112);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_12),
.B(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_20),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_20),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_40),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_27),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_22),
.A2(n_14),
.B1(n_15),
.B2(n_12),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_21),
.B1(n_13),
.B2(n_2),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_19),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_50),
.B1(n_37),
.B2(n_21),
.Y(n_61)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_23),
.B(n_29),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_53),
.C(n_50),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_22),
.B1(n_30),
.B2(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_55),
.B1(n_54),
.B2(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_13),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_39),
.B1(n_37),
.B2(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_63),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_31),
.B1(n_37),
.B2(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_46),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_57),
.C(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_73),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_62),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_64),
.C(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_81),
.B1(n_82),
.B2(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_62),
.B1(n_47),
.B2(n_51),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_44),
.B1(n_65),
.B2(n_50),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_84),
.A2(n_86),
.B(n_68),
.C(n_3),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_2),
.B(n_3),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_91),
.B(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_58),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_3),
.B(n_4),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_4),
.C(n_5),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_6),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_96),
.Y(n_99)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_83),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_80),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_102),
.B(n_80),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_88),
.B(n_81),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_106),
.C(n_105),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_99),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_79),
.C(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_108),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_88),
.A3(n_45),
.B1(n_58),
.B2(n_9),
.C1(n_6),
.C2(n_11),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_7),
.B(n_8),
.Y(n_111)
);

AOI21x1_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_110),
.B(n_10),
.Y(n_112)
);


endmodule