module real_jpeg_32392_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_249;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_210;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_283;
wire n_85;
wire n_81;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

AOI22x1_ASAP7_75t_L g43 ( 
.A1(n_0),
.A2(n_23),
.B1(n_44),
.B2(n_48),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_0),
.A2(n_23),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_0),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_0),
.B(n_75),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_0),
.A2(n_139),
.A3(n_145),
.B1(n_148),
.B2(n_157),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_0),
.A2(n_23),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_0),
.B(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_2),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_2),
.Y(n_254)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_3),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_6),
.Y(n_218)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_8),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_70),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

OAI22x1_ASAP7_75t_SL g186 ( 
.A1(n_8),
.A2(n_70),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_8),
.A2(n_70),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_9),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_9),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_221),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

AOI21x1_ASAP7_75t_SL g12 ( 
.A1(n_13),
.A2(n_195),
.B(n_220),
.Y(n_12)
);

OAI21x1_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_134),
.B(n_194),
.Y(n_13)
);

AOI21x1_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_112),
.B(n_133),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_76),
.Y(n_15)
);

NOR2xp67_ASAP7_75t_SL g133 ( 
.A(n_16),
.B(n_76),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_40),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_17),
.A2(n_40),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_17),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_24),
.B(n_29),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_23),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_30),
.B(n_35),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_23),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_23),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_23),
.B(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_23),
.A2(n_252),
.B(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_54),
.B(n_58),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_35),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_58)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_40),
.A2(n_121),
.B1(n_167),
.B2(n_193),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_40),
.B(n_137),
.C(n_193),
.Y(n_196)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22x1_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_53),
.B1(n_65),
.B2(n_75),
.Y(n_41)
);

AOI22x1_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_53),
.B1(n_75),
.B2(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_43),
.Y(n_285)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_47),
.Y(n_147)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_52),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_54),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_58),
.B(n_282),
.C(n_283),
.Y(n_281)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_97),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_77),
.B(n_98),
.C(n_102),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_77),
.B(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_130),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_85),
.B1(n_89),
.B2(n_93),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_80),
.B(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_93),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_98),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_98),
.B(n_200),
.C(n_202),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_99),
.Y(n_201)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g168 ( 
.A(n_103),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_103),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_103),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21x1_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_122),
.B(n_132),
.Y(n_112)
);

NOR2xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_119),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_114),
.B(n_203),
.C(n_210),
.Y(n_256)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_115),
.A2(n_210),
.B(n_219),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

OAI211xp5_ASAP7_75t_L g219 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.C(n_210),
.Y(n_219)
);

AOI21x1_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_129),
.B(n_131),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_136),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_166),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_163),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

BUFx4f_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_167),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_167),
.A2(n_193),
.B1(n_280),
.B2(n_286),
.Y(n_279)
);

AOI22x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_181),
.B1(n_186),
.B2(n_192),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_168),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_173),
.B1(n_176),
.B2(n_178),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_184),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_186),
.Y(n_205)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx4f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_197),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_208),
.B2(n_209),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_211),
.B(n_273),
.Y(n_272)
);

AO22x1_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_217),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_214),
.Y(n_276)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_287),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_224),
.B(n_225),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_257),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_255),
.B2(n_256),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21x1_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_233),
.B(n_243),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_240),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_273)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_279),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B(n_268),
.Y(n_260)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);


endmodule