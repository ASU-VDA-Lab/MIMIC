module fake_jpeg_1504_n_236 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_236);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_235;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_27),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_83),
.Y(n_96)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_52),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_54),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_76),
.B1(n_56),
.B2(n_67),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_68),
.B1(n_64),
.B2(n_73),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_100),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_78),
.Y(n_101)
);

AO22x1_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_85),
.B1(n_86),
.B2(n_68),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_116),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_112),
.Y(n_132)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_83),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_122),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_76),
.B1(n_79),
.B2(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_121),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_87),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_87),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_120),
.B1(n_73),
.B2(n_72),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_73),
.B(n_64),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_66),
.B1(n_59),
.B2(n_67),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_63),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_82),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_79),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_125),
.C(n_42),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_53),
.C(n_66),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_57),
.A3(n_74),
.B1(n_61),
.B2(n_69),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_140),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_129),
.A2(n_142),
.B1(n_5),
.B2(n_6),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_1),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_134),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_1),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_144),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_59),
.B1(n_94),
.B2(n_65),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_58),
.B1(n_57),
.B2(n_22),
.Y(n_158)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_104),
.B(n_103),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_65),
.B1(n_58),
.B2(n_57),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_5),
.B(n_6),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_107),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_143),
.Y(n_152)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_157),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_94),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_2),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_111),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_14),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_25),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_163),
.Y(n_186)
);

OAI211xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_167),
.B(n_10),
.C(n_12),
.Y(n_177)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_3),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_125),
.B1(n_137),
.B2(n_135),
.Y(n_164)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_124),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_8),
.Y(n_170)
);

AOI22x1_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_29),
.B1(n_50),
.B2(n_49),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_33),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_8),
.C(n_9),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_180),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_30),
.B(n_47),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_176),
.B(n_187),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_51),
.B(n_46),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_187),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_45),
.B(n_44),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_13),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_189),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_192),
.A2(n_160),
.B1(n_159),
.B2(n_158),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_198),
.Y(n_206)
);

AO221x1_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_165),
.B1(n_146),
.B2(n_153),
.C(n_160),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_201),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_183),
.A2(n_167),
.B(n_161),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_189),
.B1(n_183),
.B2(n_178),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_200),
.B1(n_186),
.B2(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_179),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_198),
.A2(n_176),
.B(n_174),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_207),
.B(n_210),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_171),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_195),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_211),
.B(n_214),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_200),
.B1(n_204),
.B2(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_172),
.C(n_190),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_190),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_205),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_216),
.A2(n_218),
.B1(n_209),
.B2(n_197),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_208),
.B(n_215),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_210),
.B1(n_203),
.B2(n_19),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_219),
.B1(n_225),
.B2(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_219),
.Y(n_230)
);

NOR2xp67_ASAP7_75t_SL g231 ( 
.A(n_230),
.B(n_228),
.Y(n_231)
);

AOI21x1_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_221),
.B(n_226),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_222),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_35),
.B(n_36),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_234),
.A2(n_38),
.B(n_17),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_16),
.Y(n_236)
);


endmodule