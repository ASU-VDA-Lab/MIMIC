module fake_jpeg_17815_n_390 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx2_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_40),
.B(n_47),
.Y(n_109)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_37),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_56),
.B(n_31),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_104),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_38),
.A2(n_18),
.B1(n_29),
.B2(n_26),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_68),
.A2(n_90),
.B1(n_93),
.B2(n_16),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_29),
.B1(n_18),
.B2(n_37),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_94),
.B(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_73),
.B(n_78),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_84),
.B(n_102),
.Y(n_162)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_28),
.Y(n_88)
);

OR2x2_ASAP7_75t_SL g152 ( 
.A(n_88),
.B(n_95),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_46),
.A2(n_18),
.B1(n_29),
.B2(n_26),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_18),
.B1(n_28),
.B2(n_23),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_48),
.B(n_14),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_42),
.B(n_36),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_39),
.A2(n_36),
.B1(n_35),
.B2(n_33),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_35),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_111),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_58),
.A2(n_32),
.B1(n_27),
.B2(n_24),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_6),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_33),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_41),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_64),
.A2(n_32),
.B1(n_27),
.B2(n_24),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_61),
.A2(n_24),
.B(n_20),
.C(n_16),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_17),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_120),
.A2(n_169),
.B1(n_142),
.B2(n_166),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_70),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_123),
.B(n_125),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_69),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_17),
.C(n_20),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_164),
.C(n_89),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_20),
.Y(n_130)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_139),
.Y(n_212)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_78),
.A2(n_0),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_9),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_99),
.A2(n_16),
.B1(n_4),
.B2(n_5),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_148),
.B1(n_165),
.B2(n_124),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_147),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_151),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_1),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_150),
.A2(n_169),
.B(n_121),
.Y(n_215)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_112),
.B(n_5),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_155),
.B(n_161),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_156),
.Y(n_206)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_165),
.Y(n_186)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_5),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_94),
.B(n_6),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

BUFx8_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_87),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_90),
.B(n_6),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_170),
.A2(n_179),
.B1(n_185),
.B2(n_199),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_173),
.A2(n_195),
.B1(n_148),
.B2(n_142),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_116),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_180),
.Y(n_216)
);

OAI22x1_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_100),
.B1(n_89),
.B2(n_116),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_107),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_137),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_119),
.A2(n_82),
.B1(n_107),
.B2(n_80),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_101),
.B1(n_92),
.B2(n_10),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_92),
.C(n_87),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_132),
.C(n_158),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_191),
.B(n_193),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_192),
.B(n_194),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_12),
.Y(n_193)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_127),
.B(n_10),
.CI(n_11),
.CON(n_194),
.SN(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_119),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_169),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_198),
.B(n_201),
.Y(n_252)
);

OAI22x1_ASAP7_75t_SL g199 ( 
.A1(n_152),
.A2(n_11),
.B1(n_12),
.B2(n_120),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_11),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_SL g250 ( 
.A1(n_205),
.A2(n_197),
.B(n_187),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_152),
.B(n_120),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_208),
.A2(n_201),
.B(n_180),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_120),
.B(n_128),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_214),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_122),
.B(n_134),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_215),
.B(n_201),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_199),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_217),
.B(n_219),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_174),
.C(n_213),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_218),
.B(n_256),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_214),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_235),
.B1(n_254),
.B2(n_256),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_186),
.A2(n_138),
.B1(n_157),
.B2(n_153),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_221),
.A2(n_224),
.B1(n_251),
.B2(n_226),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_202),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_224),
.C(n_251),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_181),
.A2(n_160),
.B1(n_131),
.B2(n_139),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_131),
.Y(n_225)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_179),
.A2(n_140),
.B(n_137),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_229),
.A2(n_228),
.B(n_221),
.C(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_223),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_208),
.B(n_193),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_233),
.A2(n_241),
.B(n_248),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_132),
.B1(n_156),
.B2(n_191),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_242),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_176),
.B(n_175),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_171),
.Y(n_239)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_253),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_184),
.B(n_195),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_205),
.A2(n_194),
.A3(n_203),
.B1(n_189),
.B2(n_192),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_171),
.B(n_177),
.Y(n_243)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_188),
.B1(n_190),
.B2(n_194),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_250),
.B1(n_226),
.B2(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_172),
.Y(n_246)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_188),
.A2(n_190),
.B(n_204),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_197),
.B(n_187),
.C(n_211),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_231),
.C(n_233),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_182),
.A2(n_213),
.B1(n_159),
.B2(n_146),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_206),
.B(n_182),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_206),
.A2(n_208),
.B1(n_170),
.B2(n_159),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_171),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_234),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_254),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_259),
.A2(n_265),
.B1(n_278),
.B2(n_229),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_227),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_264),
.B(n_266),
.Y(n_309)
);

NAND2x1_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_244),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_267),
.B(n_252),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_228),
.B1(n_241),
.B2(n_229),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_216),
.B(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_220),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_230),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_277),
.B(n_288),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_219),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_231),
.C(n_232),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_237),
.Y(n_282)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_287),
.B(n_252),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_255),
.B1(n_247),
.B2(n_234),
.Y(n_300)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_234),
.Y(n_290)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_300),
.B1(n_319),
.B2(n_288),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_296),
.B1(n_259),
.B2(n_262),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_294),
.A2(n_283),
.B1(n_289),
.B2(n_280),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_297),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_229),
.B1(n_222),
.B2(n_240),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_285),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_290),
.Y(n_302)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_286),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_279),
.C(n_280),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_305),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_257),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_308),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_257),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_271),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_261),
.B(n_260),
.Y(n_313)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_284),
.Y(n_314)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_263),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_263),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_316),
.Y(n_330)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_318),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_274),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_322),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_321),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_282),
.C(n_287),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_326),
.A2(n_327),
.B1(n_316),
.B2(n_306),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_294),
.A2(n_289),
.B1(n_259),
.B2(n_265),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_273),
.C(n_276),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_289),
.C(n_275),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_335),
.C(n_339),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_275),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_333),
.A2(n_312),
.B(n_310),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_300),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_311),
.C(n_305),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_297),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_340),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_317),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_341),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_342),
.B(n_320),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_303),
.Y(n_344)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_345),
.A2(n_351),
.B(n_354),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_325),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_350),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_293),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_356),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_326),
.A2(n_308),
.B1(n_307),
.B2(n_296),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_348),
.A2(n_331),
.B1(n_327),
.B2(n_318),
.Y(n_367)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_352),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_317),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_329),
.A2(n_311),
.B(n_303),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_329),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_309),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_353),
.A2(n_330),
.B1(n_337),
.B2(n_339),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_358),
.A2(n_354),
.B1(n_352),
.B2(n_342),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_365),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_367),
.B(n_368),
.Y(n_373)
);

AO221x1_ASAP7_75t_L g368 ( 
.A1(n_345),
.A2(n_331),
.B1(n_328),
.B2(n_323),
.C(n_295),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_359),
.A2(n_355),
.B(n_349),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_369),
.A2(n_359),
.B(n_343),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_347),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_372),
.C(n_355),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_356),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_361),
.B(n_348),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_374),
.B(n_375),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_360),
.Y(n_376)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_376),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_377),
.A2(n_363),
.B1(n_364),
.B2(n_370),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_372),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_380),
.B(n_381),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_362),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_383),
.A2(n_380),
.B(n_370),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_384),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_371),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_387),
.Y(n_388)
);

AOI221xp5_ASAP7_75t_L g389 ( 
.A1(n_388),
.A2(n_366),
.B1(n_363),
.B2(n_378),
.C(n_351),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_367),
.Y(n_390)
);


endmodule