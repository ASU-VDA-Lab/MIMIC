module fake_jpeg_8609_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx8_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_9),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_21),
.B1(n_15),
.B2(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_19),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_21),
.B1(n_17),
.B2(n_8),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_1),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_19),
.B(n_8),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_28),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_16),
.B(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OA21x2_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_35),
.B(n_20),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_20),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_25),
.B1(n_20),
.B2(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_17),
.B1(n_25),
.B2(n_18),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_20),
.Y(n_45)
);

MAJx2_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_18),
.C(n_14),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_41),
.B(n_20),
.Y(n_46)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_26),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_46),
.B(n_47),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_26),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_4),
.C(n_6),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_48),
.B1(n_26),
.B2(n_3),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_2),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_3),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_57),
.CI(n_54),
.CON(n_58),
.SN(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_53),
.C(n_55),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_58),
.Y(n_60)
);


endmodule