module fake_jpeg_18541_n_212 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_25),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_32),
.Y(n_47)
);

AND2x4_ASAP7_75t_SL g27 ( 
.A(n_18),
.B(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_6),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_24),
.Y(n_51)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_49),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_47),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_54),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_27),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_28),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_31),
.B1(n_32),
.B2(n_27),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_59),
.B1(n_42),
.B2(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_31),
.B1(n_27),
.B2(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_42),
.B1(n_36),
.B2(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_26),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_61),
.B1(n_41),
.B2(n_56),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_40),
.B(n_60),
.C(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_73),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_81),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_33),
.A3(n_25),
.B1(n_42),
.B2(n_14),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_52),
.B(n_49),
.C(n_48),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_82),
.C(n_52),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_36),
.B1(n_26),
.B2(n_37),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_62),
.B1(n_41),
.B2(n_37),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_46),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_88),
.B(n_95),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_89),
.Y(n_110)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_86),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_52),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_70),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_98),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_61),
.B1(n_41),
.B2(n_44),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_72),
.C(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_73),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_107),
.B(n_109),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_112),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_81),
.B1(n_97),
.B2(n_61),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_58),
.B1(n_14),
.B2(n_15),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_84),
.B(n_94),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_111),
.B(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_96),
.B1(n_91),
.B2(n_82),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_131),
.B1(n_114),
.B2(n_115),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_113),
.A2(n_84),
.B1(n_72),
.B2(n_76),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_105),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_84),
.B1(n_88),
.B2(n_74),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_85),
.B1(n_97),
.B2(n_69),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_129),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_81),
.B1(n_46),
.B2(n_35),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_106),
.B1(n_108),
.B2(n_104),
.Y(n_137)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_16),
.Y(n_149)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_21),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_144),
.B1(n_149),
.B2(n_150),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_143),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_145),
.Y(n_152)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_58),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_15),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_118),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_12),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_128),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_46),
.B1(n_28),
.B2(n_13),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_116),
.C(n_119),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_155),
.C(n_150),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_125),
.C(n_124),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_133),
.C(n_123),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_129),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_19),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_162),
.A2(n_136),
.B1(n_137),
.B2(n_148),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_169),
.B1(n_160),
.B2(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_149),
.B1(n_143),
.B2(n_140),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_172),
.C(n_152),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_174),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_173),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_28),
.B1(n_8),
.B2(n_9),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_176),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_19),
.B1(n_6),
.B2(n_11),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_152),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_170),
.C(n_171),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_8),
.B(n_10),
.C(n_9),
.D(n_3),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_7),
.C(n_11),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_12),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_188),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_166),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_193),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_23),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_192),
.Y(n_200)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_4),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_0),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_181),
.A3(n_184),
.B1(n_180),
.B2(n_186),
.C1(n_183),
.C2(n_20),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_197),
.B(n_199),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_187),
.B1(n_5),
.B2(n_3),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_4),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.C(n_195),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_5),
.B(n_8),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_205),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_201),
.A2(n_5),
.B(n_23),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_1),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_2),
.B(n_209),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_2),
.Y(n_212)
);


endmodule