module fake_jpeg_25182_n_250 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_30),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_14),
.B1(n_17),
.B2(n_23),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_35),
.B1(n_14),
.B2(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_14),
.B1(n_23),
.B2(n_17),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_13),
.B(n_12),
.C(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_52),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_25),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_33),
.B1(n_17),
.B2(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_32),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_60),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_67),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_40),
.B1(n_38),
.B2(n_13),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_27),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_40),
.B1(n_39),
.B2(n_16),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_63),
.B(n_72),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_36),
.B(n_60),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_94),
.B1(n_76),
.B2(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_59),
.B(n_39),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_62),
.B(n_78),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_69),
.B1(n_75),
.B2(n_78),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_71),
.B(n_77),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_60),
.B1(n_33),
.B2(n_54),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_29),
.C(n_26),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_26),
.C(n_29),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_26),
.B(n_32),
.C(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_68),
.B1(n_76),
.B2(n_65),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_107),
.B(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_102),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_113),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_86),
.B(n_91),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_71),
.A3(n_72),
.B1(n_74),
.B2(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_88),
.C(n_86),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_62),
.B1(n_68),
.B2(n_76),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_115),
.B1(n_82),
.B2(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_85),
.B(n_22),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_84),
.A2(n_65),
.B1(n_32),
.B2(n_24),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_116),
.B(n_132),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_93),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_118),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_87),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_123),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_94),
.B1(n_92),
.B2(n_96),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_126),
.B1(n_30),
.B2(n_50),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_127),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_107),
.B1(n_99),
.B2(n_111),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_104),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_133),
.C(n_136),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_81),
.C(n_92),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_81),
.B(n_82),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_79),
.B(n_50),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_20),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_143),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_101),
.B1(n_112),
.B2(n_102),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_149),
.B1(n_15),
.B2(n_21),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_113),
.C(n_97),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_146),
.C(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_152),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_97),
.C(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_148),
.B(n_156),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_79),
.Y(n_148)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_49),
.C(n_30),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_47),
.C(n_19),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_130),
.C(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_158),
.Y(n_169)
);

XOR2x2_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_22),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_157),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_162),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_10),
.B(n_1),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_118),
.C(n_120),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_153),
.C(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_168),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_125),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_119),
.B1(n_136),
.B2(n_47),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_174),
.B1(n_160),
.B2(n_168),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_24),
.B1(n_10),
.B2(n_19),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_156),
.B1(n_146),
.B2(n_154),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_144),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_186),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_157),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_21),
.C(n_24),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_16),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_193),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_24),
.B1(n_21),
.B2(n_15),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_191),
.B(n_1),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_0),
.B(n_1),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_192),
.A2(n_170),
.B1(n_173),
.B2(n_172),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_15),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_173),
.B(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

NOR2x1_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_204),
.B1(n_186),
.B2(n_193),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_170),
.B1(n_165),
.B2(n_172),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_184),
.B1(n_183),
.B2(n_180),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_204),
.Y(n_207)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_2),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_172),
.B1(n_21),
.B2(n_3),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_1),
.B(n_2),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_183),
.C(n_3),
.Y(n_211)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_210),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_215),
.B1(n_2),
.B2(n_4),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_2),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_214),
.C(n_216),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_9),
.C(n_4),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_9),
.C(n_4),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_200),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_195),
.C(n_201),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_212),
.A2(n_197),
.B1(n_199),
.B2(n_196),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_213),
.B1(n_6),
.B2(n_7),
.Y(n_228)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_5),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_226),
.C(n_216),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_202),
.B(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_223),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_224),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_4),
.C(n_5),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_219),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_222),
.C(n_225),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_5),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_233),
.B(n_234),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_6),
.B(n_7),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_238),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_232),
.B(n_219),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_223),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_239),
.A2(n_230),
.B(n_231),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_240),
.A2(n_242),
.B(n_235),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_226),
.B(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_244),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_241),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_245),
.A2(n_6),
.B(n_8),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_8),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_247),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_8),
.B(n_9),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_8),
.B(n_9),
.Y(n_250)
);


endmodule