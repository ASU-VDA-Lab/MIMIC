module fake_jpeg_24084_n_62 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_38;
wire n_36;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_1),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_37),
.B(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_0),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_44),
.B(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_19),
.B1(n_6),
.B2(n_7),
.Y(n_49)
);

AOI211xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_42),
.B(n_2),
.C(n_10),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_8),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_55),
.B(n_56),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_52),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_50),
.C(n_24),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_23),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_27),
.Y(n_62)
);


endmodule