module fake_jpeg_30729_n_360 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_360);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx11_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_48),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_59),
.Y(n_96)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_6),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_6),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_67),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_64),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_26),
.B(n_5),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_30),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_73),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_21),
.B(n_35),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_16),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_69),
.B1(n_60),
.B2(n_74),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_77),
.A2(n_90),
.B1(n_116),
.B2(n_0),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_28),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_92),
.B(n_113),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_30),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_28),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_1),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_40),
.B(n_38),
.C(n_35),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_42),
.B(n_72),
.C(n_2),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_41),
.B1(n_36),
.B2(n_43),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_30),
.B1(n_32),
.B2(n_42),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_117),
.B1(n_42),
.B2(n_31),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_32),
.CON(n_92),
.SN(n_92)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_70),
.B(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_115),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_41),
.B1(n_23),
.B2(n_43),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_97),
.A2(n_98),
.B1(n_118),
.B2(n_9),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_45),
.A2(n_41),
.B1(n_23),
.B2(n_39),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_38),
.B(n_40),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_9),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_121),
.Y(n_123)
);

HAxp5_ASAP7_75t_SL g113 ( 
.A(n_55),
.B(n_39),
.CON(n_113),
.SN(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_19),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_47),
.B(n_33),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_49),
.A2(n_19),
.B1(n_33),
.B2(n_31),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_68),
.A2(n_42),
.B1(n_31),
.B2(n_2),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_42),
.B1(n_31),
.B2(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_45),
.B(n_7),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_122),
.A2(n_86),
.B1(n_88),
.B2(n_94),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_133),
.Y(n_168)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_127),
.A2(n_130),
.B(n_140),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_5),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_78),
.B(n_0),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_138),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_92),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_157),
.B1(n_106),
.B2(n_108),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_146),
.Y(n_169)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_78),
.B(n_7),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_76),
.Y(n_165)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_78),
.B(n_7),
.C(n_8),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_80),
.B(n_8),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_159),
.Y(n_166)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_9),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_150),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_107),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_93),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_161),
.Y(n_173)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_84),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_94),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_119),
.B1(n_108),
.B2(n_88),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_163),
.A2(n_164),
.B1(n_175),
.B2(n_187),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_89),
.B1(n_113),
.B2(n_110),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_165),
.B(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_159),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_116),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_119),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_136),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_129),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_198),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_131),
.B(n_86),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_189),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_142),
.B1(n_124),
.B2(n_147),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_128),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_188),
.A2(n_156),
.B1(n_155),
.B2(n_154),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_123),
.B(n_104),
.Y(n_196)
);

NAND2x1_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_139),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_204),
.A2(n_209),
.B1(n_186),
.B2(n_197),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_136),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_211),
.C(n_220),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_206),
.B(n_207),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_173),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_139),
.B1(n_145),
.B2(n_148),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_194),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_210),
.B(n_214),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_144),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_166),
.B(n_144),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_216),
.B(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_170),
.B(n_146),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_227),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_177),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_151),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_160),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_158),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_225),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_169),
.B(n_126),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_139),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_175),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_182),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_188),
.B(n_132),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_232),
.B(n_178),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_192),
.B(n_182),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_235),
.B(n_245),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_163),
.B(n_181),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_177),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_243),
.B(n_244),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_174),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_180),
.B(n_165),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_250),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_165),
.B1(n_195),
.B2(n_197),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_231),
.A3(n_202),
.B1(n_203),
.B2(n_229),
.C1(n_211),
.C2(n_205),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_258),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_200),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_231),
.A2(n_195),
.B1(n_165),
.B2(n_186),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_204),
.B1(n_216),
.B2(n_185),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_210),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_230),
.Y(n_263)
);

OAI32xp33_ASAP7_75t_L g258 ( 
.A1(n_203),
.A2(n_206),
.A3(n_232),
.B1(n_202),
.B2(n_220),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_200),
.B(n_174),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_246),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_200),
.C(n_217),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_277),
.C(n_261),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_270),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_224),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_259),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_236),
.A2(n_201),
.B1(n_222),
.B2(n_215),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_272),
.A2(n_276),
.B1(n_260),
.B2(n_251),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_237),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_274),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_223),
.B(n_208),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_279),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_199),
.C(n_178),
.Y(n_277)
);

NAND4xp25_ASAP7_75t_SL g278 ( 
.A(n_239),
.B(n_135),
.C(n_183),
.D(n_190),
.Y(n_278)
);

NAND4xp25_ASAP7_75t_SL g295 ( 
.A(n_278),
.B(n_249),
.C(n_256),
.D(n_247),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_199),
.Y(n_280)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_280),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_234),
.B(n_183),
.Y(n_281)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_257),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

AO22x1_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_235),
.B1(n_258),
.B2(n_248),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_268),
.B(n_266),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_277),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_297),
.C(n_301),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_295),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_249),
.C(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_245),
.C(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_262),
.B(n_257),
.C(n_260),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_282),
.B1(n_268),
.B2(n_270),
.Y(n_304)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_263),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_269),
.B1(n_267),
.B2(n_283),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_304),
.A2(n_307),
.B1(n_308),
.B2(n_314),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_265),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_314),
.Y(n_323)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_286),
.B1(n_289),
.B2(n_303),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_308),
.A2(n_298),
.B1(n_288),
.B2(n_292),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_311),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_289),
.A2(n_280),
.B1(n_266),
.B2(n_279),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_310),
.A2(n_318),
.B1(n_295),
.B2(n_298),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_264),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_285),
.B1(n_292),
.B2(n_294),
.Y(n_313)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_275),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_293),
.C(n_299),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_285),
.A2(n_276),
.B1(n_273),
.B2(n_241),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_312),
.B(n_294),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_328),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_324),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_300),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_322),
.Y(n_336)
);

XNOR2x1_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_301),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_329),
.Y(n_339)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_330),
.A2(n_317),
.B(n_309),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g331 ( 
.A(n_323),
.B(n_316),
.CI(n_304),
.CON(n_331),
.SN(n_331)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_333),
.Y(n_342)
);

AOI31xp67_ASAP7_75t_SL g333 ( 
.A1(n_320),
.A2(n_293),
.A3(n_299),
.B(n_278),
.Y(n_333)
);

NAND4xp25_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_317),
.C(n_238),
.D(n_305),
.Y(n_334)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_334),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_338),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_325),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_321),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_328),
.A2(n_318),
.B(n_241),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_339),
.B(n_327),
.C(n_330),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_343),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_327),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_323),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_347),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_238),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_348),
.B(n_176),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_331),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_344),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_352),
.B(n_353),
.C(n_343),
.Y(n_356)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_350),
.A2(n_342),
.B(n_344),
.C(n_346),
.Y(n_354)
);

AOI21x1_ASAP7_75t_L g358 ( 
.A1(n_354),
.A2(n_338),
.B(n_190),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_349),
.B(n_341),
.Y(n_357)
);

OAI311xp33_ASAP7_75t_L g359 ( 
.A1(n_357),
.A2(n_358),
.A3(n_355),
.B1(n_176),
.C1(n_143),
.Y(n_359)
);

XNOR2x2_ASAP7_75t_SL g360 ( 
.A(n_359),
.B(n_134),
.Y(n_360)
);


endmodule