module real_jpeg_27944_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_0),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_0),
.A2(n_28),
.B1(n_54),
.B2(n_56),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_0),
.A2(n_28),
.B1(n_60),
.B2(n_61),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_54),
.Y(n_92)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_1),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_107),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_2),
.A2(n_54),
.B1(n_56),
.B2(n_107),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_107),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_3),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_49),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_6),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_6),
.A2(n_30),
.B(n_34),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_120),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_6),
.B(n_32),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_6),
.A2(n_60),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_6),
.B(n_60),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_6),
.B(n_74),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_6),
.A2(n_91),
.B1(n_246),
.B2(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_6),
.A2(n_33),
.B(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_7),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_105),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_7),
.A2(n_60),
.B1(n_61),
.B2(n_105),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_7),
.A2(n_54),
.B1(n_56),
.B2(n_105),
.Y(n_240)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_9),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_9),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_10),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_110),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_110),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_54),
.B1(n_56),
.B2(n_110),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_11),
.A2(n_60),
.B1(n_61),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_11),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_100),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_100),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_11),
.A2(n_54),
.B1(n_56),
.B2(n_100),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_12),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_12),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_12),
.A2(n_56),
.A3(n_60),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_13),
.A2(n_37),
.B1(n_60),
.B2(n_61),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_13),
.A2(n_37),
.B1(n_54),
.B2(n_56),
.Y(n_132)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx11_ASAP7_75t_SL g55 ( 
.A(n_16),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_17),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_116),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_17),
.A2(n_60),
.B1(n_61),
.B2(n_116),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_17),
.A2(n_54),
.B1(n_56),
.B2(n_116),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_22),
.B(n_43),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_24),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_30),
.Y(n_31)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_26),
.A2(n_35),
.B(n_120),
.C(n_121),
.Y(n_119)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_32),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_32),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_29),
.A2(n_32),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_29),
.A2(n_32),
.B1(n_106),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_29),
.A2(n_32),
.B1(n_115),
.B2(n_190),
.Y(n_189)
);

AO22x1_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_32),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_33),
.A2(n_66),
.B(n_68),
.C(n_69),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_66),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g270 ( 
.A1(n_33),
.A2(n_61),
.A3(n_70),
.B1(n_263),
.B2(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_34),
.B(n_120),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_82),
.B(n_336),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_75),
.C(n_77),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_44),
.A2(n_45),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_63),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_46),
.B(n_320),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_48),
.A2(n_79),
.B1(n_81),
.B2(n_170),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_52),
.A2(n_311),
.B1(n_313),
.B2(n_314),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_52),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_52),
.A2(n_63),
.B1(n_314),
.B2(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_58),
.B(n_62),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_58),
.B1(n_98),
.B2(n_101),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_53),
.A2(n_58),
.B1(n_101),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_53),
.A2(n_58),
.B1(n_62),
.B2(n_143),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_53),
.A2(n_58),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_53),
.A2(n_58),
.B1(n_221),
.B2(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_53),
.B(n_120),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_53),
.A2(n_58),
.B1(n_188),
.B2(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_54),
.B(n_57),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_54),
.B(n_252),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_61),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_60),
.B(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_63),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_74),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_64),
.A2(n_74),
.B1(n_111),
.B2(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_64),
.A2(n_74),
.B1(n_184),
.B2(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_64),
.A2(n_72),
.B1(n_74),
.B2(n_312),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_69),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_65),
.A2(n_69),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_65),
.A2(n_69),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_65),
.A2(n_69),
.B1(n_128),
.B2(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_65),
.A2(n_69),
.B1(n_196),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_70),
.Y(n_272)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_75),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_81),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_79),
.A2(n_81),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_329),
.B(n_335),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_305),
.A3(n_324),
.B1(n_327),
.B2(n_328),
.C(n_340),
.Y(n_83)
);

AOI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_154),
.A3(n_176),
.B1(n_299),
.B2(n_304),
.C(n_341),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_86),
.A2(n_300),
.B(n_303),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_135),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_87),
.B(n_135),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_112),
.C(n_130),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_88),
.B(n_130),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_102),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_103),
.C(n_108),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_97),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_90),
.B(n_97),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_96),
.B1(n_125),
.B2(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_91),
.A2(n_125),
.B(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_91),
.A2(n_95),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_91),
.A2(n_95),
.B1(n_240),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_91),
.A2(n_235),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_94),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_92),
.A2(n_123),
.B1(n_126),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_92),
.A2(n_126),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_95),
.B(n_120),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_99),
.A2(n_141),
.B1(n_144),
.B2(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_112),
.B(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_127),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_113),
.B(n_127),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_118),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_119),
.B(n_122),
.Y(n_191)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_SL g274 ( 
.A(n_126),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_153),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_147),
.C(n_153),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_145),
.B2(n_146),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_146),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_141),
.A2(n_144),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_146),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_145),
.A2(n_168),
.B(n_171),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_147),
.Y(n_338)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_150),
.CI(n_152),
.CON(n_147),
.SN(n_147)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_150),
.C(n_152),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_155),
.B(n_156),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_174),
.B2(n_175),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_159),
.B(n_165),
.C(n_175),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_163),
.B(n_164),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_163),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_162),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_164),
.B(n_307),
.C(n_316),
.Y(n_306)
);

FAx1_ASAP7_75t_L g326 ( 
.A(n_164),
.B(n_307),
.CI(n_316),
.CON(n_326),
.SN(n_326)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_174),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_206),
.C(n_211),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_200),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_178),
.B(n_200),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_191),
.C(n_192),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_179),
.B(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_186),
.C(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_297),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_191),
.Y(n_297)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_194),
.B(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_197),
.B(n_199),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_198),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_203),
.C(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_207),
.A2(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_208),
.B(n_209),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_293),
.B(n_298),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_279),
.B(n_292),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_256),
.B(n_278),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_236),
.B(n_255),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_226),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_216),
.B(n_226),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_217),
.A2(n_218),
.B1(n_222),
.B2(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_231),
.C(n_233),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_232),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_234),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_243),
.B(n_254),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_242),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_248),
.B(n_253),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_247),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_258),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_269),
.B1(n_276),
.B2(n_277),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_264),
.B1(n_267),
.B2(n_268),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_268),
.C(n_277),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_269),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_273),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_281),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_288),
.C(n_290),
.Y(n_294)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_288),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_317),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_317),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_315),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_309),
.B1(n_319),
.B2(n_322),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_311),
.C(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_322),
.C(n_323),
.Y(n_330)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_311),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_326),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule