module fake_jpeg_8104_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_48),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_33),
.B1(n_26),
.B2(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_54),
.B1(n_28),
.B2(n_34),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_52),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_33),
.B1(n_26),
.B2(n_28),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_69),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_26),
.B1(n_28),
.B2(n_47),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_65),
.A2(n_18),
.B1(n_34),
.B2(n_20),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_43),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_51),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_46),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_42),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_25),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_77),
.A2(n_81),
.B(n_100),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_79),
.B(n_82),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_109),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_86),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_59),
.B1(n_37),
.B2(n_8),
.Y(n_129)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_89),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_40),
.C(n_70),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_2),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_101),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_99),
.B1(n_53),
.B2(n_59),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_22),
.B(n_19),
.C(n_30),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_20),
.B(n_21),
.C(n_31),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_23),
.B1(n_31),
.B2(n_34),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_23),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_19),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_69),
.B(n_30),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_22),
.C(n_24),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_11),
.B1(n_10),
.B2(n_8),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_112),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_21),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_138),
.B(n_100),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_121),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_46),
.B1(n_43),
.B2(n_58),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_123),
.A2(n_130),
.B1(n_76),
.B2(n_108),
.Y(n_168)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_86),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_131),
.B1(n_135),
.B2(n_102),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_129),
.A2(n_139),
.B(n_143),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_75),
.A2(n_37),
.B1(n_15),
.B2(n_14),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_75),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_136),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_79),
.C(n_82),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_138)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_144),
.A2(n_152),
.B1(n_160),
.B2(n_176),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_SL g199 ( 
.A(n_145),
.B(n_157),
.C(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

AO21x2_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_99),
.B(n_100),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_155),
.B1(n_158),
.B2(n_166),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_78),
.Y(n_201)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_159),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_93),
.B(n_81),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_162),
.B(n_172),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_140),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_101),
.C(n_89),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_174),
.C(n_90),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_154),
.A2(n_115),
.B1(n_85),
.B2(n_5),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_112),
.B1(n_88),
.B2(n_83),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_117),
.B(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_77),
.B(n_81),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_135),
.B1(n_142),
.B2(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_77),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_163),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_98),
.B(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_110),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_170),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_119),
.B1(n_116),
.B2(n_130),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_133),
.B1(n_120),
.B2(n_125),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_137),
.B(n_91),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_121),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_90),
.Y(n_171)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_117),
.A2(n_91),
.B(n_95),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_175),
.B(n_177),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_125),
.C(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_169),
.B(n_161),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_147),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_179),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_193),
.C(n_203),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_174),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_190),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_182),
.Y(n_227)
);

AO22x1_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_76),
.B1(n_139),
.B2(n_126),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_184),
.A2(n_199),
.B(n_183),
.C(n_196),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_122),
.B1(n_115),
.B2(n_126),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_200),
.B1(n_148),
.B2(n_154),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_111),
.B(n_94),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_148),
.B(n_147),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_165),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_192),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_78),
.C(n_132),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_173),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_148),
.A2(n_164),
.B1(n_167),
.B2(n_158),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_7),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_149),
.B(n_78),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_145),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_187),
.C(n_193),
.Y(n_236)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_225)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_211),
.B(n_231),
.Y(n_256)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_194),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_218),
.B1(n_222),
.B2(n_202),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_200),
.A2(n_170),
.B1(n_85),
.B2(n_104),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_186),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_223),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_225),
.A2(n_238),
.B1(n_184),
.B2(n_188),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_235),
.C(n_236),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_237),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_199),
.B(n_204),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_179),
.A2(n_206),
.B1(n_197),
.B2(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_185),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_233),
.B(n_230),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_178),
.B(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_228),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_243),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_212),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_245),
.B(n_261),
.Y(n_269)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_214),
.A2(n_194),
.B1(n_180),
.B2(n_201),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_203),
.C(n_182),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_258),
.C(n_259),
.Y(n_268)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_213),
.A2(n_224),
.B1(n_238),
.B2(n_222),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_260),
.B1(n_239),
.B2(n_250),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_236),
.C(n_235),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_274),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_257),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_238),
.B1(n_215),
.B2(n_220),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_264),
.B(n_269),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_221),
.Y(n_267)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_238),
.B(n_226),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_278),
.B(n_243),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_238),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_273),
.Y(n_290)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_270),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_225),
.C(n_258),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_277),
.C(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_252),
.C(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_256),
.C(n_259),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_282),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_279),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_278),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_288),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_263),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_285),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_272),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_268),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_296),
.C(n_293),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_277),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_299),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_268),
.B(n_271),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_305),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_273),
.B1(n_292),
.B2(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_309),
.C(n_290),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_281),
.B1(n_294),
.B2(n_290),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_301),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_295),
.C(n_296),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_313),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_309),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_317),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_304),
.C(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_318),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_301),
.A2(n_306),
.B(n_309),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_307),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_319),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_314),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_313),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_326),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_322),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_320),
.B(n_328),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_323),
.Y(n_334)
);


endmodule