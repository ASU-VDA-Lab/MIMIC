module fake_jpeg_2443_n_221 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_221);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx8_ASAP7_75t_SL g74 ( 
.A(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_66),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_61),
.Y(n_100)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx4f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_66),
.Y(n_85)
);

CKINVDCx12_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_78),
.B1(n_70),
.B2(n_73),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_78),
.B1(n_70),
.B2(n_67),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_67),
.B1(n_57),
.B2(n_60),
.Y(n_106)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_71),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_68),
.B1(n_73),
.B2(n_62),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_69),
.B1(n_87),
.B2(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_107),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_57),
.B1(n_60),
.B2(n_72),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_77),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_56),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_114),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_77),
.Y(n_114)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_91),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_110),
.A2(n_87),
.B1(n_69),
.B2(n_68),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_131),
.B1(n_133),
.B2(n_102),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_58),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_75),
.B(n_62),
.C(n_98),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_104),
.B(n_9),
.C(n_11),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_69),
.B1(n_63),
.B2(n_59),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_1),
.B(n_2),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_119),
.B(n_104),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_63),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_2),
.C(n_3),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_14),
.C(n_15),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_59),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_4),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_5),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_26),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_148),
.B1(n_153),
.B2(n_134),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_119),
.B1(n_7),
.B2(n_8),
.Y(n_148)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NAND4xp25_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.D(n_161),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_162),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_R g174 ( 
.A(n_156),
.B(n_33),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_6),
.B(n_12),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_16),
.B(n_19),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_35),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_28),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_163),
.Y(n_177)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_20),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_121),
.B1(n_131),
.B2(n_124),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_124),
.C(n_138),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_184),
.C(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_173),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_175),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_174),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_34),
.B1(n_50),
.B2(n_49),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_21),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_180),
.B(n_164),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_146),
.B(n_22),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_156),
.B1(n_24),
.B2(n_25),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_40),
.C(n_46),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_192),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_179),
.A2(n_154),
.B(n_176),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_189),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_157),
.C(n_152),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_190),
.C(n_194),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_149),
.C(n_159),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_179),
.A2(n_156),
.B(n_41),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_39),
.C(n_51),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

XNOR2x2_ASAP7_75t_SL g199 ( 
.A(n_196),
.B(n_156),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

BUFx12_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_177),
.C(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_44),
.C(n_27),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_208),
.C(n_211),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_200),
.A2(n_191),
.B(n_175),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_205),
.A2(n_165),
.B1(n_181),
.B2(n_25),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_210),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_165),
.B1(n_181),
.B2(n_23),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_198),
.C(n_203),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_208),
.C(n_206),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_209),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_218),
.A2(n_215),
.B(n_212),
.Y(n_219)
);

OAI211xp5_ASAP7_75t_SL g220 ( 
.A1(n_219),
.A2(n_202),
.B(n_199),
.C(n_43),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_23),
.C(n_24),
.Y(n_221)
);


endmodule