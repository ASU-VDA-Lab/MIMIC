module fake_netlist_5_1891_n_2079 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2079);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2079;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1360;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_69),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_87),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_47),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_62),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_63),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_43),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_126),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_38),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_122),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_103),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_64),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_82),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_76),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_44),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_5),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_71),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_64),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_68),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_21),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_23),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_152),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_50),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_53),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_190),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_44),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_139),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_137),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_130),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_140),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_5),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_41),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_86),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_46),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_85),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_183),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_63),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_79),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_112),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_192),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_69),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_22),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_21),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_179),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_120),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_162),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_127),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_123),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_22),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_134),
.Y(n_254)
);

CKINVDCx11_ASAP7_75t_R g255 ( 
.A(n_95),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_20),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_104),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_153),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_16),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_167),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_90),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_155),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_143),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_19),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_144),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_61),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_52),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_35),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_12),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_129),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_169),
.Y(n_272)
);

BUFx8_ASAP7_75t_SL g273 ( 
.A(n_180),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_182),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_146),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_111),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_48),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_131),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_41),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_191),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_6),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_105),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_133),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_175),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_57),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_39),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_26),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_150),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_51),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_84),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_3),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_37),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_93),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_62),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_24),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_59),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_141),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_66),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_38),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_128),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_142),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_26),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_138),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_8),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_24),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_14),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_94),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_28),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_28),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_184),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_17),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_76),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_193),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_101),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_23),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_47),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_74),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_92),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_174),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_185),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_55),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_33),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_115),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_6),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_80),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_27),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_49),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_37),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_78),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_1),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_35),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_156),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_65),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_54),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_8),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_187),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_70),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_73),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_32),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_97),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_45),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_74),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_186),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_7),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_11),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_13),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_100),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_2),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_109),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_65),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_91),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_61),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_45),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_3),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_147),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_49),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_42),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_34),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_16),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_55),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_114),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_1),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_36),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_118),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_30),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_164),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_33),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_145),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_20),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_11),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_18),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_99),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_57),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_42),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_75),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_10),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_171),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_165),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_71),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_18),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_31),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_151),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_113),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_9),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_89),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_36),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_177),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_58),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_39),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_200),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_302),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_273),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_245),
.B(n_0),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_195),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_195),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_255),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_302),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_197),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_201),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_380),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_302),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_302),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_233),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_302),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_302),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_236),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_274),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_283),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_319),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_286),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_203),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_205),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_302),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_385),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_286),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_234),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_206),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_209),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_211),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_318),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_302),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_224),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_302),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_227),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_271),
.B(n_0),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_314),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_208),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_208),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_285),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_229),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_231),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_232),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_243),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_249),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_301),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_198),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_285),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_330),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_196),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_313),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_250),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_199),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_330),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_337),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_247),
.B(n_2),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_301),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_271),
.B(n_4),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_247),
.B(n_4),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_301),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_194),
.B(n_7),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_384),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_254),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_337),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_200),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_194),
.B(n_9),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_257),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_260),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_233),
.B(n_188),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_202),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_261),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_202),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_196),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_262),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_266),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_272),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_301),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_213),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_278),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_216),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_280),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_271),
.B(n_10),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_282),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_284),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_237),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_293),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_297),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_217),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_213),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_300),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_221),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_361),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_303),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_307),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_310),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_218),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_320),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_218),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_222),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_222),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_400),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_406),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_440),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_440),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_398),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_454),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_391),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_454),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_442),
.B(n_394),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_391),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_459),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_459),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_458),
.Y(n_504)
);

AND2x6_ASAP7_75t_L g505 ( 
.A(n_458),
.B(n_313),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_399),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_420),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_411),
.B(n_361),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_412),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_417),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_403),
.B(n_237),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_458),
.B(n_313),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_458),
.B(n_313),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_440),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_418),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_461),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_440),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_481),
.B(n_365),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_416),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_467),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_400),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_407),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_436),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_419),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_R g525 ( 
.A(n_392),
.B(n_323),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_467),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_422),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_440),
.B(n_313),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_424),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_478),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_430),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_469),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_478),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_485),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_477),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_408),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_485),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_487),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_487),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_488),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_433),
.B(n_290),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_488),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_397),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_489),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_489),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_397),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_401),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_401),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_480),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_402),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_402),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_404),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_405),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_441),
.B(n_290),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_405),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_413),
.Y(n_558)
);

INVxp33_ASAP7_75t_SL g559 ( 
.A(n_396),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_426),
.B(n_332),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_474),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_413),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_452),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_421),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_409),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_456),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_457),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_421),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_460),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_511),
.B(n_395),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_508),
.B(n_464),
.Y(n_571)
);

INVx8_ASAP7_75t_L g572 ( 
.A(n_505),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_495),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_548),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_548),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_548),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_547),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_542),
.B(n_468),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_504),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_556),
.B(n_472),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_547),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_497),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_511),
.B(n_390),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_499),
.B(n_473),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_549),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_492),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_561),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_561),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_549),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_554),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_497),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_506),
.B(n_475),
.Y(n_592)
);

AND2x2_ASAP7_75t_SL g593 ( 
.A(n_490),
.B(n_325),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_492),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_504),
.Y(n_595)
);

NAND2x1p5_ASAP7_75t_L g596 ( 
.A(n_504),
.B(n_207),
.Y(n_596)
);

OAI21xp33_ASAP7_75t_L g597 ( 
.A1(n_518),
.A2(n_448),
.B(n_445),
.Y(n_597)
);

AO22x2_ASAP7_75t_L g598 ( 
.A1(n_519),
.A2(n_393),
.B1(n_415),
.B2(n_445),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_505),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_532),
.B(n_476),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_509),
.B(n_479),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_532),
.B(n_482),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_492),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_518),
.B(n_390),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_492),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_554),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_505),
.B(n_484),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_500),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_496),
.B(n_474),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_555),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_555),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_505),
.B(n_486),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_496),
.B(n_427),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_492),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_492),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_557),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_498),
.B(n_425),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_500),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_557),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_562),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_514),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_490),
.B(n_451),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_514),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_562),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_510),
.B(n_432),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_544),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_544),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_564),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_553),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_532),
.B(n_451),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_498),
.B(n_501),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_564),
.Y(n_632)
);

INVxp67_ASAP7_75t_SL g633 ( 
.A(n_551),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_568),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_505),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_568),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_553),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_501),
.B(n_427),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_523),
.A2(n_309),
.B1(n_317),
.B2(n_311),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_505),
.B(n_425),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_558),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_558),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_514),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_558),
.Y(n_644)
);

AND2x6_ASAP7_75t_L g645 ( 
.A(n_558),
.B(n_325),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_551),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_521),
.A2(n_228),
.B1(n_415),
.B2(n_348),
.Y(n_647)
);

INVx6_ASAP7_75t_L g648 ( 
.A(n_551),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_551),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_551),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_505),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_533),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_536),
.A2(n_326),
.B1(n_327),
.B2(n_324),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_502),
.B(n_428),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_551),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_552),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_521),
.B(n_410),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_552),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_512),
.B(n_447),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_550),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_515),
.Y(n_661)
);

NAND2x1_ASAP7_75t_L g662 ( 
.A(n_512),
.B(n_368),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_552),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_552),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_524),
.B(n_434),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_552),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_552),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_502),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_514),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_494),
.Y(n_670)
);

BUFx8_ASAP7_75t_SL g671 ( 
.A(n_491),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_494),
.Y(n_672)
);

NAND2x1p5_ASAP7_75t_L g673 ( 
.A(n_503),
.B(n_207),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_527),
.B(n_463),
.Y(n_674)
);

INVx8_ASAP7_75t_L g675 ( 
.A(n_512),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_494),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_493),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_507),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_514),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_512),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_512),
.B(n_447),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_503),
.B(n_471),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_529),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_512),
.A2(n_471),
.B1(n_455),
.B2(n_450),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_512),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_522),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_532),
.B(n_483),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_516),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_516),
.B(n_368),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_513),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_531),
.B(n_465),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_560),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_520),
.B(n_428),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_514),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_517),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_520),
.B(n_429),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_563),
.B(n_470),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_566),
.Y(n_698)
);

BUFx6f_ASAP7_75t_SL g699 ( 
.A(n_513),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_517),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_537),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_517),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_526),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_526),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_517),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_567),
.B(n_439),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_517),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_530),
.B(n_210),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_530),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_569),
.B(n_439),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_534),
.B(n_210),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_513),
.B(n_423),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_534),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_517),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_559),
.B(n_462),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_513),
.B(n_423),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_513),
.B(n_239),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_493),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_513),
.B(n_252),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_535),
.B(n_462),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_513),
.B(n_340),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_493),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_571),
.B(n_493),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_583),
.A2(n_414),
.B1(n_351),
.B2(n_355),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_578),
.B(n_212),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_597),
.A2(n_214),
.B1(n_315),
.B2(n_292),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_617),
.B(n_212),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_583),
.A2(n_347),
.B1(n_372),
.B2(n_377),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_631),
.B(n_535),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_617),
.B(n_215),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_617),
.B(n_215),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_597),
.A2(n_214),
.B1(n_270),
.B2(n_292),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_604),
.B(n_342),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_604),
.B(n_223),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_588),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_574),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_617),
.B(n_219),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_599),
.B(n_301),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_682),
.B(n_219),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_599),
.B(n_301),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_631),
.B(n_538),
.Y(n_741)
);

NAND2x1_ASAP7_75t_L g742 ( 
.A(n_599),
.B(n_528),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_668),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_574),
.Y(n_744)
);

INVx8_ASAP7_75t_L g745 ( 
.A(n_671),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_579),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_682),
.B(n_220),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_708),
.A2(n_711),
.B1(n_684),
.B2(n_645),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_720),
.A2(n_315),
.B1(n_270),
.B2(n_365),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_574),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_668),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_SL g752 ( 
.A(n_639),
.B(n_346),
.C(n_338),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_644),
.A2(n_446),
.B(n_435),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_682),
.B(n_220),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_682),
.B(n_230),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_575),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_570),
.B(n_225),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_577),
.B(n_230),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_570),
.B(n_226),
.Y(n_759)
);

CKINVDCx11_ASAP7_75t_R g760 ( 
.A(n_678),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_706),
.B(n_235),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_633),
.A2(n_446),
.B(n_435),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_688),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_577),
.B(n_238),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_581),
.B(n_585),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_596),
.A2(n_349),
.B1(n_382),
.B2(n_383),
.Y(n_766)
);

AND2x6_ASAP7_75t_SL g767 ( 
.A(n_715),
.B(n_244),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_710),
.B(n_525),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_599),
.B(n_301),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_581),
.B(n_238),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_585),
.B(n_241),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_703),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_584),
.B(n_240),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_703),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_651),
.B(n_301),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_575),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_580),
.B(n_246),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_575),
.Y(n_778)
);

NOR2x2_ASAP7_75t_L g779 ( 
.A(n_639),
.B(n_653),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_576),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_589),
.B(n_241),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_642),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_589),
.B(n_242),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_587),
.B(n_393),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_609),
.B(n_590),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_642),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_609),
.B(n_538),
.Y(n_787)
);

AND2x6_ASAP7_75t_SL g788 ( 
.A(n_625),
.B(n_244),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_593),
.A2(n_378),
.B1(n_387),
.B2(n_242),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_573),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_651),
.B(n_301),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_576),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_576),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_704),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_SL g795 ( 
.A(n_692),
.B(n_565),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_579),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_579),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_590),
.B(n_248),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_606),
.B(n_248),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_647),
.B(n_264),
.C(n_256),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_704),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_661),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_651),
.B(n_251),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_606),
.B(n_251),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_610),
.B(n_263),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_610),
.B(n_611),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_593),
.A2(n_364),
.B1(n_263),
.B2(n_275),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_572),
.Y(n_808)
);

AND2x6_ASAP7_75t_SL g809 ( 
.A(n_665),
.B(n_253),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_587),
.B(n_253),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_652),
.B(n_259),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_SL g812 ( 
.A(n_692),
.B(n_357),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_618),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_709),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_708),
.A2(n_345),
.B(n_277),
.C(n_279),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_720),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_652),
.B(n_539),
.Y(n_817)
);

INVx5_ASAP7_75t_L g818 ( 
.A(n_572),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_SL g819 ( 
.A(n_683),
.B(n_371),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_611),
.B(n_275),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_708),
.A2(n_345),
.B1(n_277),
.B2(n_279),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_616),
.B(n_276),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_708),
.A2(n_352),
.B1(n_291),
.B2(n_295),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_660),
.B(n_259),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_657),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_709),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_L g827 ( 
.A(n_630),
.B(n_267),
.C(n_265),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_616),
.B(n_276),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_618),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_651),
.B(n_288),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_595),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_713),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_618),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_619),
.B(n_288),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_713),
.Y(n_835)
);

NAND2x1p5_ASAP7_75t_L g836 ( 
.A(n_635),
.B(n_329),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_711),
.A2(n_381),
.B1(n_291),
.B2(n_295),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_619),
.B(n_329),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_626),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_620),
.B(n_268),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_620),
.B(n_336),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_613),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_613),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_660),
.B(n_539),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_635),
.B(n_336),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_R g846 ( 
.A(n_698),
.B(n_269),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_635),
.B(n_349),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_628),
.B(n_364),
.Y(n_848)
);

AND3x2_ASAP7_75t_SL g849 ( 
.A(n_598),
.B(n_384),
.C(n_312),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_635),
.B(n_366),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_677),
.A2(n_446),
.B(n_435),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_628),
.B(n_281),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_626),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_632),
.B(n_287),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_595),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_595),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_635),
.B(n_366),
.Y(n_857)
);

AO221x1_ASAP7_75t_L g858 ( 
.A1(n_598),
.A2(n_376),
.B1(n_331),
.B2(n_341),
.C(n_352),
.Y(n_858)
);

AO22x1_ASAP7_75t_L g859 ( 
.A1(n_711),
.A2(n_341),
.B1(n_331),
.B2(n_354),
.Y(n_859)
);

AND2x6_ASAP7_75t_SL g860 ( 
.A(n_674),
.B(n_322),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_632),
.B(n_289),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_638),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_635),
.B(n_382),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_638),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_654),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_634),
.B(n_383),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_711),
.B(n_540),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_657),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_680),
.B(n_593),
.Y(n_869)
);

AND2x6_ASAP7_75t_SL g870 ( 
.A(n_697),
.B(n_592),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_642),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_634),
.B(n_540),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_622),
.B(n_541),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_680),
.B(n_449),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_654),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_693),
.Y(n_876)
);

NAND2x1p5_ASAP7_75t_L g877 ( 
.A(n_680),
.B(n_541),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_636),
.B(n_543),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_SL g879 ( 
.A(n_653),
.B(n_359),
.C(n_294),
.Y(n_879)
);

CKINVDCx8_ASAP7_75t_R g880 ( 
.A(n_601),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_691),
.B(n_622),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_600),
.B(n_543),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_693),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_636),
.B(n_296),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_624),
.B(n_298),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_686),
.B(n_545),
.Y(n_886)
);

HB1xp67_ASAP7_75t_SL g887 ( 
.A(n_598),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_624),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_696),
.A2(n_381),
.B(n_376),
.C(n_322),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_696),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_624),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_644),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_685),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_641),
.B(n_545),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_888),
.B(n_680),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_893),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_796),
.B(n_602),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_748),
.A2(n_690),
.B(n_685),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_733),
.B(n_687),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_893),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_735),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_790),
.B(n_701),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_825),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_892),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_818),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_802),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_893),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_787),
.B(n_785),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_888),
.B(n_680),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_725),
.B(n_596),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_813),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_777),
.B(n_596),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_SL g913 ( 
.A(n_752),
.B(n_304),
.C(n_299),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_829),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_796),
.B(n_690),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_777),
.B(n_641),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_893),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_SL g918 ( 
.A1(n_812),
.A2(n_598),
.B1(n_699),
.B2(n_572),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_SL g919 ( 
.A(n_879),
.B(n_306),
.C(n_305),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_868),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_743),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_761),
.A2(n_612),
.B1(n_607),
.B2(n_719),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_797),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_817),
.Y(n_924)
);

AND2x6_ASAP7_75t_L g925 ( 
.A(n_797),
.B(n_640),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_R g926 ( 
.A(n_795),
.B(n_699),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_751),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_745),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_818),
.B(n_680),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_785),
.B(n_673),
.Y(n_930)
);

AND2x4_ASAP7_75t_SL g931 ( 
.A(n_844),
.B(n_258),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_733),
.B(n_673),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_763),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_760),
.Y(n_934)
);

AO22x1_ASAP7_75t_L g935 ( 
.A1(n_761),
.A2(n_358),
.B1(n_308),
.B2(n_316),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_867),
.B(n_646),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_772),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_842),
.B(n_673),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_774),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_SL g940 ( 
.A(n_789),
.B(n_328),
.C(n_321),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_794),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_888),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_801),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_SL g944 ( 
.A(n_749),
.B(n_334),
.C(n_333),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_867),
.B(n_646),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_855),
.Y(n_946)
);

XNOR2xp5_ASAP7_75t_L g947 ( 
.A(n_887),
.B(n_717),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_R g948 ( 
.A(n_880),
.B(n_699),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_745),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_855),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_856),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_843),
.B(n_582),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_SL g953 ( 
.A(n_819),
.B(n_258),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_814),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_833),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_SL g956 ( 
.A(n_749),
.B(n_339),
.C(n_335),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_826),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_R g958 ( 
.A(n_745),
.B(n_572),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_839),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_888),
.B(n_712),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_853),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_856),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_746),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_746),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_768),
.B(n_816),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_SL g966 ( 
.A(n_773),
.B(n_350),
.C(n_344),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_736),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_746),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_746),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_734),
.B(n_582),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_734),
.B(n_591),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_744),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_818),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_SL g974 ( 
.A(n_773),
.B(n_356),
.C(n_353),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_750),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_729),
.B(n_649),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_756),
.Y(n_977)
);

CKINVDCx12_ASAP7_75t_R g978 ( 
.A(n_810),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_831),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_832),
.B(n_835),
.Y(n_980)
);

INVx6_ASAP7_75t_L g981 ( 
.A(n_831),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_862),
.B(n_591),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_776),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_876),
.B(n_608),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_748),
.B(n_716),
.Y(n_985)
);

AO21x2_ASAP7_75t_L g986 ( 
.A1(n_803),
.A2(n_681),
.B(n_659),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_831),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_831),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_778),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_757),
.A2(n_721),
.B1(n_667),
.B2(n_666),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_891),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_729),
.B(n_608),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_741),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_864),
.B(n_626),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_780),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_810),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_792),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_741),
.B(n_649),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_793),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_765),
.B(n_656),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_894),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_869),
.A2(n_662),
.B(n_637),
.C(n_629),
.Y(n_1002)
);

NAND2xp33_ASAP7_75t_SL g1003 ( 
.A(n_726),
.B(n_662),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_865),
.B(n_875),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_883),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_890),
.Y(n_1006)
);

XNOR2xp5_ASAP7_75t_L g1007 ( 
.A(n_784),
.B(n_77),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_810),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_806),
.B(n_656),
.Y(n_1009)
);

BUFx8_ASAP7_75t_L g1010 ( 
.A(n_873),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_757),
.B(n_664),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_818),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_759),
.B(n_664),
.Y(n_1013)
);

BUFx4f_ASAP7_75t_L g1014 ( 
.A(n_877),
.Y(n_1014)
);

INVx6_ASAP7_75t_L g1015 ( 
.A(n_886),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_869),
.B(n_650),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_872),
.Y(n_1017)
);

OR2x4_ASAP7_75t_L g1018 ( 
.A(n_759),
.B(n_354),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_878),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_SL g1020 ( 
.A(n_889),
.B(n_360),
.C(n_362),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_885),
.B(n_666),
.Y(n_1021)
);

AND2x2_ASAP7_75t_SL g1022 ( 
.A(n_807),
.B(n_726),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_758),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_732),
.B(n_627),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_885),
.B(n_667),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_SL g1026 ( 
.A(n_889),
.B(n_367),
.C(n_363),
.Y(n_1026)
);

NOR3xp33_ASAP7_75t_SL g1027 ( 
.A(n_815),
.B(n_375),
.C(n_389),
.Y(n_1027)
);

AND2x2_ASAP7_75t_SL g1028 ( 
.A(n_732),
.B(n_370),
.Y(n_1028)
);

NAND2x1p5_ASAP7_75t_L g1029 ( 
.A(n_808),
.B(n_722),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_742),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_SL g1031 ( 
.A(n_815),
.B(n_374),
.C(n_388),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_SL g1032 ( 
.A(n_840),
.B(n_386),
.C(n_379),
.Y(n_1032)
);

INVx5_ASAP7_75t_L g1033 ( 
.A(n_808),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_764),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_SL g1035 ( 
.A(n_840),
.B(n_369),
.C(n_852),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_811),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_770),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_882),
.B(n_650),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_877),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_771),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_781),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_852),
.B(n_655),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_727),
.A2(n_689),
.B1(n_645),
.B2(n_629),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_782),
.B(n_786),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_811),
.B(n_627),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_871),
.B(n_655),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_854),
.B(n_658),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_783),
.Y(n_1048)
);

NOR2x1_ASAP7_75t_L g1049 ( 
.A(n_811),
.B(n_722),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_SL g1050 ( 
.A(n_854),
.B(n_370),
.C(n_373),
.Y(n_1050)
);

BUFx2_ASAP7_75t_SL g1051 ( 
.A(n_845),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_SL g1052 ( 
.A(n_861),
.B(n_373),
.C(n_453),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_824),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_R g1054 ( 
.A(n_870),
.B(n_572),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_861),
.B(n_658),
.Y(n_1055)
);

NAND2xp33_ASAP7_75t_SL g1056 ( 
.A(n_846),
.B(n_663),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_824),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_798),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_SL g1059 ( 
.A(n_884),
.B(n_437),
.C(n_453),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_724),
.B(n_546),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_753),
.A2(n_675),
.B(n_663),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_730),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_824),
.B(n_204),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_884),
.B(n_722),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_731),
.B(n_722),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_737),
.B(n_627),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_739),
.B(n_629),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_836),
.Y(n_1068)
);

INVx4_ASAP7_75t_L g1069 ( 
.A(n_836),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_799),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_881),
.B(n_637),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_874),
.Y(n_1072)
);

INVx5_ASAP7_75t_L g1073 ( 
.A(n_767),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_874),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_723),
.B(n_675),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_747),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_804),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_754),
.B(n_637),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_755),
.A2(n_830),
.B1(n_803),
.B2(n_827),
.Y(n_1079)
);

INVx3_ASAP7_75t_SL g1080 ( 
.A(n_779),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_846),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_788),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_809),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_SL g1084 ( 
.A(n_849),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_805),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_820),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_860),
.Y(n_1087)
);

AO21x2_ASAP7_75t_L g1088 ( 
.A1(n_912),
.A2(n_830),
.B(n_828),
.Y(n_1088)
);

BUFx2_ASAP7_75t_SL g1089 ( 
.A(n_906),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1075),
.A2(n_740),
.B(n_775),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1075),
.A2(n_740),
.B(n_775),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_994),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_899),
.B(n_1015),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1019),
.B(n_728),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_994),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1016),
.A2(n_738),
.B(n_769),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_908),
.B(n_800),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_921),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_967),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_899),
.A2(n_858),
.B1(n_822),
.B2(n_834),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1022),
.A2(n_837),
.B(n_823),
.C(n_821),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_908),
.B(n_821),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_927),
.Y(n_1103)
);

NAND2x1_ASAP7_75t_L g1104 ( 
.A(n_900),
.B(n_648),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1017),
.B(n_932),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1016),
.A2(n_769),
.B(n_791),
.Y(n_1106)
);

NAND3x1_ASAP7_75t_L g1107 ( 
.A(n_1049),
.B(n_849),
.C(n_1063),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_1015),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_930),
.A2(n_766),
.A3(n_841),
.B(n_848),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_898),
.A2(n_791),
.B(n_851),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_906),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_967),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1015),
.B(n_823),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_933),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_964),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1061),
.A2(n_1002),
.B(n_1029),
.Y(n_1116)
);

O2A1O1Ixp5_ASAP7_75t_SL g1117 ( 
.A1(n_960),
.A2(n_866),
.B(n_838),
.C(n_845),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_964),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1029),
.A2(n_762),
.B(n_714),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_903),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_901),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_972),
.Y(n_1122)
);

NOR2x1_ASAP7_75t_SL g1123 ( 
.A(n_1033),
.B(n_847),
.Y(n_1123)
);

AO31x2_ASAP7_75t_L g1124 ( 
.A1(n_1011),
.A2(n_676),
.A3(n_670),
.B(n_672),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_932),
.B(n_837),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1017),
.B(n_859),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_960),
.A2(n_705),
.B(n_714),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1022),
.A2(n_863),
.B1(n_857),
.B2(n_850),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_924),
.B(n_1023),
.Y(n_1129)
);

BUFx4f_ASAP7_75t_L g1130 ( 
.A(n_920),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_972),
.Y(n_1131)
);

OA21x2_ASAP7_75t_L g1132 ( 
.A1(n_1042),
.A2(n_672),
.B(n_670),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1028),
.A2(n_546),
.B(n_857),
.C(n_850),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_985),
.A2(n_714),
.B(n_705),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_964),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1033),
.A2(n_675),
.B(n_586),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1028),
.A2(n_863),
.B(n_847),
.C(n_444),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_924),
.B(n_1034),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_985),
.A2(n_705),
.B(n_679),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_910),
.A2(n_676),
.B(n_645),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_922),
.A2(n_645),
.B(n_718),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_975),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_993),
.B(n_679),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1040),
.B(n_694),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_SL g1145 ( 
.A1(n_1062),
.A2(n_702),
.B(n_694),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1041),
.B(n_702),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1066),
.A2(n_594),
.B(n_707),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_1057),
.Y(n_1148)
);

O2A1O1Ixp5_ASAP7_75t_L g1149 ( 
.A1(n_970),
.A2(n_603),
.B(n_707),
.C(n_695),
.Y(n_1149)
);

INVx6_ASAP7_75t_SL g1150 ( 
.A(n_897),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1065),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1010),
.Y(n_1152)
);

NOR2xp67_ASAP7_75t_L g1153 ( 
.A(n_965),
.B(n_81),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_923),
.A2(n_594),
.B(n_707),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1048),
.B(n_718),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1077),
.A2(n_429),
.B(n_437),
.C(n_438),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_923),
.A2(n_621),
.B(n_707),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1079),
.A2(n_675),
.B1(n_648),
.B2(n_718),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1085),
.B(n_594),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_931),
.B(n_1004),
.Y(n_1160)
);

AO21x2_ASAP7_75t_L g1161 ( 
.A1(n_1013),
.A2(n_1025),
.B(n_1021),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_931),
.B(n_384),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_976),
.B(n_594),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1086),
.B(n_603),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1018),
.B(n_603),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_981),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1086),
.B(n_603),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_923),
.A2(n_605),
.B(n_695),
.Y(n_1168)
);

OAI22x1_ASAP7_75t_L g1169 ( 
.A1(n_1080),
.A2(n_204),
.B1(n_312),
.B2(n_444),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_993),
.B(n_605),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_993),
.B(n_605),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1080),
.B(n_438),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_975),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_902),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_946),
.A2(n_621),
.B(n_695),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_946),
.A2(n_621),
.B(n_695),
.Y(n_1176)
);

AOI221xp5_ASAP7_75t_L g1177 ( 
.A1(n_935),
.A2(n_443),
.B1(n_204),
.B2(n_312),
.C(n_384),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1005),
.A2(n_443),
.B(n_466),
.C(n_449),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1004),
.B(n_258),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1001),
.B(n_605),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1081),
.B(n_1036),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1033),
.A2(n_700),
.B(n_586),
.Y(n_1182)
);

INVxp67_ASAP7_75t_SL g1183 ( 
.A(n_964),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1033),
.A2(n_973),
.B(n_905),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_928),
.B(n_648),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1005),
.B(n_343),
.Y(n_1186)
);

NAND2x1p5_ASAP7_75t_L g1187 ( 
.A(n_969),
.B(n_614),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_916),
.A2(n_645),
.B(n_621),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1001),
.B(n_614),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1024),
.A2(n_645),
.B(n_614),
.Y(n_1190)
);

BUFx2_ASAP7_75t_R g1191 ( 
.A(n_928),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_976),
.B(n_614),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1010),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1006),
.B(n_343),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1006),
.B(n_343),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1047),
.A2(n_449),
.A3(n_466),
.B(n_689),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1037),
.B(n_645),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1062),
.A2(n_648),
.B1(n_586),
.B2(n_669),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1060),
.B(n_12),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_900),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_947),
.B(n_689),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_949),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_946),
.A2(n_466),
.B(n_689),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_900),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1037),
.B(n_689),
.Y(n_1205)
);

NOR2x1_ASAP7_75t_SL g1206 ( 
.A(n_900),
.B(n_586),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1058),
.B(n_689),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1058),
.B(n_689),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_949),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_905),
.A2(n_700),
.B(n_669),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_950),
.A2(n_700),
.B(n_669),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_996),
.B(n_1008),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1055),
.A2(n_13),
.A3(n_14),
.B(n_15),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1044),
.A2(n_669),
.B1(n_643),
.B2(n_623),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_915),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1070),
.B(n_971),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_937),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_902),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1070),
.B(n_700),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1010),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1064),
.A2(n_15),
.A3(n_17),
.B(n_19),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_977),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1072),
.B(n_700),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_907),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_950),
.A2(n_669),
.B(n_643),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_980),
.B(n_643),
.Y(n_1226)
);

O2A1O1Ixp5_ASAP7_75t_L g1227 ( 
.A1(n_1056),
.A2(n_1003),
.B(n_1071),
.C(n_1009),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_939),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1044),
.B(n_643),
.Y(n_1229)
);

OR2x6_ASAP7_75t_L g1230 ( 
.A(n_897),
.B(n_643),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1071),
.A2(n_25),
.A3(n_27),
.B(n_29),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_950),
.A2(n_623),
.B(n_615),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_897),
.B(n_25),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1000),
.A2(n_623),
.B(n_615),
.Y(n_1234)
);

NAND3x1_ASAP7_75t_L g1235 ( 
.A(n_1084),
.B(n_29),
.C(n_30),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1044),
.B(n_623),
.Y(n_1236)
);

NOR2x1_ASAP7_75t_SL g1237 ( 
.A(n_907),
.B(n_623),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1045),
.B(n_31),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_951),
.A2(n_615),
.B(n_586),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1072),
.B(n_615),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_951),
.A2(n_615),
.B(n_106),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1072),
.B(n_102),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_941),
.B(n_528),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_943),
.A2(n_32),
.A3(n_34),
.B(n_40),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_954),
.A2(n_40),
.A3(n_43),
.B(n_46),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_905),
.A2(n_528),
.B(n_116),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_973),
.A2(n_528),
.B(n_108),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_934),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1024),
.A2(n_528),
.B(n_117),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_957),
.B(n_528),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_952),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1120),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1147),
.A2(n_962),
.B(n_951),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1092),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1098),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1105),
.B(n_1076),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1199),
.A2(n_953),
.B1(n_1018),
.B2(n_1073),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1147),
.A2(n_962),
.B(n_990),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1163),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1116),
.A2(n_962),
.B(n_896),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1120),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1174),
.A2(n_1073),
.B1(n_1082),
.B2(n_1053),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1227),
.A2(n_1059),
.B(n_1052),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1193),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1094),
.A2(n_940),
.B(n_1035),
.C(n_1050),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1200),
.Y(n_1266)
);

NOR2x1_ASAP7_75t_SL g1267 ( 
.A(n_1088),
.B(n_973),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1089),
.B(n_969),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1211),
.A2(n_896),
.B(n_959),
.Y(n_1269)
);

BUFx8_ASAP7_75t_L g1270 ( 
.A(n_1181),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1099),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1097),
.A2(n_918),
.B1(n_1084),
.B2(n_1076),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1103),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1125),
.A2(n_1003),
.B(n_992),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1234),
.A2(n_1038),
.B(n_904),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1216),
.A2(n_1012),
.B(n_929),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1121),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1211),
.A2(n_961),
.B(n_959),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1163),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1111),
.Y(n_1280)
);

AOI22x1_ASAP7_75t_L g1281 ( 
.A1(n_1249),
.A2(n_938),
.B1(n_977),
.B2(n_983),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1114),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1172),
.Y(n_1283)
);

CKINVDCx9p33_ASAP7_75t_R g1284 ( 
.A(n_1093),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1102),
.B(n_938),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1225),
.A2(n_914),
.B(n_911),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1130),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1149),
.A2(n_955),
.B(n_914),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1111),
.B(n_976),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1225),
.A2(n_955),
.B(n_961),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1125),
.A2(n_952),
.B(n_982),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1092),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1151),
.A2(n_999),
.B(n_997),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1095),
.B(n_982),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1161),
.A2(n_986),
.B(n_1027),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1200),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1093),
.A2(n_1084),
.B1(n_1053),
.B2(n_998),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1112),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1101),
.A2(n_968),
.B1(n_1014),
.B2(n_981),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1112),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1122),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1122),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1131),
.Y(n_1303)
);

O2A1O1Ixp5_ASAP7_75t_L g1304 ( 
.A1(n_1110),
.A2(n_1056),
.B(n_963),
.C(n_1014),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1232),
.A2(n_1239),
.B(n_1127),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1251),
.B(n_1045),
.Y(n_1306)
);

BUFx4f_ASAP7_75t_L g1307 ( 
.A(n_1200),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1232),
.A2(n_983),
.B(n_999),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1100),
.A2(n_984),
.B(n_1043),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1239),
.A2(n_989),
.B(n_997),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1131),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1177),
.B(n_913),
.C(n_966),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1161),
.A2(n_986),
.B(n_1031),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1129),
.B(n_1083),
.Y(n_1314)
);

OA21x2_ASAP7_75t_L g1315 ( 
.A1(n_1151),
.A2(n_989),
.B(n_995),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1127),
.A2(n_995),
.B(n_963),
.Y(n_1316)
);

INVx3_ASAP7_75t_SL g1317 ( 
.A(n_1218),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1126),
.B(n_991),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_SL g1319 ( 
.A1(n_1145),
.A2(n_942),
.B(n_1069),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1142),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1212),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1165),
.B(n_974),
.C(n_1032),
.Y(n_1322)
);

AO21x2_ASAP7_75t_L g1323 ( 
.A1(n_1141),
.A2(n_1020),
.B(n_1026),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1241),
.A2(n_1046),
.B(n_895),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1101),
.A2(n_998),
.B(n_1046),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1154),
.A2(n_1168),
.B(n_1157),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1138),
.A2(n_1014),
.B1(n_981),
.B2(n_942),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1154),
.A2(n_963),
.B(n_1068),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1160),
.B(n_1082),
.Y(n_1329)
);

AOI221xp5_ASAP7_75t_L g1330 ( 
.A1(n_1169),
.A2(n_944),
.B1(n_956),
.B2(n_1082),
.C(n_1087),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1157),
.A2(n_1068),
.B(n_909),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1148),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1241),
.A2(n_1046),
.B(n_909),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1191),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1117),
.A2(n_998),
.B(n_936),
.Y(n_1335)
);

BUFx12f_ASAP7_75t_L g1336 ( 
.A(n_1152),
.Y(n_1336)
);

NOR2x1_ASAP7_75t_SL g1337 ( 
.A(n_1088),
.B(n_1012),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1217),
.Y(n_1338)
);

BUFx2_ASAP7_75t_SL g1339 ( 
.A(n_1218),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1215),
.A2(n_1113),
.B1(n_1228),
.B2(n_1230),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1220),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1215),
.A2(n_915),
.B1(n_907),
.B2(n_917),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1109),
.B(n_936),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1201),
.A2(n_945),
.B1(n_936),
.B2(n_1007),
.Y(n_1344)
);

OR2x6_ASAP7_75t_L g1345 ( 
.A(n_1230),
.B(n_1185),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1142),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1132),
.A2(n_1038),
.B(n_895),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1150),
.A2(n_1073),
.B1(n_1087),
.B2(n_1074),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1163),
.B(n_945),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1168),
.A2(n_1068),
.B(n_925),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1108),
.Y(n_1351)
);

OR2x6_ASAP7_75t_L g1352 ( 
.A(n_1230),
.B(n_979),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1175),
.A2(n_925),
.B(n_1051),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1192),
.B(n_945),
.Y(n_1354)
);

AO21x2_ASAP7_75t_L g1355 ( 
.A1(n_1140),
.A2(n_1188),
.B(n_1190),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1175),
.A2(n_925),
.B(n_1069),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1150),
.A2(n_1073),
.B1(n_1074),
.B2(n_1072),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1238),
.B(n_919),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1233),
.B(n_1074),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1128),
.A2(n_925),
.B(n_1038),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1173),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1176),
.A2(n_925),
.B(n_1069),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1248),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1173),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1150),
.A2(n_1054),
.B1(n_926),
.B2(n_1074),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1222),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1183),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1176),
.A2(n_925),
.B(n_1030),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1222),
.Y(n_1369)
);

OAI222xp33_ASAP7_75t_L g1370 ( 
.A1(n_1186),
.A2(n_1073),
.B1(n_1039),
.B2(n_978),
.C1(n_915),
.C2(n_1054),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1139),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1180),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1155),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1139),
.A2(n_1030),
.B(n_907),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1144),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1192),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1134),
.A2(n_1030),
.B(n_917),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1146),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1192),
.Y(n_1379)
);

AND2x6_ASAP7_75t_L g1380 ( 
.A(n_1200),
.B(n_917),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1108),
.B(n_988),
.Y(n_1381)
);

CKINVDCx8_ASAP7_75t_R g1382 ( 
.A(n_1204),
.Y(n_1382)
);

NOR2x1_ASAP7_75t_SL g1383 ( 
.A(n_1242),
.B(n_917),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1204),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1134),
.A2(n_1030),
.B(n_1039),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1165),
.A2(n_948),
.B1(n_988),
.B2(n_987),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1118),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1136),
.A2(n_1039),
.B(n_988),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1179),
.B(n_988),
.C(n_987),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1156),
.A2(n_948),
.B(n_958),
.C(n_52),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1229),
.A2(n_987),
.B1(n_979),
.B2(n_969),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1189),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1090),
.A2(n_987),
.B(n_979),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1090),
.A2(n_1091),
.B(n_1119),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1223),
.A2(n_958),
.B(n_969),
.Y(n_1395)
);

A2O1A1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1133),
.A2(n_979),
.B(n_51),
.C(n_53),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1194),
.A2(n_528),
.B1(n_54),
.B2(n_56),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1159),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1223),
.A2(n_121),
.B(n_173),
.Y(n_1399)
);

INVx5_ASAP7_75t_L g1400 ( 
.A(n_1204),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1220),
.A2(n_50),
.B1(n_56),
.B2(n_58),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1178),
.A2(n_59),
.B(n_60),
.Y(n_1402)
);

CKINVDCx16_ASAP7_75t_R g1403 ( 
.A(n_1202),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1124),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1162),
.B(n_60),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1091),
.A2(n_125),
.B(n_172),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1164),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1204),
.Y(n_1408)
);

INVx2_ASAP7_75t_SL g1409 ( 
.A(n_1224),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1124),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1195),
.B(n_66),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1202),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1209),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1182),
.A2(n_132),
.B(n_166),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1209),
.B(n_124),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1185),
.B(n_119),
.Y(n_1416)
);

AO31x2_ASAP7_75t_L g1417 ( 
.A1(n_1178),
.A2(n_67),
.A3(n_68),
.B(n_70),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1133),
.A2(n_67),
.B(n_72),
.C(n_73),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1124),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1255),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1273),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1401),
.A2(n_1242),
.B1(n_1153),
.B2(n_1235),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1412),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1363),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1321),
.B(n_1156),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1403),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1272),
.A2(n_1107),
.B1(n_1235),
.B2(n_1185),
.Y(n_1427)
);

NOR3xp33_ASAP7_75t_SL g1428 ( 
.A(n_1312),
.B(n_1137),
.C(n_1170),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1285),
.B(n_1107),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1277),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1339),
.Y(n_1431)
);

INVx6_ASAP7_75t_L g1432 ( 
.A(n_1268),
.Y(n_1432)
);

CKINVDCx8_ASAP7_75t_R g1433 ( 
.A(n_1339),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1265),
.A2(n_1137),
.B(n_1205),
.C(n_1207),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1405),
.A2(n_1123),
.B1(n_1231),
.B2(n_1206),
.Y(n_1435)
);

INVx8_ASAP7_75t_L g1436 ( 
.A(n_1380),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1285),
.B(n_1166),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1314),
.B(n_1166),
.Y(n_1438)
);

AOI21xp33_ASAP7_75t_L g1439 ( 
.A1(n_1322),
.A2(n_1226),
.B(n_1208),
.Y(n_1439)
);

OAI211xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1330),
.A2(n_1167),
.B(n_1143),
.C(n_1171),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1360),
.A2(n_1158),
.B(n_1214),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1389),
.A2(n_1197),
.B(n_1106),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1282),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1281),
.A2(n_1231),
.B1(n_1237),
.B2(n_1245),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1294),
.B(n_1256),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1341),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1281),
.A2(n_1274),
.B(n_1325),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1257),
.A2(n_1143),
.B1(n_1171),
.B2(n_1170),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1294),
.B(n_1236),
.Y(n_1449)
);

OR2x6_ASAP7_75t_L g1450 ( 
.A(n_1345),
.B(n_1184),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1349),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1411),
.A2(n_1358),
.B1(n_1397),
.B2(n_1309),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1338),
.Y(n_1453)
);

BUFx4f_ASAP7_75t_L g1454 ( 
.A(n_1317),
.Y(n_1454)
);

CKINVDCx6p67_ASAP7_75t_R g1455 ( 
.A(n_1317),
.Y(n_1455)
);

BUFx12f_ASAP7_75t_L g1456 ( 
.A(n_1270),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1358),
.A2(n_1240),
.B1(n_1243),
.B2(n_1250),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1412),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1382),
.Y(n_1459)
);

BUFx4f_ASAP7_75t_L g1460 ( 
.A(n_1283),
.Y(n_1460)
);

OAI221xp5_ASAP7_75t_L g1461 ( 
.A1(n_1418),
.A2(n_1240),
.B1(n_1246),
.B2(n_1247),
.C(n_1219),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1359),
.B(n_1231),
.Y(n_1462)
);

INVxp33_ASAP7_75t_SL g1463 ( 
.A(n_1287),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1261),
.Y(n_1464)
);

OAI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1318),
.A2(n_1118),
.B1(n_1135),
.B2(n_1224),
.Y(n_1465)
);

NAND2xp33_ASAP7_75t_R g1466 ( 
.A(n_1289),
.B(n_1115),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1345),
.B(n_1118),
.Y(n_1467)
);

OAI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1396),
.A2(n_1104),
.B1(n_1198),
.B2(n_1187),
.C(n_1115),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1318),
.A2(n_1096),
.B1(n_1106),
.B2(n_1135),
.Y(n_1469)
);

NOR3xp33_ASAP7_75t_SL g1470 ( 
.A(n_1370),
.B(n_1210),
.C(n_1231),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1349),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1263),
.A2(n_1256),
.B1(n_1323),
.B2(n_1291),
.Y(n_1472)
);

INVx4_ASAP7_75t_R g1473 ( 
.A(n_1413),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1254),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1375),
.B(n_1135),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1263),
.A2(n_1224),
.B1(n_1221),
.B2(n_1213),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1271),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1394),
.A2(n_1203),
.B(n_1187),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1359),
.B(n_1244),
.Y(n_1479)
);

OAI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1297),
.A2(n_1109),
.B1(n_1221),
.B2(n_1213),
.C(n_1244),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1301),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1344),
.A2(n_1109),
.B1(n_1196),
.B2(n_1124),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1365),
.A2(n_1109),
.B1(n_1196),
.B2(n_1221),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1378),
.B(n_1306),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1277),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1348),
.B(n_1196),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1304),
.A2(n_1196),
.B(n_1221),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1376),
.B(n_1213),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1292),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1376),
.B(n_1213),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1298),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1332),
.Y(n_1492)
);

AOI222xp33_ASAP7_75t_L g1493 ( 
.A1(n_1283),
.A2(n_72),
.B1(n_75),
.B2(n_1245),
.C1(n_1244),
.C2(n_98),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1298),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1373),
.B(n_1245),
.Y(n_1495)
);

INVx6_ASAP7_75t_L g1496 ( 
.A(n_1268),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1289),
.B(n_1244),
.Y(n_1497)
);

AOI21xp33_ASAP7_75t_L g1498 ( 
.A1(n_1323),
.A2(n_1245),
.B(n_96),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1289),
.B(n_83),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1394),
.A2(n_107),
.B(n_135),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1300),
.Y(n_1501)
);

AOI222xp33_ASAP7_75t_L g1502 ( 
.A1(n_1329),
.A2(n_149),
.B1(n_154),
.B2(n_157),
.C1(n_158),
.C2(n_160),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1270),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1407),
.B(n_181),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1263),
.A2(n_1323),
.B1(n_1402),
.B2(n_1398),
.Y(n_1505)
);

NAND4xp25_ASAP7_75t_L g1506 ( 
.A(n_1252),
.B(n_1280),
.C(n_1334),
.D(n_1386),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1402),
.A2(n_1340),
.B1(n_1416),
.B2(n_1343),
.Y(n_1507)
);

NAND2x1p5_ASAP7_75t_L g1508 ( 
.A(n_1400),
.B(n_1387),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1302),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1349),
.B(n_1354),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1354),
.B(n_1259),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1354),
.B(n_1252),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1259),
.B(n_1279),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1259),
.B(n_1279),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1279),
.B(n_1379),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1336),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1379),
.B(n_1351),
.Y(n_1517)
);

CKINVDCx12_ASAP7_75t_R g1518 ( 
.A(n_1268),
.Y(n_1518)
);

AOI221x1_ASAP7_75t_L g1519 ( 
.A1(n_1299),
.A2(n_1335),
.B1(n_1414),
.B2(n_1391),
.C(n_1410),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1379),
.B(n_1392),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1345),
.B(n_1352),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1402),
.A2(n_1416),
.B1(n_1343),
.B2(n_1262),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1320),
.Y(n_1523)
);

OAI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1345),
.A2(n_1372),
.B1(n_1268),
.B2(n_1352),
.Y(n_1524)
);

INVx4_ASAP7_75t_SL g1525 ( 
.A(n_1380),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1336),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1372),
.B(n_1346),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1416),
.A2(n_1270),
.B1(n_1355),
.B2(n_1264),
.Y(n_1528)
);

AO221x2_ASAP7_75t_L g1529 ( 
.A1(n_1357),
.A2(n_1284),
.B1(n_1327),
.B2(n_1417),
.C(n_1342),
.Y(n_1529)
);

CKINVDCx16_ASAP7_75t_R g1530 ( 
.A(n_1341),
.Y(n_1530)
);

NAND2xp33_ASAP7_75t_R g1531 ( 
.A(n_1415),
.B(n_1367),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1302),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1355),
.A2(n_1415),
.B1(n_1303),
.B2(n_1366),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1387),
.Y(n_1534)
);

O2A1O1Ixp5_ASAP7_75t_SL g1535 ( 
.A1(n_1303),
.A2(n_1311),
.B(n_1361),
.C(n_1366),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_SL g1536 ( 
.A(n_1390),
.B(n_1367),
.C(n_1276),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1352),
.A2(n_1382),
.B1(n_1361),
.B2(n_1311),
.Y(n_1537)
);

NAND3xp33_ASAP7_75t_L g1538 ( 
.A(n_1415),
.B(n_1381),
.C(n_1352),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1364),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1384),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1307),
.A2(n_1400),
.B1(n_1387),
.B2(n_1408),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1384),
.B(n_1408),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1400),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1383),
.A2(n_1355),
.B1(n_1399),
.B2(n_1406),
.Y(n_1544)
);

AOI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1369),
.A2(n_1313),
.B1(n_1295),
.B2(n_1419),
.C(n_1404),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1267),
.A2(n_1337),
.B(n_1353),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1369),
.B(n_1409),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1295),
.A2(n_1313),
.B1(n_1399),
.B2(n_1324),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1388),
.A2(n_1385),
.B(n_1337),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1307),
.B(n_1400),
.Y(n_1550)
);

NAND2xp33_ASAP7_75t_SL g1551 ( 
.A(n_1266),
.B(n_1296),
.Y(n_1551)
);

AO31x2_ASAP7_75t_L g1552 ( 
.A1(n_1371),
.A2(n_1267),
.A3(n_1383),
.B(n_1295),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1266),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1266),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1307),
.Y(n_1555)
);

AO31x2_ASAP7_75t_L g1556 ( 
.A1(n_1313),
.A2(n_1293),
.A3(n_1315),
.B(n_1347),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1409),
.A2(n_1275),
.B1(n_1347),
.B2(n_1417),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1399),
.A2(n_1288),
.B1(n_1293),
.B2(n_1315),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1406),
.A2(n_1380),
.B1(n_1395),
.B2(n_1333),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1266),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1380),
.A2(n_1395),
.B1(n_1324),
.B2(n_1333),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1266),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1417),
.B(n_1296),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1296),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1380),
.A2(n_1333),
.B1(n_1324),
.B2(n_1296),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1296),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1293),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_SL g1568 ( 
.A(n_1380),
.B(n_1319),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1417),
.B(n_1315),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1260),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1547),
.Y(n_1571)
);

OAI221xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1452),
.A2(n_1417),
.B1(n_1319),
.B2(n_1275),
.C(n_1258),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1452),
.A2(n_1288),
.B1(n_1258),
.B2(n_1260),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1422),
.A2(n_1288),
.B1(n_1253),
.B2(n_1350),
.C(n_1316),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1493),
.A2(n_1253),
.B1(n_1316),
.B2(n_1350),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1420),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1437),
.B(n_1393),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1542),
.B(n_1393),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1422),
.A2(n_1308),
.B1(n_1278),
.B2(n_1286),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1421),
.Y(n_1580)
);

CKINVDCx11_ASAP7_75t_R g1581 ( 
.A(n_1433),
.Y(n_1581)
);

AO31x2_ASAP7_75t_L g1582 ( 
.A1(n_1519),
.A2(n_1487),
.A3(n_1483),
.B(n_1447),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1429),
.B(n_1331),
.Y(n_1583)
);

OAI211xp5_ASAP7_75t_L g1584 ( 
.A1(n_1502),
.A2(n_1331),
.B(n_1356),
.C(n_1362),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1562),
.Y(n_1585)
);

AOI222xp33_ASAP7_75t_L g1586 ( 
.A1(n_1427),
.A2(n_1328),
.B1(n_1278),
.B2(n_1286),
.C1(n_1290),
.C2(n_1308),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1538),
.A2(n_1385),
.B1(n_1362),
.B2(n_1368),
.Y(n_1587)
);

AOI222xp33_ASAP7_75t_L g1588 ( 
.A1(n_1454),
.A2(n_1328),
.B1(n_1290),
.B2(n_1310),
.C1(n_1368),
.C2(n_1377),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1506),
.A2(n_1310),
.B1(n_1269),
.B2(n_1374),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1529),
.A2(n_1454),
.B1(n_1536),
.B2(n_1445),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1424),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1528),
.A2(n_1377),
.B1(n_1374),
.B2(n_1269),
.Y(n_1592)
);

AOI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1425),
.A2(n_1305),
.B(n_1326),
.Y(n_1593)
);

OAI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1438),
.A2(n_1326),
.B1(n_1428),
.B2(n_1448),
.C(n_1528),
.Y(n_1594)
);

CKINVDCx6p67_ASAP7_75t_R g1595 ( 
.A(n_1456),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1462),
.B(n_1479),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1529),
.A2(n_1455),
.B1(n_1451),
.B2(n_1471),
.Y(n_1597)
);

OAI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1531),
.A2(n_1484),
.B1(n_1521),
.B2(n_1466),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_SL g1599 ( 
.A(n_1555),
.B(n_1426),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1451),
.A2(n_1471),
.B1(n_1440),
.B2(n_1511),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1440),
.A2(n_1511),
.B1(n_1536),
.B2(n_1463),
.Y(n_1601)
);

OAI211xp5_ASAP7_75t_SL g1602 ( 
.A1(n_1492),
.A2(n_1464),
.B(n_1430),
.C(n_1428),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1521),
.B(n_1540),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1447),
.A2(n_1441),
.B1(n_1498),
.B2(n_1492),
.Y(n_1604)
);

AO222x2_ASAP7_75t_L g1605 ( 
.A1(n_1530),
.A2(n_1497),
.B1(n_1513),
.B2(n_1446),
.C1(n_1563),
.C2(n_1499),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1431),
.A2(n_1503),
.B1(n_1460),
.B2(n_1510),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1512),
.B(n_1517),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1448),
.A2(n_1522),
.B1(n_1507),
.B2(n_1533),
.Y(n_1608)
);

OAI211xp5_ASAP7_75t_L g1609 ( 
.A1(n_1435),
.A2(n_1480),
.B(n_1470),
.C(n_1464),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1473),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1459),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1441),
.A2(n_1453),
.B1(n_1443),
.B2(n_1449),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1513),
.A2(n_1522),
.B1(n_1504),
.B2(n_1524),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1488),
.B(n_1490),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1423),
.Y(n_1615)
);

AOI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1439),
.A2(n_1482),
.B1(n_1472),
.B2(n_1507),
.C(n_1470),
.Y(n_1616)
);

O2A1O1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1434),
.A2(n_1486),
.B(n_1485),
.C(n_1468),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1520),
.B(n_1475),
.Y(n_1618)
);

AOI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1537),
.A2(n_1524),
.B(n_1465),
.C(n_1461),
.Y(n_1619)
);

AOI21xp33_ASAP7_75t_L g1620 ( 
.A1(n_1457),
.A2(n_1435),
.B(n_1465),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1432),
.A2(n_1496),
.B1(n_1436),
.B2(n_1459),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1527),
.B(n_1515),
.Y(n_1622)
);

OR2x6_ASAP7_75t_L g1623 ( 
.A(n_1450),
.B(n_1436),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1472),
.A2(n_1495),
.B1(n_1516),
.B2(n_1526),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_SL g1625 ( 
.A1(n_1432),
.A2(n_1496),
.B1(n_1436),
.B2(n_1459),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1537),
.A2(n_1505),
.B1(n_1533),
.B2(n_1557),
.C(n_1476),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1518),
.A2(n_1458),
.B1(n_1555),
.B2(n_1496),
.Y(n_1627)
);

AOI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1514),
.A2(n_1442),
.B(n_1505),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1432),
.A2(n_1467),
.B1(n_1469),
.B2(n_1541),
.Y(n_1629)
);

OAI211xp5_ASAP7_75t_SL g1630 ( 
.A1(n_1476),
.A2(n_1444),
.B(n_1469),
.C(n_1544),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1467),
.A2(n_1543),
.B1(n_1550),
.B2(n_1450),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1467),
.A2(n_1543),
.B1(n_1450),
.B2(n_1444),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1474),
.A2(n_1489),
.B1(n_1532),
.B2(n_1509),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1535),
.A2(n_1544),
.B(n_1500),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1491),
.A2(n_1501),
.B1(n_1494),
.B2(n_1539),
.Y(n_1635)
);

OAI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1543),
.A2(n_1565),
.B1(n_1477),
.B2(n_1481),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1523),
.B(n_1534),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1553),
.Y(n_1638)
);

OA21x2_ASAP7_75t_L g1639 ( 
.A1(n_1548),
.A2(n_1545),
.B(n_1558),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1554),
.B(n_1564),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1560),
.B(n_1566),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1568),
.A2(n_1569),
.B1(n_1551),
.B2(n_1534),
.Y(n_1642)
);

BUFx8_ASAP7_75t_L g1643 ( 
.A(n_1525),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1525),
.A2(n_1559),
.B1(n_1561),
.B2(n_1508),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1559),
.A2(n_1561),
.B(n_1508),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1525),
.A2(n_1567),
.B1(n_1570),
.B2(n_1558),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1546),
.Y(n_1647)
);

AOI21xp33_ASAP7_75t_L g1648 ( 
.A1(n_1570),
.A2(n_1546),
.B(n_1567),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1552),
.A2(n_953),
.B1(n_1531),
.B2(n_1401),
.Y(n_1649)
);

AOI222xp33_ASAP7_75t_L g1650 ( 
.A1(n_1478),
.A2(n_1556),
.B1(n_752),
.B2(n_899),
.C1(n_879),
.C2(n_1401),
.Y(n_1650)
);

AOI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1556),
.A2(n_899),
.B1(n_1401),
.B2(n_761),
.C(n_752),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1422),
.A2(n_1452),
.B1(n_899),
.B2(n_1272),
.Y(n_1652)
);

OAI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_953),
.B2(n_761),
.C(n_773),
.Y(n_1653)
);

OAI31xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1427),
.A2(n_899),
.A3(n_1401),
.B(n_1257),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_953),
.B2(n_761),
.C(n_773),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1422),
.A2(n_1452),
.B1(n_899),
.B2(n_1272),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1437),
.B(n_1542),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1424),
.B(n_686),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1531),
.A2(n_953),
.B1(n_1401),
.B2(n_899),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_1401),
.B2(n_761),
.C(n_752),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1547),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1531),
.A2(n_953),
.B1(n_1401),
.B2(n_899),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1530),
.A2(n_899),
.B1(n_880),
.B2(n_1218),
.Y(n_1663)
);

OAI21xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1502),
.A2(n_1022),
.B(n_1422),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1446),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_1401),
.B2(n_761),
.C(n_752),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1484),
.B(n_1445),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_1022),
.B2(n_1401),
.Y(n_1668)
);

AOI222xp33_ASAP7_75t_L g1669 ( 
.A1(n_1452),
.A2(n_752),
.B1(n_899),
.B2(n_879),
.C1(n_1401),
.C2(n_593),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_953),
.B2(n_665),
.Y(n_1670)
);

OAI221xp5_ASAP7_75t_L g1671 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_953),
.B2(n_761),
.C(n_773),
.Y(n_1671)
);

NOR2xp67_ASAP7_75t_L g1672 ( 
.A(n_1492),
.B(n_906),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1422),
.A2(n_1452),
.B1(n_899),
.B2(n_1272),
.Y(n_1673)
);

AOI222xp33_ASAP7_75t_L g1674 ( 
.A1(n_1452),
.A2(n_752),
.B1(n_899),
.B2(n_879),
.C1(n_1401),
.C2(n_593),
.Y(n_1674)
);

OAI21x1_ASAP7_75t_SL g1675 ( 
.A1(n_1427),
.A2(n_1383),
.B(n_1390),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_1401),
.B2(n_761),
.C(n_752),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_1401),
.B2(n_761),
.C(n_752),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1424),
.B(n_686),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1422),
.A2(n_1452),
.B1(n_899),
.B2(n_1272),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1484),
.B(n_1445),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1484),
.B(n_1445),
.Y(n_1681)
);

AOI211xp5_ASAP7_75t_L g1682 ( 
.A1(n_1427),
.A2(n_899),
.B(n_1401),
.C(n_953),
.Y(n_1682)
);

INVx5_ASAP7_75t_SL g1683 ( 
.A(n_1459),
.Y(n_1683)
);

OAI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_953),
.B2(n_761),
.C(n_773),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_1022),
.B2(n_1401),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1422),
.A2(n_1452),
.B1(n_899),
.B2(n_1272),
.Y(n_1686)
);

BUFx12f_ASAP7_75t_L g1687 ( 
.A(n_1426),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_1401),
.B2(n_761),
.C(n_752),
.Y(n_1688)
);

OAI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1531),
.A2(n_953),
.B1(n_1401),
.B2(n_899),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1484),
.B(n_1445),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1422),
.A2(n_1452),
.B1(n_899),
.B2(n_1272),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_1022),
.B2(n_1401),
.Y(n_1692)
);

AO21x2_ASAP7_75t_L g1693 ( 
.A1(n_1549),
.A2(n_1487),
.B(n_1498),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1445),
.B(n_1462),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_953),
.B2(n_665),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1424),
.B(n_686),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1452),
.A2(n_899),
.B1(n_953),
.B2(n_665),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1623),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1612),
.B(n_1667),
.Y(n_1699)
);

NOR2xp67_ASAP7_75t_L g1700 ( 
.A(n_1647),
.B(n_1645),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1576),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1580),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1612),
.B(n_1680),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_SL g1704 ( 
.A(n_1623),
.B(n_1609),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1681),
.B(n_1690),
.Y(n_1705)
);

BUFx12f_ASAP7_75t_L g1706 ( 
.A(n_1581),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1596),
.B(n_1582),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1582),
.B(n_1639),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1582),
.B(n_1639),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1577),
.B(n_1578),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1614),
.B(n_1693),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1587),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1640),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1693),
.B(n_1648),
.Y(n_1715)
);

INVx5_ASAP7_75t_L g1716 ( 
.A(n_1641),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1694),
.B(n_1618),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1592),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1571),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1633),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1632),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1661),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1633),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1622),
.B(n_1607),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1646),
.B(n_1644),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1634),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1635),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1660),
.A2(n_1666),
.B1(n_1677),
.B2(n_1676),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1653),
.B(n_1655),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1646),
.B(n_1644),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1572),
.B(n_1608),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1573),
.B(n_1616),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1604),
.B(n_1573),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1635),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1629),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1603),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1637),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1574),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1636),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1604),
.B(n_1624),
.Y(n_1740)
);

INVx2_ASAP7_75t_SL g1741 ( 
.A(n_1643),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1626),
.B(n_1593),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1594),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1586),
.B(n_1628),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1643),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1590),
.B(n_1624),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1636),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1575),
.B(n_1642),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1630),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1590),
.B(n_1619),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1575),
.B(n_1579),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1579),
.B(n_1657),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1598),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1589),
.B(n_1588),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1675),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1589),
.B(n_1620),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1631),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1617),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1613),
.B(n_1597),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1638),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1611),
.Y(n_1761)
);

OR2x6_ASAP7_75t_L g1762 ( 
.A(n_1698),
.B(n_1584),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1712),
.B(n_1591),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1711),
.B(n_1625),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1716),
.B(n_1611),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1712),
.B(n_1598),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1711),
.B(n_1625),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1728),
.A2(n_1685),
.B1(n_1668),
.B2(n_1692),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1711),
.B(n_1621),
.Y(n_1769)
);

AOI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1749),
.A2(n_1671),
.B1(n_1684),
.B2(n_1659),
.C(n_1689),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1716),
.B(n_1610),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1701),
.Y(n_1772)
);

AND2x4_ASAP7_75t_SL g1773 ( 
.A(n_1736),
.B(n_1601),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1707),
.B(n_1621),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1729),
.A2(n_1728),
.B1(n_1688),
.B2(n_1669),
.Y(n_1775)
);

OAI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1750),
.A2(n_1697),
.B1(n_1695),
.B2(n_1670),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1707),
.B(n_1585),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1729),
.A2(n_1674),
.B1(n_1673),
.B2(n_1691),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1716),
.B(n_1600),
.Y(n_1779)
);

AOI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1749),
.A2(n_1686),
.B1(n_1679),
.B2(n_1656),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1750),
.A2(n_1659),
.B1(n_1662),
.B2(n_1689),
.C(n_1651),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1756),
.A2(n_1652),
.B1(n_1650),
.B2(n_1692),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1758),
.B(n_1699),
.Y(n_1783)
);

OR2x6_ASAP7_75t_SL g1784 ( 
.A(n_1731),
.B(n_1605),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1701),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1708),
.B(n_1615),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1714),
.Y(n_1787)
);

OAI33xp33_ASAP7_75t_L g1788 ( 
.A1(n_1731),
.A2(n_1662),
.A3(n_1649),
.B1(n_1602),
.B2(n_1663),
.B3(n_1627),
.Y(n_1788)
);

BUFx10_ASAP7_75t_L g1789 ( 
.A(n_1741),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1717),
.B(n_1724),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1708),
.B(n_1606),
.Y(n_1791)
);

INVxp67_ASAP7_75t_SL g1792 ( 
.A(n_1712),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1716),
.B(n_1672),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1702),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1704),
.A2(n_1649),
.B(n_1664),
.Y(n_1795)
);

INVxp67_ASAP7_75t_L g1796 ( 
.A(n_1724),
.Y(n_1796)
);

INVx4_ASAP7_75t_SL g1797 ( 
.A(n_1741),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1719),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1708),
.B(n_1683),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1752),
.B(n_1683),
.Y(n_1800)
);

OAI33xp33_ASAP7_75t_L g1801 ( 
.A1(n_1731),
.A2(n_1654),
.A3(n_1665),
.B1(n_1682),
.B2(n_1685),
.B3(n_1658),
.Y(n_1801)
);

NAND4xp25_ASAP7_75t_L g1802 ( 
.A(n_1758),
.B(n_1678),
.C(n_1696),
.D(n_1599),
.Y(n_1802)
);

OAI31xp33_ASAP7_75t_L g1803 ( 
.A1(n_1740),
.A2(n_1595),
.A3(n_1683),
.B(n_1687),
.Y(n_1803)
);

NAND2xp33_ASAP7_75t_R g1804 ( 
.A(n_1753),
.B(n_1726),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1746),
.A2(n_1753),
.B1(n_1743),
.B2(n_1739),
.Y(n_1805)
);

AOI33xp33_ASAP7_75t_L g1806 ( 
.A1(n_1744),
.A2(n_1742),
.A3(n_1732),
.B1(n_1743),
.B2(n_1756),
.B3(n_1754),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1717),
.B(n_1705),
.Y(n_1807)
);

AOI31xp33_ASAP7_75t_L g1808 ( 
.A1(n_1746),
.A2(n_1740),
.A3(n_1743),
.B(n_1721),
.Y(n_1808)
);

OAI31xp33_ASAP7_75t_L g1809 ( 
.A1(n_1740),
.A2(n_1753),
.A3(n_1756),
.B(n_1739),
.Y(n_1809)
);

NAND4xp25_ASAP7_75t_L g1810 ( 
.A(n_1742),
.B(n_1726),
.C(n_1744),
.D(n_1732),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1705),
.B(n_1699),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1722),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1703),
.B(n_1737),
.Y(n_1813)
);

OA222x2_ASAP7_75t_L g1814 ( 
.A1(n_1733),
.A2(n_1703),
.B1(n_1734),
.B2(n_1727),
.C1(n_1720),
.C2(n_1723),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1722),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1772),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1772),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1774),
.B(n_1709),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1789),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1785),
.Y(n_1820)
);

INVxp67_ASAP7_75t_L g1821 ( 
.A(n_1813),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1785),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1774),
.B(n_1786),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1794),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1792),
.B(n_1715),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1794),
.Y(n_1826)
);

NAND2xp33_ASAP7_75t_R g1827 ( 
.A(n_1793),
.B(n_1726),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1777),
.B(n_1709),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1764),
.B(n_1710),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1798),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1764),
.B(n_1710),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1763),
.B(n_1715),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1767),
.B(n_1713),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1765),
.B(n_1716),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1763),
.B(n_1715),
.Y(n_1835)
);

NOR2x1_ASAP7_75t_L g1836 ( 
.A(n_1810),
.B(n_1700),
.Y(n_1836)
);

INVx4_ASAP7_75t_SL g1837 ( 
.A(n_1793),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1798),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1767),
.B(n_1713),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1769),
.B(n_1716),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1769),
.B(n_1716),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1811),
.B(n_1738),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1789),
.Y(n_1843)
);

OR2x6_ASAP7_75t_L g1844 ( 
.A(n_1779),
.B(n_1698),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1796),
.B(n_1738),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1799),
.B(n_1791),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1766),
.B(n_1714),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1766),
.B(n_1718),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1787),
.B(n_1742),
.Y(n_1849)
);

OAI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1775),
.A2(n_1744),
.B(n_1732),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1812),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1790),
.B(n_1737),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1816),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1816),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1818),
.B(n_1814),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1837),
.B(n_1793),
.Y(n_1856)
);

INVx3_ASAP7_75t_SL g1857 ( 
.A(n_1843),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1818),
.B(n_1814),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1817),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1817),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1842),
.B(n_1783),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1842),
.B(n_1808),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1851),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1820),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1818),
.B(n_1800),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1851),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1820),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1829),
.B(n_1831),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1822),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1822),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1851),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1845),
.B(n_1808),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1824),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1850),
.B(n_1706),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1824),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1829),
.B(n_1800),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1845),
.B(n_1807),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1829),
.B(n_1771),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1821),
.B(n_1810),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1850),
.B(n_1706),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1847),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1826),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1826),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1830),
.Y(n_1884)
);

AOI322xp5_ASAP7_75t_L g1885 ( 
.A1(n_1836),
.A2(n_1778),
.A3(n_1782),
.B1(n_1780),
.B2(n_1776),
.C1(n_1781),
.C2(n_1770),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1821),
.B(n_1809),
.Y(n_1886)
);

NOR2x1_ASAP7_75t_SL g1887 ( 
.A(n_1844),
.B(n_1762),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1848),
.B(n_1815),
.Y(n_1888)
);

OR2x6_ASAP7_75t_L g1889 ( 
.A(n_1836),
.B(n_1795),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1847),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1838),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1848),
.B(n_1815),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1881),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1889),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1853),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1853),
.Y(n_1896)
);

NOR2xp67_ASAP7_75t_L g1897 ( 
.A(n_1856),
.B(n_1706),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1854),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1866),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1890),
.B(n_1848),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1866),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1854),
.Y(n_1902)
);

AND2x2_ASAP7_75t_SL g1903 ( 
.A(n_1874),
.B(n_1806),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1866),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1879),
.B(n_1886),
.Y(n_1905)
);

NOR2x1_ASAP7_75t_L g1906 ( 
.A(n_1889),
.B(n_1849),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1856),
.B(n_1837),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1861),
.B(n_1849),
.Y(n_1908)
);

NAND2xp33_ASAP7_75t_R g1909 ( 
.A(n_1889),
.B(n_1739),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1889),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1889),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1862),
.B(n_1833),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1857),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1888),
.B(n_1832),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1859),
.Y(n_1915)
);

NAND2xp33_ASAP7_75t_SL g1916 ( 
.A(n_1857),
.B(n_1804),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1888),
.B(n_1832),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1868),
.B(n_1837),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_SL g1919 ( 
.A(n_1880),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1872),
.B(n_1784),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1859),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1868),
.B(n_1837),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1860),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1860),
.Y(n_1924)
);

AOI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1855),
.A2(n_1801),
.B1(n_1768),
.B2(n_1805),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1877),
.B(n_1833),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1865),
.Y(n_1927)
);

NOR3xp33_ASAP7_75t_L g1928 ( 
.A(n_1855),
.B(n_1802),
.C(n_1788),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1865),
.B(n_1847),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1892),
.B(n_1832),
.Y(n_1930)
);

NOR2xp67_ASAP7_75t_L g1931 ( 
.A(n_1856),
.B(n_1840),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1892),
.B(n_1835),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1856),
.B(n_1858),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1864),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1864),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1876),
.B(n_1835),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1876),
.B(n_1833),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1893),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1895),
.Y(n_1939)
);

INVxp67_ASAP7_75t_SL g1940 ( 
.A(n_1909),
.Y(n_1940)
);

AOI31xp33_ASAP7_75t_L g1941 ( 
.A1(n_1920),
.A2(n_1858),
.A3(n_1741),
.B(n_1745),
.Y(n_1941)
);

NAND3xp33_ASAP7_75t_L g1942 ( 
.A(n_1920),
.B(n_1885),
.C(n_1809),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1896),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1928),
.B(n_1839),
.Y(n_1944)
);

AOI322xp5_ASAP7_75t_L g1945 ( 
.A1(n_1925),
.A2(n_1839),
.A3(n_1831),
.B1(n_1784),
.B2(n_1885),
.C1(n_1721),
.C2(n_1828),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1898),
.Y(n_1946)
);

NAND4xp75_ASAP7_75t_L g1947 ( 
.A(n_1906),
.B(n_1803),
.C(n_1745),
.D(n_1700),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1919),
.A2(n_1805),
.B1(n_1857),
.B2(n_1795),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1903),
.B(n_1839),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1903),
.A2(n_1802),
.B(n_1803),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1905),
.B(n_1823),
.Y(n_1951)
);

AOI21xp33_ASAP7_75t_L g1952 ( 
.A1(n_1909),
.A2(n_1827),
.B(n_1757),
.Y(n_1952)
);

NAND3xp33_ASAP7_75t_SL g1953 ( 
.A(n_1916),
.B(n_1754),
.C(n_1760),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1916),
.A2(n_1827),
.B1(n_1754),
.B2(n_1725),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1905),
.A2(n_1844),
.B1(n_1748),
.B2(n_1762),
.Y(n_1955)
);

AOI21xp33_ASAP7_75t_L g1956 ( 
.A1(n_1910),
.A2(n_1757),
.B(n_1835),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1908),
.B(n_1852),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1902),
.Y(n_1958)
);

INVx1_ASAP7_75t_SL g1959 ( 
.A(n_1913),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1915),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1908),
.B(n_1852),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1937),
.B(n_1823),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1933),
.Y(n_1963)
);

O2A1O1Ixp33_ASAP7_75t_SL g1964 ( 
.A1(n_1911),
.A2(n_1745),
.B(n_1760),
.C(n_1819),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1926),
.B(n_1823),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1897),
.A2(n_1730),
.B1(n_1725),
.B2(n_1748),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1921),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1912),
.B(n_1825),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1927),
.B(n_1846),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_SL g1970 ( 
.A(n_1894),
.B(n_1907),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1907),
.A2(n_1725),
.B(n_1730),
.Y(n_1971)
);

OAI321xp33_ASAP7_75t_L g1972 ( 
.A1(n_1933),
.A2(n_1762),
.A3(n_1733),
.B1(n_1730),
.B2(n_1751),
.C(n_1755),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_1900),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1907),
.B(n_1887),
.Y(n_1974)
);

AOI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1942),
.A2(n_1748),
.B1(n_1735),
.B2(n_1751),
.Y(n_1975)
);

AOI211xp5_ASAP7_75t_SL g1976 ( 
.A1(n_1940),
.A2(n_1931),
.B(n_1918),
.C(n_1922),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1974),
.B(n_1918),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1974),
.B(n_1922),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1938),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1938),
.Y(n_1980)
);

INVx1_ASAP7_75t_SL g1981 ( 
.A(n_1959),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1945),
.B(n_1900),
.Y(n_1982)
);

AOI221xp5_ASAP7_75t_L g1983 ( 
.A1(n_1940),
.A2(n_1924),
.B1(n_1923),
.B2(n_1934),
.C(n_1935),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1939),
.Y(n_1984)
);

OAI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1950),
.A2(n_1929),
.B1(n_1936),
.B2(n_1844),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1963),
.B(n_1887),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1963),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1943),
.Y(n_1988)
);

AOI211xp5_ASAP7_75t_L g1989 ( 
.A1(n_1953),
.A2(n_1948),
.B(n_1944),
.C(n_1952),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1946),
.Y(n_1990)
);

OAI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1941),
.A2(n_1844),
.B1(n_1834),
.B2(n_1748),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1973),
.B(n_1878),
.Y(n_1992)
);

AOI222xp33_ASAP7_75t_L g1993 ( 
.A1(n_1953),
.A2(n_1751),
.B1(n_1748),
.B2(n_1735),
.C1(n_1759),
.C2(n_1718),
.Y(n_1993)
);

OAI21xp33_ASAP7_75t_L g1994 ( 
.A1(n_1949),
.A2(n_1733),
.B(n_1759),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1958),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1960),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1971),
.B(n_1846),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1972),
.A2(n_1704),
.B(n_1760),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1967),
.Y(n_1999)
);

INVxp67_ASAP7_75t_L g2000 ( 
.A(n_1970),
.Y(n_2000)
);

O2A1O1Ixp33_ASAP7_75t_L g2001 ( 
.A1(n_1964),
.A2(n_1747),
.B(n_1825),
.C(n_1901),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1980),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1977),
.B(n_1951),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1979),
.B(n_1969),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1981),
.B(n_1966),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1982),
.A2(n_1989),
.B(n_1994),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1977),
.B(n_1954),
.Y(n_2007)
);

XNOR2xp5_ASAP7_75t_L g2008 ( 
.A(n_1975),
.B(n_1947),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1979),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1987),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_2000),
.A2(n_1955),
.B1(n_1964),
.B2(n_1956),
.Y(n_2011)
);

INVxp67_ASAP7_75t_SL g2012 ( 
.A(n_2001),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1993),
.B(n_1957),
.Y(n_2013)
);

OAI21xp5_ASAP7_75t_SL g2014 ( 
.A1(n_1975),
.A2(n_1968),
.B(n_1773),
.Y(n_2014)
);

BUFx2_ASAP7_75t_L g2015 ( 
.A(n_1987),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1996),
.Y(n_2016)
);

INVx1_ASAP7_75t_SL g2017 ( 
.A(n_1978),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1978),
.B(n_1962),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1996),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1994),
.B(n_1961),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1999),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1999),
.Y(n_2022)
);

OAI221xp5_ASAP7_75t_L g2023 ( 
.A1(n_2008),
.A2(n_1976),
.B1(n_1983),
.B2(n_1985),
.C(n_1998),
.Y(n_2023)
);

NOR2x1_ASAP7_75t_SL g2024 ( 
.A(n_2002),
.B(n_1984),
.Y(n_2024)
);

OAI21xp33_ASAP7_75t_L g2025 ( 
.A1(n_2006),
.A2(n_1992),
.B(n_1997),
.Y(n_2025)
);

AND4x1_ASAP7_75t_L g2026 ( 
.A(n_2005),
.B(n_1995),
.C(n_1984),
.D(n_1988),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_2015),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_2012),
.A2(n_1991),
.B1(n_1992),
.B2(n_1986),
.Y(n_2028)
);

NAND3xp33_ASAP7_75t_L g2029 ( 
.A(n_2008),
.B(n_1995),
.C(n_1988),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2017),
.B(n_1986),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2007),
.B(n_1990),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_2020),
.B(n_1990),
.Y(n_2032)
);

NOR3xp33_ASAP7_75t_L g2033 ( 
.A(n_2014),
.B(n_1965),
.C(n_1904),
.Y(n_2033)
);

NOR2x1_ASAP7_75t_SL g2034 ( 
.A(n_2004),
.B(n_1760),
.Y(n_2034)
);

AOI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_2023),
.A2(n_2013),
.B1(n_2009),
.B2(n_2007),
.C(n_2019),
.Y(n_2035)
);

O2A1O1Ixp33_ASAP7_75t_L g2036 ( 
.A1(n_2029),
.A2(n_2013),
.B(n_2009),
.C(n_2022),
.Y(n_2036)
);

NOR2x1_ASAP7_75t_L g2037 ( 
.A(n_2029),
.B(n_2027),
.Y(n_2037)
);

AOI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_2032),
.A2(n_2021),
.B1(n_2016),
.B2(n_2011),
.C(n_2015),
.Y(n_2038)
);

NAND3xp33_ASAP7_75t_SL g2039 ( 
.A(n_2026),
.B(n_2004),
.C(n_2010),
.Y(n_2039)
);

AOI222xp33_ASAP7_75t_SL g2040 ( 
.A1(n_2024),
.A2(n_2003),
.B1(n_2018),
.B2(n_1904),
.C1(n_1901),
.C2(n_1899),
.Y(n_2040)
);

OAI321xp33_ASAP7_75t_L g2041 ( 
.A1(n_2025),
.A2(n_2003),
.A3(n_2018),
.B1(n_1917),
.B2(n_1932),
.C(n_1930),
.Y(n_2041)
);

AOI221xp5_ASAP7_75t_L g2042 ( 
.A1(n_2031),
.A2(n_1899),
.B1(n_1867),
.B2(n_1869),
.C(n_1870),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_2030),
.B(n_1914),
.Y(n_2043)
);

AOI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2028),
.A2(n_1882),
.B1(n_1875),
.B2(n_1873),
.C(n_1870),
.Y(n_2044)
);

O2A1O1Ixp33_ASAP7_75t_L g2045 ( 
.A1(n_2033),
.A2(n_1932),
.B(n_1917),
.C(n_1914),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_2037),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2035),
.A2(n_1797),
.B1(n_1834),
.B2(n_1841),
.Y(n_2047)
);

AOI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_2036),
.A2(n_2034),
.B(n_1871),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_2039),
.B(n_1930),
.Y(n_2049)
);

NOR2xp67_ASAP7_75t_L g2050 ( 
.A(n_2041),
.B(n_1871),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_2043),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2046),
.B(n_2038),
.Y(n_2052)
);

NOR2x1_ASAP7_75t_L g2053 ( 
.A(n_2051),
.B(n_2045),
.Y(n_2053)
);

AND2x4_ASAP7_75t_L g2054 ( 
.A(n_2049),
.B(n_2040),
.Y(n_2054)
);

OAI211xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2047),
.A2(n_2044),
.B(n_2042),
.C(n_1825),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2050),
.Y(n_2056)
);

BUFx12f_ASAP7_75t_L g2057 ( 
.A(n_2048),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2046),
.Y(n_2058)
);

NOR3xp33_ASAP7_75t_L g2059 ( 
.A(n_2052),
.B(n_1841),
.C(n_1840),
.Y(n_2059)
);

NAND3xp33_ASAP7_75t_SL g2060 ( 
.A(n_2056),
.B(n_1840),
.C(n_1841),
.Y(n_2060)
);

AOI31xp33_ASAP7_75t_SL g2061 ( 
.A1(n_2053),
.A2(n_1871),
.A3(n_1863),
.B(n_1761),
.Y(n_2061)
);

AND2x4_ASAP7_75t_L g2062 ( 
.A(n_2058),
.B(n_1837),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_2054),
.A2(n_1797),
.B1(n_1834),
.B2(n_1837),
.Y(n_2063)
);

NAND4xp25_ASAP7_75t_L g2064 ( 
.A(n_2054),
.B(n_1793),
.C(n_1834),
.D(n_1759),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2059),
.B(n_2057),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2062),
.B(n_1878),
.Y(n_2066)
);

OAI221xp5_ASAP7_75t_L g2067 ( 
.A1(n_2063),
.A2(n_2055),
.B1(n_1819),
.B2(n_1844),
.C(n_1875),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_2060),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2068),
.Y(n_2069)
);

OAI21xp33_ASAP7_75t_L g2070 ( 
.A1(n_2069),
.A2(n_2064),
.B(n_2065),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2070),
.Y(n_2071)
);

CKINVDCx20_ASAP7_75t_R g2072 ( 
.A(n_2070),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_2071),
.A2(n_2067),
.B(n_2066),
.Y(n_2073)
);

OAI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_2072),
.A2(n_2061),
.B(n_1863),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2074),
.Y(n_2075)
);

AOI221xp5_ASAP7_75t_L g2076 ( 
.A1(n_2073),
.A2(n_1882),
.B1(n_1867),
.B2(n_1869),
.C(n_1873),
.Y(n_2076)
);

INVxp67_ASAP7_75t_SL g2077 ( 
.A(n_2075),
.Y(n_2077)
);

AOI221xp5_ASAP7_75t_L g2078 ( 
.A1(n_2077),
.A2(n_2076),
.B1(n_1883),
.B2(n_1891),
.C(n_1884),
.Y(n_2078)
);

AOI211xp5_ASAP7_75t_L g2079 ( 
.A1(n_2078),
.A2(n_1883),
.B(n_1891),
.C(n_1884),
.Y(n_2079)
);


endmodule