module fake_aes_1176_n_1273 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1273);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1273;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_411;
wire n_860;
wire n_1208;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_7), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_14), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_288), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_34), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_80), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_315), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_7), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_53), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_143), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_237), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_236), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_159), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_272), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_67), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_121), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_163), .Y(n_335) );
INVxp33_ASAP7_75t_L g336 ( .A(n_281), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_264), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_145), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_197), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_242), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_199), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_301), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_188), .Y(n_343) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_319), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_100), .Y(n_345) );
NOR2xp67_ASAP7_75t_L g346 ( .A(n_214), .B(n_171), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_311), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_273), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_61), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_81), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_232), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_278), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_148), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_126), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_26), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_286), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_179), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_147), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_310), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_67), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_146), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_19), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_202), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_102), .Y(n_364) );
INVxp33_ASAP7_75t_L g365 ( .A(n_261), .Y(n_365) );
CKINVDCx14_ASAP7_75t_R g366 ( .A(n_204), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_157), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_133), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_213), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_98), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_30), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_183), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_275), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_140), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_112), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_122), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_175), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_230), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_114), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_17), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_72), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_42), .Y(n_382) );
CKINVDCx16_ASAP7_75t_R g383 ( .A(n_172), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_184), .Y(n_384) );
BUFx5_ASAP7_75t_L g385 ( .A(n_176), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_131), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_309), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_33), .Y(n_388) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_38), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_249), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_39), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_50), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_72), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_37), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_2), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_0), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_123), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_218), .Y(n_398) );
CKINVDCx14_ASAP7_75t_R g399 ( .A(n_40), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_190), .B(n_70), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_285), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_127), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_52), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_266), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_262), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_151), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_56), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_305), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_120), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_246), .Y(n_410) );
CKINVDCx14_ASAP7_75t_R g411 ( .A(n_225), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_79), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_160), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_60), .Y(n_414) );
NOR2xp67_ASAP7_75t_L g415 ( .A(n_292), .B(n_36), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_86), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_43), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_24), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_297), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_289), .Y(n_420) );
CKINVDCx14_ASAP7_75t_R g421 ( .A(n_189), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_25), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_318), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_174), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_101), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_201), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_209), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_47), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_166), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_110), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_260), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_71), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_233), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_191), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_6), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_215), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_68), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_75), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_193), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_2), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_103), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_299), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_13), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_274), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_83), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_251), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_222), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_200), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_267), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_39), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_280), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_149), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_279), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_287), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_156), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_51), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_84), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_164), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_139), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_68), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_6), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_256), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_226), .Y(n_463) );
BUFx10_ASAP7_75t_L g464 ( .A(n_51), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_115), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_259), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_20), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_86), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_303), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_141), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_40), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_194), .Y(n_472) );
BUFx2_ASAP7_75t_L g473 ( .A(n_282), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_15), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_153), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_206), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_219), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_15), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_63), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_41), .Y(n_480) );
INVxp33_ASAP7_75t_SL g481 ( .A(n_271), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_24), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_399), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_464), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_385), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_385), .Y(n_486) );
NAND2xp33_ASAP7_75t_L g487 ( .A(n_385), .B(n_113), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_385), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_385), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_351), .Y(n_490) );
BUFx8_ASAP7_75t_L g491 ( .A(n_384), .Y(n_491) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_473), .B(n_317), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_382), .Y(n_493) );
AOI22x1_ASAP7_75t_SL g494 ( .A1(n_320), .A2(n_3), .B1(n_0), .B2(n_1), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_351), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_385), .Y(n_496) );
OAI22x1_ASAP7_75t_R g497 ( .A1(n_320), .A2(n_5), .B1(n_1), .B2(n_4), .Y(n_497) );
AND2x2_ASAP7_75t_SL g498 ( .A(n_328), .B(n_316), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_376), .B(n_321), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_382), .Y(n_500) );
NAND2xp33_ASAP7_75t_L g501 ( .A(n_385), .B(n_116), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_435), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_351), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_435), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_351), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_450), .Y(n_506) );
NAND2xp33_ASAP7_75t_SL g507 ( .A(n_336), .B(n_4), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_413), .Y(n_508) );
INVx3_ASAP7_75t_L g509 ( .A(n_327), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_413), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_450), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_480), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g513 ( .A1(n_407), .A2(n_9), .B1(n_5), .B2(n_8), .Y(n_513) );
OAI22x1_ASAP7_75t_R g514 ( .A1(n_407), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_413), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_413), .Y(n_516) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_325), .A2(n_118), .B(n_117), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_336), .B(n_11), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_327), .B(n_11), .Y(n_520) );
INVx5_ASAP7_75t_L g521 ( .A(n_419), .Y(n_521) );
INVx5_ASAP7_75t_L g522 ( .A(n_419), .Y(n_522) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_419), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_419), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_520), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_485), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_509), .B(n_365), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_483), .B(n_365), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_485), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_485), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_498), .A2(n_324), .B1(n_333), .B2(n_326), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_490), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_509), .B(n_325), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_486), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_499), .B(n_366), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_490), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_484), .B(n_465), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_490), .Y(n_538) );
INVx4_ASAP7_75t_SL g539 ( .A(n_520), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_486), .Y(n_540) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_497), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_490), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_499), .B(n_366), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_486), .Y(n_544) );
BUFx3_ASAP7_75t_L g545 ( .A(n_509), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_487), .B(n_331), .C(n_322), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_490), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_490), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_491), .B(n_383), .Y(n_549) );
INVx4_ASAP7_75t_L g550 ( .A(n_520), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_495), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_509), .B(n_330), .Y(n_552) );
INVx3_ASAP7_75t_L g553 ( .A(n_520), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_498), .A2(n_350), .B1(n_360), .B2(n_345), .Y(n_554) );
BUFx3_ASAP7_75t_L g555 ( .A(n_517), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_495), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_493), .B(n_330), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_488), .B(n_489), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_498), .A2(n_362), .B1(n_371), .B2(n_364), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_488), .Y(n_560) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_495), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_493), .B(n_404), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_491), .B(n_444), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_495), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_491), .B(n_472), .Y(n_565) );
AND2x6_ASAP7_75t_L g566 ( .A(n_519), .B(n_339), .Y(n_566) );
AND2x6_ASAP7_75t_L g567 ( .A(n_488), .B(n_339), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_500), .B(n_404), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_535), .B(n_492), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_555), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_527), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_535), .B(n_492), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_535), .B(n_492), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_531), .A2(n_507), .B1(n_399), .B2(n_491), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_543), .B(n_489), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_543), .B(n_489), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_541), .B(n_513), .C(n_418), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_528), .B(n_389), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_527), .A2(n_430), .B1(n_471), .B2(n_437), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_528), .B(n_464), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_557), .Y(n_581) );
INVx4_ASAP7_75t_L g582 ( .A(n_539), .Y(n_582) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_550), .B(n_380), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_528), .B(n_481), .Y(n_584) );
BUFx8_ASAP7_75t_L g585 ( .A(n_566), .Y(n_585) );
NAND2x1p5_ASAP7_75t_L g586 ( .A(n_550), .B(n_381), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_550), .B(n_354), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_525), .B(n_496), .Y(n_588) );
NOR3xp33_ASAP7_75t_L g589 ( .A(n_549), .B(n_513), .C(n_443), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_531), .A2(n_344), .B1(n_420), .B2(n_347), .Y(n_590) );
BUFx2_ASAP7_75t_L g591 ( .A(n_539), .Y(n_591) );
NOR2x1p5_ASAP7_75t_L g592 ( .A(n_563), .B(n_323), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_568), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_545), .Y(n_594) );
BUFx12f_ASAP7_75t_L g595 ( .A(n_567), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_568), .Y(n_596) );
OR2x6_ASAP7_75t_L g597 ( .A(n_565), .B(n_514), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_554), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_539), .B(n_354), .Y(n_599) );
BUFx2_ASAP7_75t_L g600 ( .A(n_539), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_559), .A2(n_431), .B1(n_355), .B2(n_422), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_525), .Y(n_602) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_555), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_533), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_525), .B(n_496), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_539), .B(n_387), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_525), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_553), .B(n_496), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_537), .B(n_553), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_555), .A2(n_501), .B(n_517), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_553), .B(n_387), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_553), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_559), .A2(n_414), .B1(n_403), .B2(n_411), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_553), .B(n_436), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_526), .B(n_436), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_533), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_566), .B(n_453), .Y(n_617) );
NAND2xp33_ASAP7_75t_L g618 ( .A(n_566), .B(n_455), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_552), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_526), .B(n_455), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_562), .B(n_464), .Y(n_622) );
OR2x6_ASAP7_75t_L g623 ( .A(n_546), .B(n_514), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_567), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_566), .A2(n_414), .B1(n_403), .B2(n_411), .Y(n_625) );
AND2x4_ASAP7_75t_SL g626 ( .A(n_529), .B(n_437), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_566), .B(n_421), .Y(n_627) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_567), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_558), .Y(n_629) );
OR2x6_ASAP7_75t_L g630 ( .A(n_530), .B(n_494), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_566), .A2(n_421), .B1(n_388), .B2(n_392), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_566), .A2(n_457), .B1(n_393), .B2(n_417), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_566), .Y(n_633) );
NAND2xp33_ASAP7_75t_L g634 ( .A(n_566), .B(n_329), .Y(n_634) );
INVx5_ASAP7_75t_L g635 ( .A(n_567), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_530), .B(n_517), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_534), .A2(n_391), .B1(n_395), .B2(n_394), .Y(n_637) );
INVx4_ASAP7_75t_L g638 ( .A(n_560), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_560), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_560), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_610), .A2(n_544), .B(n_540), .Y(n_641) );
CKINVDCx8_ASAP7_75t_R g642 ( .A(n_597), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_590), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_581), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_604), .B(n_334), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_626), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_578), .B(n_471), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_571), .B(n_540), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_590), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_582), .B(n_400), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_620), .B(n_338), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_583), .Y(n_652) );
OA22x2_ASAP7_75t_L g653 ( .A1(n_597), .A2(n_494), .B1(n_457), .B2(n_456), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_636), .A2(n_544), .B(n_560), .Y(n_654) );
INVxp67_ASAP7_75t_L g655 ( .A(n_580), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_SL g656 ( .A1(n_609), .A2(n_335), .B(n_337), .C(n_332), .Y(n_656) );
BUFx8_ASAP7_75t_SL g657 ( .A(n_630), .Y(n_657) );
INVx1_ASAP7_75t_SL g658 ( .A(n_616), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_593), .A2(n_396), .B(n_425), .C(n_416), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_569), .A2(n_567), .B1(n_428), .B2(n_432), .Y(n_660) );
INVx3_ASAP7_75t_L g661 ( .A(n_582), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_592), .B(n_370), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_596), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_619), .B(n_343), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_575), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_588), .A2(n_341), .B(n_340), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_572), .A2(n_567), .B1(n_440), .B2(n_441), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_598), .A2(n_438), .B1(n_460), .B2(n_445), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_622), .B(n_461), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_575), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_572), .B(n_474), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_586), .B(n_368), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_576), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_573), .A2(n_468), .B(n_478), .C(n_467), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_584), .B(n_479), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_576), .A2(n_504), .B(n_506), .C(n_502), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_601), .A2(n_374), .B(n_372), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_602), .A2(n_415), .B(n_504), .C(n_502), .Y(n_678) );
OAI21x1_ASAP7_75t_L g679 ( .A1(n_588), .A2(n_536), .B(n_532), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_589), .A2(n_511), .B(n_512), .C(n_506), .Y(n_680) );
NAND3xp33_ASAP7_75t_SL g681 ( .A(n_574), .B(n_379), .C(n_348), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_SL g682 ( .A1(n_633), .A2(n_352), .B(n_353), .C(n_342), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_638), .Y(n_683) );
AND2x4_ASAP7_75t_L g684 ( .A(n_591), .B(n_511), .Y(n_684) );
INVx2_ASAP7_75t_SL g685 ( .A(n_586), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_605), .A2(n_357), .B(n_356), .Y(n_686) );
NAND2x1p5_ASAP7_75t_L g687 ( .A(n_600), .B(n_512), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_615), .B(n_377), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_605), .A2(n_359), .B(n_358), .Y(n_689) );
NAND3xp33_ASAP7_75t_SL g690 ( .A(n_577), .B(n_408), .C(n_398), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_607), .A2(n_518), .B(n_361), .C(n_367), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_608), .A2(n_614), .B(n_611), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_621), .B(n_423), .Y(n_693) );
OAI22xp5_ASAP7_75t_SL g694 ( .A1(n_630), .A2(n_451), .B1(n_476), .B2(n_448), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_608), .A2(n_369), .B(n_363), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_621), .B(n_477), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_611), .B(n_349), .Y(n_697) );
O2A1O1Ixp5_ASAP7_75t_L g698 ( .A1(n_599), .A2(n_433), .B(n_463), .C(n_424), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_632), .A2(n_373), .B(n_378), .C(n_375), .Y(n_699) );
O2A1O1Ixp5_ASAP7_75t_L g700 ( .A1(n_606), .A2(n_475), .B(n_390), .C(n_401), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_614), .B(n_349), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_613), .A2(n_402), .B1(n_406), .B2(n_397), .Y(n_702) );
OR2x6_ASAP7_75t_L g703 ( .A(n_623), .B(n_349), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_612), .A2(n_410), .B(n_409), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_638), .Y(n_705) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_570), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_587), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_595), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_631), .A2(n_426), .B1(n_429), .B2(n_427), .Y(n_709) );
BUFx2_ASAP7_75t_L g710 ( .A(n_585), .Y(n_710) );
INVx4_ASAP7_75t_L g711 ( .A(n_635), .Y(n_711) );
NOR2xp67_ASAP7_75t_L g712 ( .A(n_637), .B(n_12), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_570), .B(n_434), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_SL g714 ( .A1(n_625), .A2(n_503), .B(n_510), .C(n_508), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_617), .B(n_412), .Y(n_715) );
O2A1O1Ixp33_ASAP7_75t_L g716 ( .A1(n_618), .A2(n_442), .B(n_446), .C(n_439), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_627), .A2(n_449), .B(n_447), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_634), .A2(n_454), .B(n_452), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_629), .A2(n_459), .B(n_458), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_570), .B(n_462), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_639), .B(n_412), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g722 ( .A1(n_640), .A2(n_466), .B(n_470), .C(n_469), .Y(n_722) );
AO32x1_ASAP7_75t_L g723 ( .A1(n_594), .A2(n_508), .A3(n_515), .B1(n_510), .B2(n_503), .Y(n_723) );
NOR2xp33_ASAP7_75t_SL g724 ( .A(n_603), .B(n_346), .Y(n_724) );
AO32x2_ASAP7_75t_L g725 ( .A1(n_585), .A2(n_516), .A3(n_523), .B1(n_505), .B2(n_495), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_628), .Y(n_726) );
INVx3_ASAP7_75t_L g727 ( .A(n_628), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_624), .A2(n_475), .B(n_532), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_635), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_635), .B(n_482), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g731 ( .A1(n_581), .A2(n_405), .B(n_386), .C(n_503), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_569), .A2(n_482), .B1(n_405), .B2(n_386), .Y(n_732) );
INVx1_ASAP7_75t_SL g733 ( .A(n_604), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_572), .B(n_12), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_638), .Y(n_735) );
NAND2xp33_ASAP7_75t_SL g736 ( .A(n_590), .B(n_508), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_638), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_604), .B(n_521), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_610), .A2(n_538), .B(n_536), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_610), .A2(n_542), .B(n_538), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_610), .A2(n_542), .B(n_538), .Y(n_741) );
BUFx2_ASAP7_75t_L g742 ( .A(n_583), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_604), .B(n_521), .Y(n_743) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_590), .Y(n_744) );
O2A1O1Ixp33_ASAP7_75t_L g745 ( .A1(n_572), .A2(n_515), .B(n_524), .C(n_510), .Y(n_745) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_570), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g747 ( .A1(n_581), .A2(n_524), .B(n_515), .C(n_505), .Y(n_747) );
OAI21xp5_ASAP7_75t_L g748 ( .A1(n_692), .A2(n_524), .B(n_542), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_733), .B(n_13), .Y(n_749) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_706), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g751 ( .A1(n_734), .A2(n_505), .B(n_516), .C(n_495), .Y(n_751) );
OAI21x1_ASAP7_75t_L g752 ( .A1(n_679), .A2(n_548), .B(n_547), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_658), .Y(n_753) );
NAND2x1p5_ASAP7_75t_L g754 ( .A(n_733), .B(n_521), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_644), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g756 ( .A1(n_674), .A2(n_516), .B(n_523), .C(n_505), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_641), .A2(n_548), .B(n_547), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_655), .B(n_16), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_654), .A2(n_564), .B(n_547), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_663), .Y(n_760) );
AO21x1_ASAP7_75t_L g761 ( .A1(n_697), .A2(n_523), .B(n_516), .Y(n_761) );
AO31x2_ASAP7_75t_L g762 ( .A1(n_678), .A2(n_731), .A3(n_747), .B(n_691), .Y(n_762) );
INVxp67_ASAP7_75t_L g763 ( .A(n_647), .Y(n_763) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_706), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_665), .A2(n_522), .B1(n_521), .B2(n_18), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g766 ( .A1(n_659), .A2(n_18), .B(n_16), .C(n_17), .Y(n_766) );
INVx3_ASAP7_75t_SL g767 ( .A(n_646), .Y(n_767) );
OR2x6_ASAP7_75t_L g768 ( .A(n_703), .B(n_19), .Y(n_768) );
OA21x2_ASAP7_75t_L g769 ( .A1(n_739), .A2(n_522), .B(n_551), .Y(n_769) );
AND2x4_ASAP7_75t_L g770 ( .A(n_673), .B(n_20), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_740), .A2(n_556), .B(n_551), .Y(n_771) );
NOR2xp33_ASAP7_75t_SL g772 ( .A(n_657), .B(n_522), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_652), .B(n_21), .Y(n_773) );
O2A1O1Ixp33_ASAP7_75t_SL g774 ( .A1(n_714), .A2(n_124), .B(n_125), .C(n_119), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_670), .B(n_22), .Y(n_775) );
A2O1A1Ixp33_ASAP7_75t_L g776 ( .A1(n_676), .A2(n_522), .B(n_561), .C(n_556), .Y(n_776) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_717), .A2(n_129), .B(n_128), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g778 ( .A(n_685), .B(n_551), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_648), .Y(n_779) );
CKINVDCx11_ASAP7_75t_R g780 ( .A(n_642), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_741), .A2(n_556), .B(n_551), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_643), .B(n_23), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_SL g783 ( .A1(n_701), .A2(n_132), .B(n_134), .C(n_130), .Y(n_783) );
A2O1A1Ixp33_ASAP7_75t_L g784 ( .A1(n_716), .A2(n_556), .B(n_561), .C(n_551), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_744), .B(n_25), .Y(n_785) );
OAI21x1_ASAP7_75t_L g786 ( .A1(n_728), .A2(n_136), .B(n_135), .Y(n_786) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_706), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_666), .A2(n_138), .B(n_137), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_650), .A2(n_28), .B1(n_26), .B2(n_27), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_715), .A2(n_561), .B(n_144), .Y(n_790) );
INVx1_ASAP7_75t_SL g791 ( .A(n_742), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_688), .A2(n_150), .B(n_142), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_693), .A2(n_154), .B(n_152), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_SL g794 ( .A1(n_722), .A2(n_185), .B(n_314), .C(n_313), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_650), .A2(n_29), .B1(n_31), .B2(n_32), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g796 ( .A1(n_696), .A2(n_158), .B(n_155), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_671), .B(n_31), .Y(n_797) );
AO32x2_ASAP7_75t_L g798 ( .A1(n_702), .A2(n_32), .A3(n_33), .B1(n_34), .B2(n_35), .Y(n_798) );
AO31x2_ASAP7_75t_L g799 ( .A1(n_709), .A2(n_35), .A3(n_36), .B(n_37), .Y(n_799) );
AOI221x1_ASAP7_75t_L g800 ( .A1(n_681), .A2(n_38), .B1(n_41), .B2(n_42), .C(n_43), .Y(n_800) );
INVx3_ASAP7_75t_L g801 ( .A(n_687), .Y(n_801) );
NAND2xp5_ASAP7_75t_SL g802 ( .A(n_687), .B(n_44), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_718), .A2(n_162), .B(n_161), .Y(n_803) );
AO21x2_ASAP7_75t_L g804 ( .A1(n_682), .A2(n_167), .B(n_165), .Y(n_804) );
AND2x4_ASAP7_75t_L g805 ( .A(n_710), .B(n_45), .Y(n_805) );
A2O1A1Ixp33_ASAP7_75t_L g806 ( .A1(n_686), .A2(n_45), .B(n_46), .C(n_47), .Y(n_806) );
A2O1A1Ixp33_ASAP7_75t_L g807 ( .A1(n_689), .A2(n_46), .B(n_48), .C(n_49), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_669), .B(n_48), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_713), .A2(n_169), .B(n_168), .Y(n_809) );
A2O1A1Ixp33_ASAP7_75t_L g810 ( .A1(n_695), .A2(n_49), .B(n_50), .C(n_52), .Y(n_810) );
AOI21x1_ASAP7_75t_L g811 ( .A1(n_721), .A2(n_173), .B(n_170), .Y(n_811) );
O2A1O1Ixp33_ASAP7_75t_SL g812 ( .A1(n_720), .A2(n_207), .B(n_312), .C(n_308), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_703), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_813) );
BUFx3_ASAP7_75t_L g814 ( .A(n_708), .Y(n_814) );
INVx8_ASAP7_75t_L g815 ( .A(n_662), .Y(n_815) );
AO31x2_ASAP7_75t_L g816 ( .A1(n_709), .A2(n_54), .A3(n_55), .B(n_56), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_653), .A2(n_57), .B1(n_58), .B2(n_59), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_694), .Y(n_818) );
OAI21x1_ASAP7_75t_L g819 ( .A1(n_698), .A2(n_178), .B(n_177), .Y(n_819) );
BUFx12f_ASAP7_75t_L g820 ( .A(n_662), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_712), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_821) );
O2A1O1Ixp33_ASAP7_75t_SL g822 ( .A1(n_745), .A2(n_217), .B(n_307), .C(n_306), .Y(n_822) );
INVx3_ASAP7_75t_SL g823 ( .A(n_653), .Y(n_823) );
INVxp67_ASAP7_75t_SL g824 ( .A(n_746), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_684), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_707), .B(n_64), .Y(n_826) );
OAI21xp5_ASAP7_75t_L g827 ( .A1(n_719), .A2(n_181), .B(n_180), .Y(n_827) );
O2A1O1Ixp33_ASAP7_75t_L g828 ( .A1(n_656), .A2(n_64), .B(n_65), .C(n_66), .Y(n_828) );
AO31x2_ASAP7_75t_L g829 ( .A1(n_730), .A2(n_65), .A3(n_66), .B(n_69), .Y(n_829) );
OAI21x1_ASAP7_75t_L g830 ( .A1(n_700), .A2(n_186), .B(n_182), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_683), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_690), .A2(n_69), .B1(n_71), .B2(n_73), .Y(n_832) );
OAI221xp5_ASAP7_75t_SL g833 ( .A1(n_699), .A2(n_73), .B1(n_74), .B2(n_75), .C(n_76), .Y(n_833) );
AO31x2_ASAP7_75t_L g834 ( .A1(n_704), .A2(n_77), .A3(n_78), .B(n_80), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_677), .B(n_77), .Y(n_835) );
OAI21xp5_ASAP7_75t_L g836 ( .A1(n_667), .A2(n_229), .B(n_304), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_680), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_664), .B(n_78), .Y(n_838) );
AND2x4_ASAP7_75t_L g839 ( .A(n_672), .B(n_81), .Y(n_839) );
O2A1O1Ixp33_ASAP7_75t_L g840 ( .A1(n_645), .A2(n_82), .B(n_85), .C(n_87), .Y(n_840) );
AOI221xp5_ASAP7_75t_L g841 ( .A1(n_660), .A2(n_85), .B1(n_87), .B2(n_88), .C(n_89), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_651), .B(n_88), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_705), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_735), .Y(n_844) );
AOI21xp5_ASAP7_75t_L g845 ( .A1(n_723), .A2(n_238), .B(n_302), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_737), .Y(n_846) );
OAI21x1_ASAP7_75t_L g847 ( .A1(n_738), .A2(n_235), .B(n_300), .Y(n_847) );
A2O1A1Ixp33_ASAP7_75t_L g848 ( .A1(n_732), .A2(n_89), .B(n_90), .C(n_91), .Y(n_848) );
OAI21xp5_ASAP7_75t_L g849 ( .A1(n_743), .A2(n_239), .B(n_298), .Y(n_849) );
AND2x4_ASAP7_75t_L g850 ( .A(n_661), .B(n_92), .Y(n_850) );
OA21x2_ASAP7_75t_L g851 ( .A1(n_723), .A2(n_241), .B(n_296), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_725), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_723), .A2(n_240), .B(n_295), .Y(n_853) );
O2A1O1Ixp33_ASAP7_75t_SL g854 ( .A1(n_726), .A2(n_234), .B(n_294), .C(n_293), .Y(n_854) );
A2O1A1Ixp33_ASAP7_75t_L g855 ( .A1(n_724), .A2(n_93), .B(n_94), .C(n_95), .Y(n_855) );
INVx2_ASAP7_75t_SL g856 ( .A(n_729), .Y(n_856) );
NAND2xp5_ASAP7_75t_SL g857 ( .A(n_711), .B(n_93), .Y(n_857) );
AO32x2_ASAP7_75t_L g858 ( .A1(n_725), .A2(n_94), .A3(n_95), .B1(n_96), .B2(n_97), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_725), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g860 ( .A1(n_727), .A2(n_231), .B(n_291), .Y(n_860) );
AO32x2_ASAP7_75t_L g861 ( .A1(n_711), .A2(n_96), .A3(n_97), .B1(n_98), .B2(n_99), .Y(n_861) );
A2O1A1Ixp33_ASAP7_75t_L g862 ( .A1(n_734), .A2(n_99), .B(n_100), .C(n_101), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_692), .A2(n_247), .B(n_290), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_736), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_864) );
INVx1_ASAP7_75t_SL g865 ( .A(n_791), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_755), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_760), .Y(n_867) );
INVx4_ASAP7_75t_L g868 ( .A(n_768), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_779), .B(n_106), .Y(n_869) );
AND2x4_ASAP7_75t_L g870 ( .A(n_801), .B(n_107), .Y(n_870) );
INVx6_ASAP7_75t_L g871 ( .A(n_820), .Y(n_871) );
AO22x1_ASAP7_75t_L g872 ( .A1(n_805), .A2(n_108), .B1(n_109), .B2(n_111), .Y(n_872) );
AO31x2_ASAP7_75t_L g873 ( .A1(n_761), .A2(n_109), .A3(n_111), .B(n_187), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_763), .B(n_192), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_753), .Y(n_875) );
OR2x2_ASAP7_75t_L g876 ( .A(n_808), .B(n_195), .Y(n_876) );
BUFx6f_ASAP7_75t_L g877 ( .A(n_750), .Y(n_877) );
OAI22xp33_ASAP7_75t_L g878 ( .A1(n_768), .A2(n_196), .B1(n_198), .B2(n_203), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_770), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_782), .B(n_205), .Y(n_880) );
OAI21xp33_ASAP7_75t_L g881 ( .A1(n_864), .A2(n_208), .B(n_210), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_770), .A2(n_211), .B1(n_212), .B2(n_216), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_773), .B(n_220), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_850), .A2(n_221), .B1(n_223), .B2(n_224), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_775), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_850), .A2(n_227), .B1(n_228), .B2(n_243), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_823), .A2(n_244), .B1(n_245), .B2(n_248), .Y(n_887) );
AOI21x1_ASAP7_75t_L g888 ( .A1(n_852), .A2(n_250), .B(n_252), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_815), .B(n_253), .Y(n_889) );
NAND3xp33_ASAP7_75t_L g890 ( .A(n_800), .B(n_254), .C(n_255), .Y(n_890) );
AOI21xp33_ASAP7_75t_L g891 ( .A1(n_828), .A2(n_257), .B(n_258), .Y(n_891) );
BUFx3_ASAP7_75t_L g892 ( .A(n_767), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_749), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_773), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_831), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_789), .Y(n_896) );
BUFx4f_ASAP7_75t_SL g897 ( .A(n_814), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_825), .B(n_263), .Y(n_898) );
BUFx3_ASAP7_75t_L g899 ( .A(n_780), .Y(n_899) );
A2O1A1Ixp33_ASAP7_75t_L g900 ( .A1(n_766), .A2(n_265), .B(n_268), .C(n_269), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_758), .B(n_284), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_844), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_815), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_785), .B(n_270), .Y(n_904) );
INVx3_ASAP7_75t_L g905 ( .A(n_801), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_837), .B(n_283), .Y(n_906) );
OA21x2_ASAP7_75t_L g907 ( .A1(n_859), .A2(n_276), .B(n_277), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_846), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_795), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_843), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_826), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_799), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_799), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_799), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_818), .B(n_839), .Y(n_915) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_856), .Y(n_916) );
AOI22xp5_ASAP7_75t_L g917 ( .A1(n_813), .A2(n_821), .B1(n_817), .B2(n_835), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g918 ( .A1(n_759), .A2(n_748), .B(n_757), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_816), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_802), .A2(n_797), .B1(n_838), .B2(n_842), .Y(n_920) );
AO31x2_ASAP7_75t_L g921 ( .A1(n_784), .A2(n_776), .A3(n_751), .B(n_756), .Y(n_921) );
CKINVDCx16_ASAP7_75t_R g922 ( .A(n_772), .Y(n_922) );
A2O1A1Ixp33_ASAP7_75t_L g923 ( .A1(n_840), .A2(n_862), .B(n_807), .C(n_810), .Y(n_923) );
INVx4_ASAP7_75t_L g924 ( .A(n_750), .Y(n_924) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_833), .B(n_857), .Y(n_925) );
AO31x2_ASAP7_75t_L g926 ( .A1(n_845), .A2(n_853), .A3(n_863), .B(n_765), .Y(n_926) );
INVx3_ASAP7_75t_L g927 ( .A(n_750), .Y(n_927) );
O2A1O1Ixp33_ASAP7_75t_L g928 ( .A1(n_806), .A2(n_832), .B(n_848), .C(n_855), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_816), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_841), .A2(n_754), .B1(n_836), .B2(n_827), .Y(n_930) );
AOI21xp5_ASAP7_75t_L g931 ( .A1(n_769), .A2(n_774), .B(n_752), .Y(n_931) );
AOI22xp33_ASAP7_75t_SL g932 ( .A1(n_788), .A2(n_777), .B1(n_849), .B2(n_804), .Y(n_932) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_778), .B(n_824), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_798), .Y(n_934) );
OR2x6_ASAP7_75t_L g935 ( .A(n_764), .B(n_787), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_798), .Y(n_936) );
OA21x2_ASAP7_75t_L g937 ( .A1(n_819), .A2(n_830), .B(n_786), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_798), .Y(n_938) );
AOI21x1_ASAP7_75t_L g939 ( .A1(n_811), .A2(n_851), .B(n_790), .Y(n_939) );
OAI21xp5_ASAP7_75t_L g940 ( .A1(n_803), .A2(n_793), .B(n_792), .Y(n_940) );
AOI21xp33_ASAP7_75t_L g941 ( .A1(n_847), .A2(n_796), .B(n_764), .Y(n_941) );
OA21x2_ASAP7_75t_L g942 ( .A1(n_860), .A2(n_809), .B(n_822), .Y(n_942) );
AND2x4_ASAP7_75t_L g943 ( .A(n_787), .B(n_762), .Y(n_943) );
OAI21xp5_ASAP7_75t_L g944 ( .A1(n_794), .A2(n_783), .B(n_854), .Y(n_944) );
AOI21xp5_ASAP7_75t_L g945 ( .A1(n_812), .A2(n_762), .B(n_858), .Y(n_945) );
AOI21xp5_ASAP7_75t_L g946 ( .A1(n_762), .A2(n_858), .B(n_834), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_861), .B(n_834), .Y(n_947) );
AOI21xp5_ASAP7_75t_L g948 ( .A1(n_829), .A2(n_610), .B(n_771), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_829), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_829), .Y(n_950) );
AOI21xp33_ASAP7_75t_L g951 ( .A1(n_861), .A2(n_782), .B(n_828), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_791), .B(n_733), .Y(n_952) );
A2O1A1Ixp33_ASAP7_75t_L g953 ( .A1(n_779), .A2(n_658), .B(n_734), .C(n_782), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_779), .B(n_733), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_779), .B(n_733), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_771), .A2(n_610), .B(n_781), .Y(n_956) );
AND2x4_ASAP7_75t_L g957 ( .A(n_779), .B(n_658), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_779), .B(n_733), .Y(n_958) );
AOI21xp5_ASAP7_75t_L g959 ( .A1(n_771), .A2(n_610), .B(n_781), .Y(n_959) );
OR2x2_ASAP7_75t_L g960 ( .A(n_791), .B(n_733), .Y(n_960) );
AO31x2_ASAP7_75t_L g961 ( .A1(n_761), .A2(n_852), .A3(n_859), .B(n_784), .Y(n_961) );
BUFx6f_ASAP7_75t_L g962 ( .A(n_750), .Y(n_962) );
NAND2xp5_ASAP7_75t_SL g963 ( .A(n_753), .B(n_733), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_773), .B(n_733), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_773), .B(n_733), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_755), .Y(n_966) );
A2O1A1Ixp33_ASAP7_75t_L g967 ( .A1(n_779), .A2(n_658), .B(n_734), .C(n_782), .Y(n_967) );
OAI21xp5_ASAP7_75t_L g968 ( .A1(n_837), .A2(n_692), .B(n_641), .Y(n_968) );
BUFx3_ASAP7_75t_L g969 ( .A(n_767), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_773), .B(n_733), .Y(n_970) );
OAI21xp5_ASAP7_75t_L g971 ( .A1(n_837), .A2(n_692), .B(n_641), .Y(n_971) );
NAND2x1_ASAP7_75t_L g972 ( .A(n_768), .B(n_801), .Y(n_972) );
INVx2_ASAP7_75t_SL g973 ( .A(n_791), .Y(n_973) );
NAND2xp5_ASAP7_75t_SL g974 ( .A(n_753), .B(n_733), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g975 ( .A1(n_763), .A2(n_668), .B1(n_579), .B2(n_675), .C(n_578), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_755), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_943), .Y(n_977) );
INVx1_ASAP7_75t_SL g978 ( .A(n_897), .Y(n_978) );
HB1xp67_ASAP7_75t_L g979 ( .A(n_957), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_867), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_943), .Y(n_981) );
AND2x4_ASAP7_75t_L g982 ( .A(n_935), .B(n_924), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_964), .B(n_965), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_970), .B(n_954), .Y(n_984) );
OR2x2_ASAP7_75t_L g985 ( .A(n_952), .B(n_960), .Y(n_985) );
BUFx3_ASAP7_75t_L g986 ( .A(n_903), .Y(n_986) );
INVx2_ASAP7_75t_L g987 ( .A(n_875), .Y(n_987) );
AND2x4_ASAP7_75t_L g988 ( .A(n_935), .B(n_924), .Y(n_988) );
AO21x2_ASAP7_75t_L g989 ( .A1(n_931), .A2(n_948), .B(n_945), .Y(n_989) );
AND2x4_ASAP7_75t_L g990 ( .A(n_935), .B(n_927), .Y(n_990) );
INVxp67_ASAP7_75t_L g991 ( .A(n_916), .Y(n_991) );
INVx2_ASAP7_75t_SL g992 ( .A(n_972), .Y(n_992) );
OR2x2_ASAP7_75t_L g993 ( .A(n_955), .B(n_958), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_966), .B(n_976), .Y(n_994) );
INVx3_ASAP7_75t_L g995 ( .A(n_877), .Y(n_995) );
OA21x2_ASAP7_75t_L g996 ( .A1(n_946), .A2(n_956), .B(n_959), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_910), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_870), .Y(n_998) );
OAI21xp5_ASAP7_75t_L g999 ( .A1(n_923), .A2(n_928), .B(n_925), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_869), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_895), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_902), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_896), .B(n_909), .Y(n_1003) );
INVx1_ASAP7_75t_SL g1004 ( .A(n_865), .Y(n_1004) );
OR2x2_ASAP7_75t_L g1005 ( .A(n_865), .B(n_973), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_908), .Y(n_1006) );
BUFx3_ASAP7_75t_L g1007 ( .A(n_892), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_885), .B(n_947), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_894), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_911), .B(n_893), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_879), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1012 ( .A(n_868), .B(n_915), .Y(n_1012) );
AOI21xp5_ASAP7_75t_SL g1013 ( .A1(n_884), .A2(n_886), .B(n_882), .Y(n_1013) );
AOI33xp33_ASAP7_75t_L g1014 ( .A1(n_949), .A2(n_950), .A3(n_929), .B1(n_913), .B2(n_914), .B3(n_919), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_874), .B(n_876), .Y(n_1015) );
OR2x6_ASAP7_75t_L g1016 ( .A(n_884), .B(n_886), .Y(n_1016) );
OR2x6_ASAP7_75t_L g1017 ( .A(n_883), .B(n_882), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_963), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_974), .Y(n_1019) );
AND2x4_ASAP7_75t_L g1020 ( .A(n_927), .B(n_905), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_877), .Y(n_1021) );
AOI21xp5_ASAP7_75t_SL g1022 ( .A1(n_930), .A2(n_878), .B(n_881), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_872), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_912), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_917), .B(n_922), .Y(n_1025) );
BUFx3_ASAP7_75t_L g1026 ( .A(n_969), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_934), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_905), .B(n_889), .Y(n_1028) );
AOI21xp5_ASAP7_75t_L g1029 ( .A1(n_944), .A2(n_918), .B(n_940), .Y(n_1029) );
INVx2_ASAP7_75t_L g1030 ( .A(n_961), .Y(n_1030) );
AO21x2_ASAP7_75t_L g1031 ( .A1(n_951), .A2(n_944), .B(n_939), .Y(n_1031) );
OAI21xp5_ASAP7_75t_L g1032 ( .A1(n_890), .A2(n_951), .B(n_920), .Y(n_1032) );
OR2x6_ASAP7_75t_L g1033 ( .A(n_871), .B(n_899), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_936), .B(n_938), .Y(n_1034) );
OR2x2_ASAP7_75t_L g1035 ( .A(n_904), .B(n_906), .Y(n_1035) );
INVx3_ASAP7_75t_L g1036 ( .A(n_962), .Y(n_1036) );
HB1xp67_ASAP7_75t_L g1037 ( .A(n_962), .Y(n_1037) );
AO21x2_ASAP7_75t_L g1038 ( .A1(n_891), .A2(n_968), .B(n_971), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_873), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_871), .Y(n_1040) );
INVxp67_ASAP7_75t_L g1041 ( .A(n_933), .Y(n_1041) );
AND2x4_ASAP7_75t_L g1042 ( .A(n_962), .B(n_971), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_968), .B(n_873), .Y(n_1043) );
NOR2xp33_ASAP7_75t_L g1044 ( .A(n_880), .B(n_901), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_898), .B(n_873), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_907), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_900), .B(n_891), .Y(n_1047) );
OA21x2_ASAP7_75t_L g1048 ( .A1(n_940), .A2(n_888), .B(n_941), .Y(n_1048) );
INVx3_ASAP7_75t_L g1049 ( .A(n_921), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_887), .B(n_921), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_907), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1052 ( .A(n_921), .Y(n_1052) );
INVx2_ASAP7_75t_L g1053 ( .A(n_937), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_926), .B(n_932), .Y(n_1054) );
OR2x6_ASAP7_75t_L g1055 ( .A(n_942), .B(n_972), .Y(n_1055) );
AO21x2_ASAP7_75t_L g1056 ( .A1(n_931), .A2(n_948), .B(n_945), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_866), .Y(n_1057) );
INVx2_ASAP7_75t_L g1058 ( .A(n_943), .Y(n_1058) );
AO21x2_ASAP7_75t_L g1059 ( .A1(n_931), .A2(n_948), .B(n_945), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_896), .A2(n_909), .B1(n_649), .B2(n_736), .Y(n_1060) );
AND2x4_ASAP7_75t_L g1061 ( .A(n_957), .B(n_935), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_868), .A2(n_590), .B1(n_768), .B2(n_649), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_866), .Y(n_1063) );
OAI21xp5_ASAP7_75t_L g1064 ( .A1(n_953), .A2(n_967), .B(n_923), .Y(n_1064) );
INVxp67_ASAP7_75t_SL g1065 ( .A(n_957), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_943), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_866), .Y(n_1067) );
AO21x2_ASAP7_75t_L g1068 ( .A1(n_931), .A2(n_948), .B(n_945), .Y(n_1068) );
AO21x2_ASAP7_75t_L g1069 ( .A1(n_931), .A2(n_948), .B(n_945), .Y(n_1069) );
INVx2_ASAP7_75t_SL g1070 ( .A(n_897), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_866), .Y(n_1071) );
INVx1_ASAP7_75t_SL g1072 ( .A(n_897), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_975), .B(n_733), .Y(n_1073) );
AOI21xp5_ASAP7_75t_R g1074 ( .A1(n_1062), .A2(n_1061), .B(n_988), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1053), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1008), .B(n_1034), .Y(n_1076) );
NOR2x1_ASAP7_75t_SL g1077 ( .A(n_1016), .B(n_1017), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1010), .B(n_984), .Y(n_1078) );
OR2x2_ASAP7_75t_L g1079 ( .A(n_1008), .B(n_1025), .Y(n_1079) );
BUFx2_ASAP7_75t_L g1080 ( .A(n_1016), .Y(n_1080) );
INVx4_ASAP7_75t_L g1081 ( .A(n_1016), .Y(n_1081) );
OR2x2_ASAP7_75t_L g1082 ( .A(n_979), .B(n_1003), .Y(n_1082) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_982), .Y(n_1083) );
OR2x6_ASAP7_75t_L g1084 ( .A(n_1013), .B(n_1017), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1034), .B(n_1043), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1043), .B(n_977), .Y(n_1086) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_979), .B(n_1024), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_977), .B(n_981), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1089 ( .A(n_985), .B(n_1065), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1014), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g1091 ( .A(n_1004), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_981), .B(n_1058), .Y(n_1092) );
BUFx2_ASAP7_75t_SL g1093 ( .A(n_992), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g1094 ( .A(n_1005), .Y(n_1094) );
AO21x2_ASAP7_75t_L g1095 ( .A1(n_1029), .A2(n_1032), .B(n_1051), .Y(n_1095) );
INVx2_ASAP7_75t_SL g1096 ( .A(n_982), .Y(n_1096) );
AOI22xp33_ASAP7_75t_SL g1097 ( .A1(n_1023), .A2(n_992), .B1(n_998), .B2(n_1061), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_980), .Y(n_1098) );
AOI221xp5_ASAP7_75t_L g1099 ( .A1(n_999), .A2(n_1064), .B1(n_1073), .B2(n_1000), .C(n_991), .Y(n_1099) );
AND2x4_ASAP7_75t_SL g1100 ( .A(n_1033), .B(n_1061), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1066), .B(n_983), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1027), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1039), .Y(n_1103) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_1060), .A2(n_1015), .B1(n_1044), .B2(n_1041), .C(n_1012), .Y(n_1104) );
INVxp67_ASAP7_75t_L g1105 ( .A(n_1007), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1054), .B(n_987), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_1044), .A2(n_1060), .B1(n_1035), .B2(n_1033), .Y(n_1107) );
AO22x1_ASAP7_75t_L g1108 ( .A1(n_982), .A2(n_988), .B1(n_990), .B2(n_1026), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1057), .Y(n_1109) );
INVx3_ASAP7_75t_L g1110 ( .A(n_1042), .Y(n_1110) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_997), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1030), .Y(n_1112) );
AND2x4_ASAP7_75t_L g1113 ( .A(n_1055), .B(n_988), .Y(n_1113) );
INVx5_ASAP7_75t_L g1114 ( .A(n_995), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_993), .B(n_1067), .Y(n_1115) );
AND2x4_ASAP7_75t_L g1116 ( .A(n_1055), .B(n_1049), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1063), .B(n_1071), .Y(n_1117) );
BUFx3_ASAP7_75t_L g1118 ( .A(n_1026), .Y(n_1118) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_1001), .Y(n_1119) );
OAI211xp5_ASAP7_75t_L g1120 ( .A1(n_1022), .A2(n_1040), .B(n_1028), .C(n_1019), .Y(n_1120) );
INVx1_ASAP7_75t_SL g1121 ( .A(n_986), .Y(n_1121) );
AND2x2_ASAP7_75t_SL g1122 ( .A(n_1050), .B(n_1022), .Y(n_1122) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_994), .B(n_1052), .Y(n_1123) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1075), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1103), .Y(n_1125) );
AOI221xp5_ASAP7_75t_L g1126 ( .A1(n_1099), .A2(n_1011), .B1(n_1009), .B2(n_1018), .C(n_1006), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1103), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1085), .B(n_1049), .Y(n_1128) );
NAND3xp33_ASAP7_75t_SL g1129 ( .A(n_1121), .B(n_978), .C(n_1072), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1076), .B(n_1002), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1102), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1085), .B(n_1049), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1076), .B(n_1020), .Y(n_1133) );
OR2x2_ASAP7_75t_L g1134 ( .A(n_1079), .B(n_996), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1102), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1086), .B(n_1031), .Y(n_1136) );
INVx6_ASAP7_75t_L g1137 ( .A(n_1118), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1086), .B(n_1031), .Y(n_1138) );
BUFx2_ASAP7_75t_L g1139 ( .A(n_1084), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1106), .B(n_1038), .Y(n_1140) );
INVx3_ASAP7_75t_L g1141 ( .A(n_1116), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1106), .B(n_1038), .Y(n_1142) );
NAND2xp33_ASAP7_75t_SL g1143 ( .A(n_1081), .B(n_1070), .Y(n_1143) );
HB1xp67_ASAP7_75t_L g1144 ( .A(n_1119), .Y(n_1144) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_1079), .B(n_1056), .Y(n_1145) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_1104), .A2(n_1070), .B1(n_986), .B2(n_1020), .C(n_1047), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1084), .B(n_989), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1112), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1084), .B(n_989), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1084), .B(n_1069), .Y(n_1150) );
HB1xp67_ASAP7_75t_L g1151 ( .A(n_1111), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1088), .B(n_1069), .Y(n_1152) );
INVx3_ASAP7_75t_L g1153 ( .A(n_1113), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1088), .B(n_1068), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1092), .B(n_1068), .Y(n_1155) );
OR2x2_ASAP7_75t_L g1156 ( .A(n_1123), .B(n_1059), .Y(n_1156) );
INVx4_ASAP7_75t_L g1157 ( .A(n_1114), .Y(n_1157) );
AND2x4_ASAP7_75t_L g1158 ( .A(n_1077), .B(n_1056), .Y(n_1158) );
INVx6_ASAP7_75t_L g1159 ( .A(n_1118), .Y(n_1159) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1123), .B(n_1045), .Y(n_1160) );
AND2x4_ASAP7_75t_L g1161 ( .A(n_1077), .B(n_1046), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1087), .B(n_1037), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1101), .B(n_990), .Y(n_1163) );
HB1xp67_ASAP7_75t_L g1164 ( .A(n_1091), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1087), .B(n_1021), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1080), .B(n_1048), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1131), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1145), .B(n_1094), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1131), .Y(n_1169) );
NAND4xp75_ASAP7_75t_L g1170 ( .A(n_1146), .B(n_1107), .C(n_1122), .D(n_1074), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1128), .B(n_1080), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1124), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1132), .B(n_1081), .Y(n_1173) );
NAND2xp5_ASAP7_75t_SL g1174 ( .A(n_1143), .B(n_1105), .Y(n_1174) );
INVx2_ASAP7_75t_SL g1175 ( .A(n_1137), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1145), .B(n_1082), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1135), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1135), .Y(n_1178) );
INVx2_ASAP7_75t_L g1179 ( .A(n_1124), .Y(n_1179) );
AND2x2_ASAP7_75t_SL g1180 ( .A(n_1139), .B(n_1122), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1136), .B(n_1138), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1125), .Y(n_1182) );
NOR2x1_ASAP7_75t_L g1183 ( .A(n_1129), .B(n_1093), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1125), .Y(n_1184) );
INVxp67_ASAP7_75t_L g1185 ( .A(n_1144), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1127), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1134), .B(n_1090), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1188 ( .A(n_1151), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1134), .B(n_1109), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1152), .B(n_1110), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1148), .Y(n_1191) );
NOR2x1_ASAP7_75t_R g1192 ( .A(n_1157), .B(n_1093), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1140), .B(n_1098), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1154), .B(n_1110), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1140), .B(n_1095), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1154), .B(n_1095), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1181), .B(n_1142), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1167), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1167), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1181), .B(n_1160), .Y(n_1200) );
AND2x6_ASAP7_75t_L g1201 ( .A(n_1192), .B(n_1161), .Y(n_1201) );
BUFx2_ASAP7_75t_L g1202 ( .A(n_1192), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1169), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1172), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1169), .Y(n_1205) );
INVxp67_ASAP7_75t_L g1206 ( .A(n_1188), .Y(n_1206) );
INVx2_ASAP7_75t_L g1207 ( .A(n_1172), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1187), .B(n_1164), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1189), .Y(n_1209) );
OAI32xp33_ASAP7_75t_L g1210 ( .A1(n_1174), .A2(n_1157), .A3(n_1130), .B1(n_1133), .B2(n_1165), .Y(n_1210) );
AOI21xp33_ASAP7_75t_SL g1211 ( .A1(n_1180), .A2(n_1108), .B(n_1158), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1189), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1190), .B(n_1166), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1168), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1168), .Y(n_1215) );
NAND3xp33_ASAP7_75t_L g1216 ( .A(n_1183), .B(n_1126), .C(n_1120), .Y(n_1216) );
OAI32xp33_ASAP7_75t_L g1217 ( .A1(n_1185), .A2(n_1165), .A3(n_1162), .B1(n_1153), .B2(n_1078), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1177), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1187), .B(n_1155), .Y(n_1219) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1179), .Y(n_1220) );
INVxp67_ASAP7_75t_L g1221 ( .A(n_1208), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1197), .B(n_1196), .Y(n_1222) );
NAND3x2_ASAP7_75t_L g1223 ( .A(n_1202), .B(n_1139), .C(n_1176), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1224 ( .A(n_1200), .B(n_1195), .Y(n_1224) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1204), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1209), .B(n_1196), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1212), .B(n_1193), .Y(n_1227) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1204), .Y(n_1228) );
INVxp67_ASAP7_75t_SL g1229 ( .A(n_1206), .Y(n_1229) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_1216), .A2(n_1170), .B1(n_1171), .B2(n_1173), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1214), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1215), .Y(n_1232) );
NOR3xp33_ASAP7_75t_L g1233 ( .A(n_1210), .B(n_1097), .C(n_1175), .Y(n_1233) );
AOI221x1_ASAP7_75t_L g1234 ( .A1(n_1211), .A2(n_1117), .B1(n_1158), .B2(n_1115), .C(n_1191), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1222), .B(n_1213), .Y(n_1235) );
O2A1O1Ixp33_ASAP7_75t_L g1236 ( .A1(n_1229), .A2(n_1217), .B(n_1219), .C(n_1203), .Y(n_1236) );
AOI221x1_ASAP7_75t_L g1237 ( .A1(n_1233), .A2(n_1203), .B1(n_1218), .B2(n_1198), .C(n_1199), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1222), .B(n_1194), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1229), .Y(n_1239) );
AOI211xp5_ASAP7_75t_SL g1240 ( .A1(n_1230), .A2(n_1201), .B(n_1150), .C(n_1147), .Y(n_1240) );
OAI21xp5_ASAP7_75t_L g1241 ( .A1(n_1223), .A2(n_1201), .B(n_1149), .Y(n_1241) );
NOR2xp33_ASAP7_75t_L g1242 ( .A(n_1221), .B(n_1205), .Y(n_1242) );
OAI21xp5_ASAP7_75t_L g1243 ( .A1(n_1234), .A2(n_1201), .B(n_1161), .Y(n_1243) );
AOI221xp5_ASAP7_75t_L g1244 ( .A1(n_1236), .A2(n_1232), .B1(n_1231), .B2(n_1227), .C(n_1226), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1239), .Y(n_1245) );
OAI211xp5_ASAP7_75t_SL g1246 ( .A1(n_1240), .A2(n_1224), .B(n_1089), .C(n_1141), .Y(n_1246) );
OAI21xp33_ASAP7_75t_SL g1247 ( .A1(n_1243), .A2(n_1228), .B(n_1225), .Y(n_1247) );
BUFx2_ASAP7_75t_L g1248 ( .A(n_1241), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1242), .Y(n_1249) );
OR3x1_ASAP7_75t_L g1250 ( .A(n_1246), .B(n_1237), .C(n_1182), .Y(n_1250) );
INVxp67_ASAP7_75t_L g1251 ( .A(n_1245), .Y(n_1251) );
NAND3xp33_ASAP7_75t_L g1252 ( .A(n_1244), .B(n_1235), .C(n_1238), .Y(n_1252) );
INVxp67_ASAP7_75t_L g1253 ( .A(n_1249), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1248), .B(n_1235), .Y(n_1254) );
NOR2xp33_ASAP7_75t_L g1255 ( .A(n_1247), .B(n_1238), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1249), .B(n_1178), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1254), .B(n_1156), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1255), .B(n_1141), .Y(n_1258) );
OAI211xp5_ASAP7_75t_SL g1259 ( .A1(n_1253), .A2(n_1162), .B(n_1163), .C(n_1083), .Y(n_1259) );
INVx1_ASAP7_75t_SL g1260 ( .A(n_1256), .Y(n_1260) );
INVx2_ASAP7_75t_SL g1261 ( .A(n_1252), .Y(n_1261) );
AO21x2_ASAP7_75t_L g1262 ( .A1(n_1258), .A2(n_1251), .B(n_1250), .Y(n_1262) );
INVx1_ASAP7_75t_SL g1263 ( .A(n_1260), .Y(n_1263) );
OR5x1_ASAP7_75t_L g1264 ( .A(n_1261), .B(n_1100), .C(n_1159), .D(n_1137), .E(n_1096), .Y(n_1264) );
AND2x4_ASAP7_75t_L g1265 ( .A(n_1257), .B(n_1100), .Y(n_1265) );
OAI22xp5_ASAP7_75t_SL g1266 ( .A1(n_1263), .A2(n_1159), .B1(n_1259), .B2(n_1096), .Y(n_1266) );
HB1xp67_ASAP7_75t_L g1267 ( .A(n_1262), .Y(n_1267) );
XNOR2xp5_ASAP7_75t_L g1268 ( .A(n_1264), .B(n_1083), .Y(n_1268) );
OAI22xp5_ASAP7_75t_SL g1269 ( .A1(n_1267), .A2(n_1265), .B1(n_1159), .B2(n_1161), .Y(n_1269) );
AOI21xp5_ASAP7_75t_L g1270 ( .A1(n_1269), .A2(n_1268), .B(n_1266), .Y(n_1270) );
OA21x2_ASAP7_75t_L g1271 ( .A1(n_1270), .A2(n_1186), .B(n_1184), .Y(n_1271) );
OAI21xp5_ASAP7_75t_L g1272 ( .A1(n_1271), .A2(n_1114), .B(n_1036), .Y(n_1272) );
AOI21xp5_ASAP7_75t_L g1273 ( .A1(n_1272), .A2(n_1220), .B(n_1207), .Y(n_1273) );
endmodule