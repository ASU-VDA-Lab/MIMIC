module fake_jpeg_4973_n_240 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_240);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_240;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_114;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

CKINVDCx9p33_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_31),
.B1(n_22),
.B2(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_32),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_46),
.B(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_24),
.B(n_0),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_31),
.B1(n_30),
.B2(n_23),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_75),
.B1(n_5),
.B2(n_7),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_60),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_31),
.B1(n_27),
.B2(n_30),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_64),
.B1(n_79),
.B2(n_2),
.Y(n_91)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_65),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_33),
.A2(n_15),
.B1(n_23),
.B2(n_21),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_15),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_77),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_36),
.A2(n_25),
.B1(n_20),
.B2(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_39),
.A2(n_26),
.B1(n_20),
.B2(n_19),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_37),
.A2(n_26),
.B(n_16),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_4),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_16),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_37),
.B(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_3),
.Y(n_100)
);

OR2x4_ASAP7_75t_SL g87 ( 
.A(n_38),
.B(n_2),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_3),
.B(n_4),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_91),
.A2(n_95),
.B1(n_108),
.B2(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_66),
.B1(n_74),
.B2(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_53),
.B1(n_52),
.B2(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_8),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_101),
.A2(n_10),
.B(n_54),
.C(n_78),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_10),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_12),
.C(n_14),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_5),
.C(n_8),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_5),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_72),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_129),
.B1(n_115),
.B2(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_122),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_124),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_87),
.B(n_76),
.C(n_66),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_127),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_77),
.B1(n_76),
.B2(n_67),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_76),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_143),
.B(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_142),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_65),
.B1(n_78),
.B2(n_76),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_117),
.B1(n_62),
.B2(n_67),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_49),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_10),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_54),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_100),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_72),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_144),
.B(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_154),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_130),
.B1(n_133),
.B2(n_144),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_95),
.B(n_99),
.C(n_83),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_160),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_168),
.B(n_130),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_110),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_106),
.C(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_131),
.B1(n_62),
.B2(n_83),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_125),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_129),
.B(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_122),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_181),
.B1(n_185),
.B2(n_186),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_90),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_180),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_174),
.B1(n_172),
.B2(n_188),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_93),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_151),
.B1(n_158),
.B2(n_168),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_183),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_131),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_184),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_124),
.B1(n_121),
.B2(n_126),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_155),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_162),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_154),
.C(n_147),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_195),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_197),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_183),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_161),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_159),
.B(n_166),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_153),
.C(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_203),
.B(n_163),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_189),
.B1(n_179),
.B2(n_194),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_208),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_171),
.B1(n_152),
.B2(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_189),
.A2(n_149),
.B1(n_187),
.B2(n_164),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_159),
.A3(n_170),
.B1(n_166),
.B2(n_163),
.C1(n_165),
.C2(n_146),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_214),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_202),
.C(n_200),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_192),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_209),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_215),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_205),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_114),
.B(n_145),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_210),
.B(n_212),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_205),
.C(n_221),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_225),
.B(n_226),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_219),
.A2(n_210),
.B(n_214),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_222),
.A2(n_213),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_217),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_231),
.B(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_193),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_218),
.B1(n_216),
.B2(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_236),
.C(n_165),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_232),
.A2(n_207),
.B(n_123),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_238),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_123),
.Y(n_240)
);


endmodule