module fake_jpeg_2101_n_386 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_386);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_386;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_12),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_79),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_56),
.Y(n_147)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_60),
.B(n_66),
.Y(n_139)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_12),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

CKINVDCx6p67_ASAP7_75t_R g152 ( 
.A(n_69),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g171 ( 
.A(n_70),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_12),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_71),
.B(n_72),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_19),
.B(n_16),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_73),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_11),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_74),
.B(n_83),
.Y(n_158)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_76),
.A2(n_34),
.B1(n_73),
.B2(n_89),
.Y(n_155)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_10),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_87),
.Y(n_134)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_90),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_18),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_40),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_95),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_93),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_34),
.B1(n_53),
.B2(n_33),
.Y(n_125)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_97),
.Y(n_124)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_105),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_17),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_101),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_18),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_25),
.B1(n_52),
.B2(n_51),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_42),
.B(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_42),
.B(n_5),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_107),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_28),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

AND2x4_ASAP7_75t_SL g108 ( 
.A(n_22),
.B(n_5),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g168 ( 
.A(n_108),
.B(n_76),
.CON(n_168),
.SN(n_168)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_110),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_28),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_115),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_116),
.A2(n_122),
.B1(n_135),
.B2(n_161),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_63),
.A2(n_52),
.B1(n_51),
.B2(n_25),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_118),
.A2(n_138),
.B1(n_157),
.B2(n_166),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_107),
.B1(n_104),
.B2(n_93),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_54),
.A2(n_31),
.B1(n_32),
.B2(n_47),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_129),
.A2(n_136),
.B1(n_151),
.B2(n_164),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_90),
.B(n_50),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_133),
.B(n_127),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_61),
.A2(n_31),
.B1(n_32),
.B2(n_47),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_56),
.A2(n_30),
.B1(n_44),
.B2(n_29),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_92),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_50),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_156),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_56),
.A2(n_44),
.B1(n_27),
.B2(n_26),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_64),
.B(n_6),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_150),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_155),
.A2(n_168),
.B(n_152),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_70),
.B(n_6),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_84),
.A2(n_34),
.B1(n_33),
.B2(n_53),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_99),
.A2(n_34),
.B1(n_33),
.B2(n_53),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_70),
.B(n_7),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_172),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_82),
.A2(n_7),
.B1(n_8),
.B2(n_98),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_105),
.A2(n_80),
.B1(n_78),
.B2(n_110),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_165),
.A2(n_170),
.B1(n_152),
.B2(n_147),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_101),
.A2(n_8),
.B1(n_109),
.B2(n_65),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_105),
.A2(n_18),
.B1(n_45),
.B2(n_24),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_173),
.B1(n_123),
.B2(n_140),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_59),
.A2(n_85),
.B1(n_18),
.B2(n_39),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_66),
.B(n_91),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_61),
.A2(n_73),
.B1(n_84),
.B2(n_89),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_66),
.B(n_91),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_174),
.B(n_175),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_66),
.B(n_91),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_113),
.A2(n_143),
.B(n_168),
.C(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_179),
.B(n_181),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_119),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_180),
.B(n_183),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_121),
.A2(n_114),
.B(n_158),
.C(n_115),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_119),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_188),
.B(n_196),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_124),
.A2(n_153),
.B1(n_161),
.B2(n_154),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_189),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_173),
.B1(n_135),
.B2(n_131),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_211),
.B1(n_215),
.B2(n_223),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_120),
.B(n_134),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_194),
.B(n_199),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_131),
.A2(n_142),
.B1(n_132),
.B2(n_166),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_195),
.A2(n_190),
.B1(n_178),
.B2(n_194),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_117),
.Y(n_197)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_203),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_134),
.B(n_128),
.Y(n_203)
);

AO22x1_ASAP7_75t_SL g205 ( 
.A1(n_134),
.A2(n_155),
.B1(n_111),
.B2(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_132),
.A2(n_142),
.B(n_138),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_208),
.C(n_228),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_152),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_208),
.B(n_216),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_233),
.B1(n_185),
.B2(n_215),
.Y(n_234)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_130),
.A2(n_150),
.B1(n_177),
.B2(n_111),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

OR2x6_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_205),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_137),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_155),
.A2(n_167),
.B1(n_144),
.B2(n_146),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_155),
.B(n_126),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_137),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_218),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_146),
.B(n_162),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_160),
.A2(n_162),
.B(n_123),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_160),
.B(n_167),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_145),
.A2(n_112),
.B1(n_140),
.B2(n_176),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_176),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_225),
.Y(n_260)
);

AOI32xp33_ASAP7_75t_L g225 ( 
.A1(n_112),
.A2(n_113),
.A3(n_114),
.B1(n_139),
.B2(n_148),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_154),
.B(n_158),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_201),
.Y(n_269)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_197),
.Y(n_266)
);

BUFx12_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_231),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_172),
.B(n_174),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_204),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_161),
.A2(n_54),
.B1(n_57),
.B2(n_56),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_235),
.B(n_250),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_189),
.A2(n_216),
.B1(n_229),
.B2(n_190),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_262),
.B1(n_192),
.B2(n_225),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_266),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_210),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_255),
.C(n_257),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_196),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_252),
.B(n_268),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_181),
.B(n_179),
.C(n_191),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_182),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_195),
.A2(n_205),
.B1(n_178),
.B2(n_206),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_185),
.A2(n_209),
.B1(n_223),
.B2(n_191),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_202),
.B(n_198),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_220),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_199),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_200),
.B(n_203),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_271),
.A2(n_285),
.B(n_244),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_267),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_282),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_275),
.B1(n_276),
.B2(n_238),
.Y(n_302)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_259),
.A2(n_230),
.B1(n_186),
.B2(n_187),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_217),
.B1(n_214),
.B2(n_187),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_279),
.A2(n_243),
.B1(n_246),
.B2(n_252),
.Y(n_305)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_284),
.Y(n_317)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_180),
.B(n_183),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_287),
.B(n_292),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_290),
.Y(n_319)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_251),
.C(n_264),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_219),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_296),
.Y(n_315)
);

OAI22x1_ASAP7_75t_L g294 ( 
.A1(n_246),
.A2(n_184),
.B1(n_231),
.B2(n_227),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_294),
.A2(n_239),
.B1(n_253),
.B2(n_250),
.Y(n_316)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_226),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_298),
.C(n_254),
.Y(n_318)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_271),
.A2(n_256),
.B(n_260),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_301),
.A2(n_309),
.B(n_311),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_302),
.A2(n_305),
.B1(n_314),
.B2(n_276),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_312),
.C(n_288),
.Y(n_331)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_258),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_310),
.B(n_266),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_286),
.A2(n_248),
.B(n_235),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_264),
.C(n_269),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_297),
.A2(n_248),
.B1(n_243),
.B2(n_266),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_316),
.A2(n_294),
.B1(n_295),
.B2(n_277),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_286),
.A2(n_248),
.B(n_237),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_302),
.A2(n_273),
.B1(n_275),
.B2(n_279),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_321),
.A2(n_308),
.B1(n_313),
.B2(n_300),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_304),
.B(n_278),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_323),
.C(n_325),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_283),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_303),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_337),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_280),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_326),
.B(n_314),
.Y(n_342)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_311),
.B(n_255),
.CI(n_257),
.CON(n_327),
.SN(n_327)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_328),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_317),
.B(n_284),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_306),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_330),
.B(n_334),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_335),
.C(n_338),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_332),
.A2(n_321),
.B1(n_333),
.B2(n_336),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_306),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_254),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_336),
.A2(n_285),
.B(n_305),
.Y(n_343)
);

OAI32xp33_ASAP7_75t_L g337 ( 
.A1(n_317),
.A2(n_248),
.A3(n_295),
.B1(n_277),
.B2(n_282),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_248),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_309),
.B(n_301),
.Y(n_339)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_327),
.B(n_332),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_342),
.B(n_338),
.Y(n_354)
);

NOR3xp33_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_337),
.C(n_325),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_349),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_318),
.Y(n_348)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_348),
.Y(n_357)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_335),
.B(n_308),
.Y(n_351)
);

OAI21x1_ASAP7_75t_L g362 ( 
.A1(n_351),
.A2(n_327),
.B(n_326),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_323),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_354),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_352),
.B(n_341),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_363),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_358),
.A2(n_339),
.B(n_348),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_322),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_362),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_340),
.B(n_331),
.Y(n_363)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_360),
.A2(n_340),
.B(n_347),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_366),
.Y(n_376)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_357),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_355),
.A2(n_346),
.B1(n_345),
.B2(n_347),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_370),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_349),
.Y(n_370)
);

NAND4xp25_ASAP7_75t_SL g372 ( 
.A(n_368),
.B(n_315),
.C(n_245),
.D(n_351),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_364),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_369),
.B(n_359),
.C(n_344),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_307),
.C(n_376),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_377),
.B(n_378),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_370),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_371),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_380),
.C(n_342),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_342),
.Y(n_383)
);

BUFx24_ASAP7_75t_SL g384 ( 
.A(n_383),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_384),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_381),
.Y(n_386)
);


endmodule