module fake_jpeg_13647_n_627 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_627);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_627;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_483;
wire n_236;
wire n_291;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_16),
.B(n_8),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_9),
.B(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_25),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g168 ( 
.A(n_61),
.Y(n_168)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_64),
.B(n_65),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_27),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_66),
.B(n_84),
.Y(n_134)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_71),
.B(n_78),
.Y(n_140)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_73),
.Y(n_206)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_75),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_76),
.Y(n_209)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_0),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_81),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_82),
.B(n_86),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_0),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_85),
.B(n_91),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_1),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_90),
.B(n_97),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_28),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_92),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_28),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_93),
.B(n_94),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_23),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_95),
.B(n_96),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_30),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_23),
.B(n_1),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_98),
.B(n_113),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_60),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_116),
.B(n_48),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_26),
.B(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_2),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_119),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_42),
.Y(n_120)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_121),
.Y(n_146)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_66),
.B(n_84),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_128),
.B(n_136),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_63),
.A2(n_22),
.B(n_21),
.C(n_56),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_133),
.A2(n_182),
.B(n_57),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_79),
.B(n_56),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_141),
.B(n_199),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_62),
.A2(n_54),
.B(n_44),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_153),
.B(n_177),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_158),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_70),
.A2(n_52),
.B1(n_48),
.B2(n_42),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_162),
.A2(n_70),
.B1(n_100),
.B2(n_122),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_94),
.B(n_33),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_170),
.B(n_195),
.Y(n_235)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_72),
.Y(n_175)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_104),
.Y(n_177)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_48),
.Y(n_182)
);

INVx4_ASAP7_75t_SL g184 ( 
.A(n_124),
.Y(n_184)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_123),
.Y(n_191)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_42),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_110),
.B(n_33),
.Y(n_195)
);

CKINVDCx12_ASAP7_75t_R g197 ( 
.A(n_73),
.Y(n_197)
);

CKINVDCx12_ASAP7_75t_R g257 ( 
.A(n_197),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_115),
.B(n_34),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_120),
.B(n_40),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_200),
.B(n_204),
.Y(n_253)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_67),
.B(n_34),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g205 ( 
.A(n_125),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_205),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_108),
.B(n_32),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_207),
.B(n_32),
.Y(n_262)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_162),
.A2(n_136),
.B1(n_172),
.B2(n_164),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_210),
.A2(n_214),
.B1(n_246),
.B2(n_263),
.Y(n_305)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_213),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_134),
.A2(n_75),
.B1(n_74),
.B2(n_126),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_99),
.B1(n_117),
.B2(n_76),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_215),
.A2(n_265),
.B1(n_173),
.B2(n_196),
.Y(n_300)
);

OR2x2_ASAP7_75t_SL g216 ( 
.A(n_133),
.B(n_169),
.Y(n_216)
);

NOR2x1_ASAP7_75t_R g320 ( 
.A(n_216),
.B(n_146),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_176),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_217),
.B(n_252),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_218),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_219),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_223),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_224),
.Y(n_311)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

BUFx2_ASAP7_75t_SL g306 ( 
.A(n_225),
.Y(n_306)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_228),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_148),
.A2(n_48),
.B1(n_42),
.B2(n_114),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_229),
.A2(n_258),
.B(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_SL g230 ( 
.A(n_163),
.B(n_54),
.C(n_22),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_230),
.B(n_236),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_131),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_234),
.Y(n_292)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_237),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_238),
.B(n_264),
.Y(n_323)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_137),
.Y(n_240)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_240),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_37),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_241),
.B(n_248),
.Y(n_333)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_183),
.A2(n_83),
.B1(n_88),
.B2(n_87),
.Y(n_246)
);

AO22x2_ASAP7_75t_L g247 ( 
.A1(n_129),
.A2(n_68),
.B1(n_121),
.B2(n_119),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g317 ( 
.A1(n_247),
.A2(n_249),
.B1(n_185),
.B2(n_178),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_140),
.B(n_37),
.Y(n_248)
);

AOI22x1_ASAP7_75t_L g249 ( 
.A1(n_161),
.A2(n_102),
.B1(n_89),
.B2(n_109),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_158),
.Y(n_250)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_186),
.Y(n_251)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_168),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_158),
.Y(n_255)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_155),
.B(n_44),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_256),
.B(n_268),
.Y(n_331)
);

NAND2xp33_ASAP7_75t_SL g258 ( 
.A(n_161),
.B(n_112),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_138),
.Y(n_259)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_138),
.Y(n_260)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_260),
.Y(n_324)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_132),
.Y(n_261)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_261),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_275),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_135),
.A2(n_69),
.B1(n_57),
.B2(n_40),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_174),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_173),
.A2(n_107),
.B1(n_58),
.B2(n_45),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_143),
.Y(n_266)
);

INVx4_ASAP7_75t_SL g318 ( 
.A(n_266),
.Y(n_318)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_129),
.Y(n_267)
);

INVx11_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_168),
.B(n_131),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_161),
.A2(n_114),
.B1(n_92),
.B2(n_58),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_269),
.A2(n_272),
.B1(n_273),
.B2(n_280),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_180),
.A2(n_45),
.B(n_41),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_143),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_166),
.A2(n_92),
.B1(n_41),
.B2(n_26),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_130),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_274),
.A2(n_278),
.B1(n_156),
.B2(n_198),
.Y(n_322)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_154),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_201),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_276),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_184),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_279),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_147),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_150),
.B(n_7),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_151),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_165),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_282),
.Y(n_319)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_167),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_171),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_283),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_232),
.B(n_152),
.C(n_144),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_289),
.B(n_307),
.C(n_313),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_215),
.A2(n_224),
.B1(n_216),
.B2(n_265),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_293),
.A2(n_315),
.B1(n_327),
.B2(n_336),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_221),
.B(n_201),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_294),
.B(n_301),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_253),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_314),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_300),
.B(n_317),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_235),
.B(n_159),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_220),
.B(n_190),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_222),
.B(n_151),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_308),
.B(n_310),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_226),
.B(n_202),
.Y(n_310)
);

XNOR2x1_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_157),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_228),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_210),
.B(n_146),
.C(n_166),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_231),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_249),
.A2(n_178),
.B1(n_202),
.B2(n_196),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_320),
.B(n_240),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_322),
.A2(n_332),
.B1(n_211),
.B2(n_242),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_227),
.B(n_156),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_326),
.B(n_334),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_273),
.A2(n_198),
.B1(n_142),
.B2(n_145),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_246),
.A2(n_185),
.B1(n_181),
.B2(n_179),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_329),
.A2(n_255),
.B1(n_250),
.B2(n_280),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_254),
.A2(n_145),
.B1(n_205),
.B2(n_191),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_243),
.B(n_142),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_269),
.A2(n_181),
.B1(n_206),
.B2(n_10),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_247),
.A2(n_206),
.B1(n_9),
.B2(n_10),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_337),
.A2(n_219),
.B(n_223),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_231),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_338),
.B(n_245),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_247),
.A2(n_206),
.B1(n_12),
.B2(n_13),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_341),
.A2(n_233),
.B1(n_212),
.B2(n_242),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_309),
.B(n_271),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_343),
.B(n_348),
.Y(n_399)
);

INVx11_ASAP7_75t_L g344 ( 
.A(n_335),
.Y(n_344)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_344),
.Y(n_404)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_247),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_363),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_331),
.B(n_233),
.Y(n_348)
);

AO22x2_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_258),
.B1(n_212),
.B2(n_266),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_384),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_350),
.A2(n_337),
.B1(n_317),
.B2(n_312),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g352 ( 
.A1(n_293),
.A2(n_259),
.B(n_260),
.Y(n_352)
);

OAI21xp33_ASAP7_75t_SL g395 ( 
.A1(n_352),
.A2(n_367),
.B(n_287),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_353),
.A2(n_346),
.B1(n_352),
.B2(n_359),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_233),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_SL g393 ( 
.A(n_356),
.B(n_359),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_287),
.B(n_270),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_294),
.B(n_244),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_361),
.B(n_362),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_237),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_264),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_311),
.A2(n_276),
.B1(n_267),
.B2(n_272),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_364),
.A2(n_339),
.B1(n_296),
.B2(n_328),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_257),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_368),
.Y(n_398)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_284),
.B(n_340),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_377),
.Y(n_417)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

NAND2x1p5_ASAP7_75t_L g371 ( 
.A(n_323),
.B(n_218),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_371),
.A2(n_372),
.B(n_290),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_373),
.Y(n_418)
);

INVx13_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_374),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_304),
.Y(n_425)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

BUFx12_ASAP7_75t_L g377 ( 
.A(n_297),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_340),
.B(n_8),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_381),
.Y(n_419)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_298),
.Y(n_380)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_380),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_286),
.B(n_12),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_323),
.B(n_12),
.C(n_13),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_323),
.C(n_307),
.Y(n_389)
);

AO22x1_ASAP7_75t_SL g384 ( 
.A1(n_305),
.A2(n_13),
.B1(n_317),
.B2(n_315),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_292),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_288),
.Y(n_420)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_386),
.Y(n_413)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_334),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_302),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_395),
.B(n_400),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_397),
.A2(n_401),
.B(n_409),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_357),
.A2(n_305),
.B1(n_311),
.B2(n_322),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_372),
.A2(n_289),
.B(n_330),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_402),
.A2(n_414),
.B1(n_415),
.B2(n_424),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_354),
.B(n_301),
.C(n_340),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_405),
.B(n_356),
.C(n_371),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_406),
.Y(n_435)
);

OAI32xp33_ASAP7_75t_L g407 ( 
.A1(n_355),
.A2(n_319),
.A3(n_324),
.B1(n_302),
.B2(n_295),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_410),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_372),
.A2(n_336),
.B(n_324),
.Y(n_409)
);

AOI22x1_ASAP7_75t_L g415 ( 
.A1(n_346),
.A2(n_295),
.B1(n_318),
.B2(n_288),
.Y(n_415)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_420),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_303),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_422),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_383),
.B(n_325),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_376),
.B(n_325),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_358),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_346),
.A2(n_384),
.B1(n_359),
.B2(n_387),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_375),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_410),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_428),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_351),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_427),
.B(n_437),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_423),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_399),
.B(n_419),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_430),
.B(n_440),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_388),
.A2(n_357),
.B1(n_370),
.B2(n_386),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_432),
.A2(n_441),
.B1(n_447),
.B2(n_454),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_404),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_433),
.B(n_434),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_422),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_385),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_411),
.Y(n_438)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_438),
.Y(n_463)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_411),
.Y(n_439)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_439),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_361),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_388),
.A2(n_384),
.B1(n_367),
.B2(n_355),
.Y(n_441)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

BUFx5_ASAP7_75t_L g444 ( 
.A(n_392),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_444),
.B(n_390),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_421),
.B(n_413),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_457),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_402),
.A2(n_354),
.B1(n_347),
.B2(n_352),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_398),
.B(n_343),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_448),
.B(n_436),
.Y(n_490)
);

BUFx8_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_451),
.B(n_461),
.Y(n_464)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_412),
.Y(n_452)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_391),
.A2(n_350),
.B1(n_371),
.B2(n_349),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_412),
.Y(n_455)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_425),
.C(n_393),
.Y(n_480)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_366),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_459),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_417),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_408),
.B(n_403),
.Y(n_460)
);

NOR2x1_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_408),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_403),
.B(n_356),
.Y(n_461)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_462),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_405),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_466),
.B(n_468),
.C(n_480),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_446),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_381),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_470),
.B(n_473),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_460),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_430),
.B(n_459),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_474),
.B(n_475),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_427),
.B(n_348),
.Y(n_475)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_477),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_437),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_479),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_393),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_494),
.C(n_443),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_431),
.A2(n_397),
.B1(n_409),
.B2(n_394),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_454),
.Y(n_495)
);

AOI221xp5_ASAP7_75t_L g485 ( 
.A1(n_440),
.A2(n_401),
.B1(n_407),
.B2(n_400),
.C(n_406),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_485),
.A2(n_490),
.B1(n_435),
.B2(n_426),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_431),
.B(n_389),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_486),
.B(n_492),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_449),
.A2(n_394),
.B1(n_353),
.B2(n_415),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_489),
.A2(n_450),
.B(n_349),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_447),
.B(n_382),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_453),
.A2(n_396),
.B(n_349),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_493),
.A2(n_429),
.B(n_435),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_378),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_495),
.A2(n_489),
.B1(n_488),
.B2(n_481),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_499),
.A2(n_514),
.B(n_517),
.Y(n_527)
);

OAI21xp33_ASAP7_75t_L g501 ( 
.A1(n_491),
.A2(n_429),
.B(n_445),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_501),
.B(n_469),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_502),
.B(n_471),
.Y(n_529)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_463),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_503),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_465),
.A2(n_434),
.B1(n_428),
.B2(n_442),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_504),
.B(n_513),
.Y(n_544)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_477),
.Y(n_506)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_506),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_442),
.Y(n_507)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_507),
.Y(n_537)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_509),
.B(n_510),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_432),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_494),
.Y(n_526)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_478),
.Y(n_511)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_468),
.B(n_480),
.C(n_464),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_523),
.C(n_486),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_483),
.A2(n_436),
.B1(n_439),
.B2(n_455),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_493),
.A2(n_450),
.B(n_458),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_465),
.A2(n_438),
.B1(n_452),
.B2(n_441),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_515),
.A2(n_518),
.B1(n_519),
.B2(n_488),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_472),
.A2(n_450),
.B(n_457),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_487),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_471),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_469),
.B(n_444),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_520),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_484),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_464),
.B(n_396),
.C(n_433),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_524),
.B(n_528),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_525),
.B(n_521),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_533),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_509),
.B(n_492),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_529),
.A2(n_500),
.B1(n_497),
.B2(n_506),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_498),
.B(n_482),
.C(n_476),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_534),
.Y(n_553)
);

NOR2xp67_ASAP7_75t_L g558 ( 
.A(n_531),
.B(n_505),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_498),
.B(n_476),
.C(n_472),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_535),
.Y(n_555)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_538),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_481),
.C(n_467),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_539),
.B(n_545),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_512),
.B(n_467),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_542),
.B(n_547),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_495),
.B(n_463),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_SL g554 ( 
.A(n_543),
.B(n_520),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_380),
.C(n_404),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_505),
.B(n_345),
.Y(n_546)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_546),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_516),
.B(n_297),
.C(n_316),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_534),
.A2(n_500),
.B(n_522),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_549),
.B(n_562),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_552),
.A2(n_504),
.B1(n_540),
.B2(n_541),
.Y(n_571)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_554),
.Y(n_584)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_558),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_559),
.B(n_564),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_542),
.B(n_499),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_561),
.B(n_539),
.C(n_533),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_544),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_536),
.Y(n_563)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_563),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_548),
.A2(n_497),
.B1(n_519),
.B2(n_518),
.Y(n_564)
);

BUFx12_ASAP7_75t_L g565 ( 
.A(n_527),
.Y(n_565)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_565),
.Y(n_585)
);

A2O1A1O1Ixp25_ASAP7_75t_L g566 ( 
.A1(n_530),
.A2(n_514),
.B(n_507),
.C(n_511),
.D(n_508),
.Y(n_566)
);

AOI21xp33_ASAP7_75t_L g580 ( 
.A1(n_566),
.A2(n_525),
.B(n_517),
.Y(n_580)
);

BUFx24_ASAP7_75t_SL g568 ( 
.A(n_537),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_568),
.B(n_496),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_569),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_571),
.B(n_349),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_SL g572 ( 
.A1(n_555),
.A2(n_496),
.B1(n_532),
.B2(n_503),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_572),
.A2(n_576),
.B1(n_547),
.B2(n_532),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_574),
.B(n_575),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_553),
.B(n_543),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_555),
.A2(n_550),
.B1(n_545),
.B2(n_559),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_560),
.B(n_526),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_577),
.B(n_579),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_567),
.B(n_524),
.C(n_528),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_580),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_556),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_581),
.B(n_567),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_561),
.B(n_418),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_583),
.B(n_551),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_570),
.A2(n_566),
.B(n_565),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_587),
.B(n_598),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_SL g604 ( 
.A1(n_589),
.A2(n_599),
.B1(n_588),
.B2(n_584),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_585),
.A2(n_565),
.B1(n_554),
.B2(n_418),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_590),
.Y(n_601)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_591),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_592),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_593),
.B(n_579),
.Y(n_605)
);

A2O1A1Ixp33_ASAP7_75t_SL g595 ( 
.A1(n_585),
.A2(n_344),
.B(n_551),
.C(n_390),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_595),
.B(n_597),
.C(n_571),
.Y(n_603)
);

AOI21x1_ASAP7_75t_L g597 ( 
.A1(n_573),
.A2(n_557),
.B(n_321),
.Y(n_597)
);

NOR2x1_ASAP7_75t_L g598 ( 
.A(n_569),
.B(n_373),
.Y(n_598)
);

INVx6_ASAP7_75t_L g599 ( 
.A(n_581),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_582),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_600),
.A2(n_608),
.B(n_590),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_596),
.B(n_582),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_602),
.B(n_604),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_603),
.B(n_605),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_594),
.B(n_576),
.Y(n_608)
);

AOI322xp5_ASAP7_75t_L g610 ( 
.A1(n_601),
.A2(n_607),
.A3(n_609),
.B1(n_600),
.B2(n_606),
.C1(n_584),
.C2(n_602),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_610),
.B(n_611),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_601),
.Y(n_611)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_612),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_600),
.A2(n_586),
.B(n_595),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_613),
.A2(n_614),
.B(n_296),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_600),
.A2(n_595),
.B(n_592),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_616),
.B(n_578),
.C(n_373),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_619),
.B(n_620),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_617),
.A2(n_615),
.B(n_610),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_621),
.A2(n_618),
.B(n_316),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_623),
.B(n_622),
.C(n_291),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_SL g625 ( 
.A(n_624),
.B(n_377),
.C(n_374),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_625),
.B(n_321),
.C(n_304),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_626),
.A2(n_339),
.B1(n_306),
.B2(n_318),
.Y(n_627)
);


endmodule