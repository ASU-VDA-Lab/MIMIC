module fake_jpeg_15634_n_27 (n_3, n_2, n_1, n_0, n_4, n_5, n_27);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_27;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

HAxp5_ASAP7_75t_SL g6 ( 
.A(n_0),
.B(n_3),
.CON(n_6),
.SN(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_3),
.Y(n_7)
);

BUFx2_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_5),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_0),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_14),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_1),
.C(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_12),
.B(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_6),
.B(n_2),
.CI(n_7),
.CON(n_16),
.SN(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_18),
.B1(n_10),
.B2(n_8),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_18),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_23),
.B(n_19),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_17),
.C(n_14),
.Y(n_23)
);

AOI322xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_25),
.A3(n_19),
.B1(n_13),
.B2(n_20),
.C1(n_16),
.C2(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_16),
.Y(n_27)
);


endmodule