module real_jpeg_17377_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AND2x2_ASAP7_75t_L g60 ( 
.A(n_0),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_0),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_0),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_0),
.B(n_134),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_0),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_0),
.B(n_410),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_1),
.B(n_37),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_1),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_33),
.Y(n_32)
);

AOI22x1_ASAP7_75t_L g40 ( 
.A1(n_2),
.A2(n_9),
.B1(n_41),
.B2(n_45),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_2),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_2),
.B(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_2),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_2),
.B(n_134),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_3),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_3),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_3),
.B(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_3),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_3),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_3),
.B(n_330),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_4),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_4),
.Y(n_312)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_5),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_5),
.Y(n_365)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_5),
.Y(n_407)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_6),
.Y(n_292)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_7),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_7),
.Y(n_199)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_7),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_8),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_8),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_8),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_8),
.B(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_8),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_8),
.B(n_44),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_8),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_9),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_9),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_9),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_9),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_9),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_9),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_9),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_9),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_10),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_10),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_10),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_10),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_10),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_10),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_10),
.B(n_370),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_11),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_28),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g67 ( 
.A(n_12),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_12),
.B(n_83),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_12),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_80),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_12),
.B(n_33),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_12),
.B(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_14),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_14),
.B(n_422),
.Y(n_421)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_15),
.Y(n_155)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_381),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_206),
.B(n_380),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_170),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_20),
.B(n_170),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_96),
.Y(n_20)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_21),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_64),
.C(n_85),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2x1_ASAP7_75t_SL g172 ( 
.A(n_23),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.C(n_50),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_24),
.B(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_26),
.B(n_143),
.Y(n_395)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_27),
.B(n_32),
.C(n_36),
.Y(n_87)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_37),
.Y(n_192)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_38),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_39),
.A2(n_40),
.B1(n_50),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_40),
.A2(n_223),
.B(n_231),
.Y(n_222)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_49),
.Y(n_230)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_49),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_49),
.Y(n_414)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_50),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.C(n_60),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_51),
.A2(n_52),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_51),
.A2(n_52),
.B1(n_60),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g396 ( 
.A(n_52),
.B(n_104),
.C(n_152),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_55),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_56),
.B(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_59),
.Y(n_196)
);

INVx11_ASAP7_75t_SL g184 ( 
.A(n_60),
.Y(n_184)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_65),
.A2(n_85),
.B1(n_86),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_65),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_78),
.C(n_81),
.Y(n_65)
);

XOR2x2_ASAP7_75t_L g200 ( 
.A(n_66),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.C(n_75),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_67),
.A2(n_75),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_67),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_67),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_71),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_72),
.B(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx13_ASAP7_75t_SL g221 ( 
.A(n_75),
.Y(n_221)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_77),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_80),
.Y(n_285)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2x1_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_89),
.C(n_92),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_89),
.A2(n_90),
.B1(n_241),
.B2(n_242),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_90),
.B(n_238),
.C(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_148),
.B1(n_168),
.B2(n_169),
.Y(n_96)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_138),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_98),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_109),
.C(n_124),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_99),
.B(n_109),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_104),
.C(n_105),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_107),
.Y(n_328)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_108),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.C(n_119),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_110),
.A2(n_119),
.B1(n_120),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_115),
.B(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_118),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_119),
.B(n_259),
.C(n_263),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_119),
.A2(n_120),
.B1(n_263),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_129),
.C(n_133),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_139),
.B(n_389),
.C(n_390),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_140),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_142),
.B(n_145),
.C(n_147),
.Y(n_399)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_148),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_149),
.B(n_157),
.C(n_158),
.Y(n_400)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_152),
.A2(n_404),
.B1(n_405),
.B2(n_408),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_152),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_153),
.B(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_159),
.B(n_162),
.C(n_163),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_168),
.B(n_385),
.C(n_386),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.C(n_178),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_175),
.Y(n_212)
);

XOR2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_200),
.C(n_203),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_193),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_182),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_185),
.B(n_193),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_186),
.B(n_191),
.Y(n_268)
);

NOR2x1_ASAP7_75t_R g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_190),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_194),
.A2(n_197),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_197),
.B(n_342),
.C(n_344),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_197),
.A2(n_256),
.B1(n_344),
.B2(n_345),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_198),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_273),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.C(n_248),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_211),
.B(n_214),
.Y(n_379)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.C(n_245),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_215),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_245),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.C(n_237),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_222),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_220),
.B(n_308),
.C(n_313),
.Y(n_307)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_238),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_240),
.Y(n_282)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_239),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_239),
.A2(n_351),
.B1(n_352),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_244),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_271),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_271),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.C(n_269),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_269),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.C(n_267),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_268),
.Y(n_280)
);

XOR2x2_ASAP7_75t_L g317 ( 
.A(n_259),
.B(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.C(n_379),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_298),
.B(n_378),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_296),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_277),
.B(n_296),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.C(n_293),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_279),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_293),
.B1(n_294),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.C(n_286),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_283),
.Y(n_306)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.Y(n_286)
);

AO22x1_ASAP7_75t_SL g332 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_291),
.Y(n_333)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_292),
.Y(n_331)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_292),
.Y(n_354)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_320),
.B(n_377),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g377 ( 
.A(n_300),
.B(n_304),
.Y(n_377)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.C(n_316),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_317),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_313),
.Y(n_324)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI21x1_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_336),
.B(n_376),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_334),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_322),
.B(n_334),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.C(n_332),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_325),
.A2(n_326),
.B1(n_332),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_327),
.B(n_329),
.Y(n_343)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_332),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_369),
.Y(n_368)
);

AOI21x1_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_348),
.B(n_375),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_341),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_341),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_342),
.A2(n_343),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_358),
.B(n_374),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_355),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_350),
.B(n_355),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_368),
.B(n_373),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_366),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_366),
.Y(n_373)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_426),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g426 ( 
.A(n_384),
.B(n_387),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_401),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_400),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_399),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_396),
.B1(n_397),
.B2(n_398),
.Y(n_394)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_395),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_396),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_415),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_409),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);


endmodule