module fake_jpeg_25792_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_0),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_24),
.B1(n_33),
.B2(n_28),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_66),
.B1(n_68),
.B2(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_63),
.Y(n_88)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_24),
.B1(n_23),
.B2(n_33),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_70),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_38),
.Y(n_73)
);

OR2x4_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_18),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_76),
.Y(n_110)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_23),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_31),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_31),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_87),
.B(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_94),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_17),
.C(n_31),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_56),
.C(n_82),
.Y(n_117)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_93),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_97),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_29),
.B1(n_22),
.B2(n_31),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_114),
.B1(n_82),
.B2(n_67),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_99),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_2),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_34),
.B1(n_22),
.B2(n_27),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_104),
.Y(n_126)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_71),
.B(n_27),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_1),
.B(n_2),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_79),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_15),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_4),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_18),
.B1(n_30),
.B2(n_27),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_55),
.A2(n_27),
.B1(n_30),
.B2(n_26),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_117),
.Y(n_146)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_64),
.B1(n_69),
.B2(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_138),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_26),
.B(n_11),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_96),
.C(n_114),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_56),
.B1(n_83),
.B2(n_4),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_92),
.B1(n_100),
.B2(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_2),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_102),
.B1(n_85),
.B2(n_108),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_R g134 ( 
.A(n_93),
.B(n_3),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_6),
.B(n_8),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_105),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_3),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_85),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_5),
.Y(n_144)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_86),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_93),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_163),
.B(n_120),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_151),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_119),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_100),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_102),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_153),
.B(n_125),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_161),
.B1(n_125),
.B2(n_121),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_95),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_103),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_6),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_163),
.B(n_134),
.C(n_162),
.D(n_138),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_94),
.B1(n_7),
.B2(n_8),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_169),
.B(n_172),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_117),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_175),
.C(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_182),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_122),
.B(n_126),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_126),
.B(n_116),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_174),
.B(n_177),
.C(n_162),
.Y(n_201)
);

XOR2x2_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_127),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_139),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_115),
.B(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_161),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_121),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_137),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_184),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_200),
.B(n_201),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_189),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_150),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_147),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_197),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_157),
.C(n_156),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_175),
.C(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_198),
.A2(n_169),
.B1(n_174),
.B2(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_166),
.B(n_162),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_208),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_191),
.Y(n_219)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_159),
.B1(n_145),
.B2(n_154),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_213),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_164),
.B1(n_177),
.B2(n_149),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_172),
.C(n_142),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_142),
.B(n_160),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_214),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_217),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_186),
.C(n_195),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_221),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_192),
.B(n_189),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_212),
.B1(n_187),
.B2(n_210),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_230),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_208),
.B1(n_204),
.B2(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_197),
.B1(n_206),
.B2(n_208),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_203),
.B(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_231),
.B(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_204),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_233),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_202),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_238),
.B(n_239),
.Y(n_241)
);

OAI321xp33_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_202),
.A3(n_220),
.B1(n_211),
.B2(n_217),
.C(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_226),
.C(n_219),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_226),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_244),
.A2(n_245),
.B(n_243),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_241),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_221),
.Y(n_247)
);


endmodule