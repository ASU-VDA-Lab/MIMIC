module real_jpeg_32478_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_578;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_0),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_0),
.Y(n_389)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_0),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_1),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_1),
.B(n_63),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_1),
.B(n_142),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_1),
.B(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_SL g342 ( 
.A(n_1),
.B(n_256),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_1),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_1),
.B(n_387),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_3),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_3),
.B(n_317),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_3),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_3),
.B(n_349),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_3),
.B(n_337),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_3),
.B(n_475),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_3),
.B(n_387),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_21),
.B(n_22),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_5),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_5),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_5),
.B(n_227),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g258 ( 
.A(n_5),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_5),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_5),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_5),
.B(n_73),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_5),
.B(n_478),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_6),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_6),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_6),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_6),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_6),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_6),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_6),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_6),
.B(n_329),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_7),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_9),
.Y(n_187)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_9),
.Y(n_527)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_10),
.Y(n_257)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_10),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_244),
.Y(n_243)
);

NAND2x1_ASAP7_75t_L g321 ( 
.A(n_11),
.B(n_97),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_11),
.B(n_349),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_11),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_11),
.B(n_490),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g525 ( 
.A(n_11),
.B(n_526),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_11),
.B(n_533),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_12),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_12),
.B(n_432),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_12),
.B(n_63),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_12),
.B(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_12),
.B(n_206),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_12),
.B(n_539),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_12),
.B(n_547),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_23),
.Y(n_22)
);

NAND2x1_ASAP7_75t_SL g36 ( 
.A(n_14),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_14),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_14),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_14),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_14),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_14),
.B(n_99),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_14),
.B(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_15),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_69),
.Y(n_68)
);

NAND2x1_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_16),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_16),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_16),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_16),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_16),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_17),
.Y(n_133)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_17),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_18),
.B(n_190),
.Y(n_189)
);

NAND2x1_ASAP7_75t_L g229 ( 
.A(n_18),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_18),
.B(n_259),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_18),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_18),
.B(n_452),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_18),
.B(n_495),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_18),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_18),
.B(n_522),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_19),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_19),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_19),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_19),
.B(n_185),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_19),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_19),
.B(n_387),
.Y(n_386)
);

O2A1O1Ixp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_299),
.B(n_574),
.C(n_588),
.Y(n_23)
);

OAI211xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_175),
.B(n_283),
.C(n_284),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g571 ( 
.A(n_25),
.B(n_572),
.Y(n_571)
);

NOR2xp67_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_146),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_26),
.B(n_146),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_108),
.C(n_123),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_27),
.B(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_76),
.B(n_107),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_28),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_47),
.C(n_60),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_29),
.B(n_47),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_30),
.B(n_36),
.C(n_40),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_34),
.Y(n_171)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_34),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_34),
.Y(n_231)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_34),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_41),
.B2(n_46),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_44),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_45),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.C(n_54),
.Y(n_47)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_48),
.B(n_51),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_50),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_53),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_54),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_56),
.B(n_324),
.Y(n_471)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g533 ( 
.A(n_58),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_59),
.Y(n_346)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_60),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_66),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_67),
.C(n_75),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_65),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_75),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_68),
.B1(n_111),
.B2(n_114),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_67),
.B(n_111),
.C(n_115),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_96),
.C(n_98),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_72),
.A2(n_75),
.B1(n_98),
.B2(n_188),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_74),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_74),
.Y(n_475)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_74),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_94),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_94),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_77),
.A2(n_78),
.B1(n_94),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2x1_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_90),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_89),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_83),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_89),
.C(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_87),
.Y(n_456)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_88),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_92),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_93),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_94),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.C(n_106),
.Y(n_94)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_97),
.Y(n_297)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_98),
.A2(n_184),
.B1(n_188),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_101),
.B(n_106),
.Y(n_198)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_103),
.Y(n_292)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_103),
.Y(n_341)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_106),
.B(n_200),
.C(n_208),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_106),
.B(n_209),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_108),
.B(n_123),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_121),
.C(n_122),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_109),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_111),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_114),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_157),
.C(n_158),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_113),
.Y(n_236)
);

NOR2xp67_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_121),
.B(n_122),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_135),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_145),
.C(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_130),
.C(n_134),
.Y(n_148)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_144),
.B2(n_145),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_173),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_148),
.B(n_149),
.C(n_173),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_159),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_151),
.B(n_156),
.C(n_159),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_157),
.B(n_162),
.C(n_168),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_168),
.B1(n_169),
.B2(n_172),
.Y(n_159)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_161),
.A2(n_162),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_161),
.B(n_290),
.C(n_295),
.Y(n_584)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_277),
.B(n_282),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_266),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_177),
.B(n_266),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_R g177 ( 
.A(n_178),
.B(n_214),
.C(n_217),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_178),
.A2(n_179),
.B1(n_214),
.B2(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_195),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_180),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_192),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_181),
.B(n_183),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_189),
.Y(n_183)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_187),
.Y(n_384)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_192),
.B(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_196),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_SL g267 ( 
.A(n_199),
.B(n_268),
.C(n_270),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_200),
.B(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.C(n_205),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_202),
.Y(n_240)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_213),
.Y(n_582)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_214),
.Y(n_361)
);

XNOR2x2_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_218),
.B(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_241),
.C(n_263),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.C(n_239),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_220),
.B(n_224),
.C(n_239),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_224),
.Y(n_372)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B(n_237),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_229),
.B(n_238),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_232),
.Y(n_402)
);

INVx3_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_239),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_241),
.B(n_264),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_252),
.B(n_262),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.C(n_250),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_243),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_SL g354 ( 
.A(n_243),
.B(n_247),
.C(n_250),
.Y(n_354)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_247),
.A2(n_250),
.B1(n_251),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_SL g262 ( 
.A(n_253),
.B(n_258),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_253),
.B(n_258),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_253),
.B(n_258),
.Y(n_355)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_257),
.Y(n_400)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_257),
.Y(n_496)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_272),
.C(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_277),
.B(n_573),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_280),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_285),
.B(n_286),
.Y(n_587)
);

BUFx24_ASAP7_75t_SL g592 ( 
.A(n_286),
.Y(n_592)
);

FAx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_288),
.CI(n_289),
.CON(n_286),
.SN(n_286)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_294),
.A2(n_295),
.B1(n_578),
.B2(n_579),
.Y(n_577)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_298),
.B(n_580),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_571),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_410),
.B(n_568),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_362),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_302),
.A2(n_569),
.B(n_570),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_359),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_L g570 ( 
.A(n_303),
.B(n_359),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.C(n_357),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_305),
.B(n_357),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_308),
.B(n_409),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_332),
.C(n_350),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_366),
.Y(n_365)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.C(n_326),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_311),
.B(n_313),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_314),
.A2(n_315),
.B1(n_326),
.B2(n_327),
.Y(n_437)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_319),
.B(n_322),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_316),
.B(n_377),
.Y(n_376)
);

AOI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_323),
.B(n_325),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_319),
.A2(n_320),
.B1(n_325),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OA21x2_ASAP7_75t_SL g421 ( 
.A1(n_327),
.A2(n_328),
.B(n_331),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_333),
.A2(n_351),
.B1(n_352),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_343),
.C(n_347),
.Y(n_333)
);

XOR2x1_ASAP7_75t_L g406 ( 
.A(n_334),
.B(n_407),
.Y(n_406)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_340),
.C(n_342),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_335),
.A2(n_336),
.B1(n_342),
.B2(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_338),
.Y(n_492)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_340),
.B(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_342),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_343),
.A2(n_344),
.B1(n_347),
.B2(n_348),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_352)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_354),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_408),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_363),
.B(n_408),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_368),
.C(n_373),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_365),
.B(n_369),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_373),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_401),
.C(n_404),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_374),
.A2(n_375),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.C(n_390),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_376),
.B(n_460),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_379),
.A2(n_390),
.B1(n_391),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_385),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_380),
.A2(n_381),
.B1(n_385),
.B2(n_386),
.Y(n_457)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_389),
.Y(n_549)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_396),
.C(n_397),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_392),
.A2(n_393),
.B1(n_397),
.B2(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_396),
.B(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_400),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_401),
.A2(n_405),
.B1(n_406),
.B2(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_401),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_464),
.B(n_566),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_438),
.B(n_441),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_412),
.B(n_438),
.C(n_567),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_417),
.C(n_434),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_413),
.B(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_417),
.B(n_435),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.C(n_422),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_421),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_422),
.B(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_428),
.C(n_430),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_423),
.B(n_480),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_424),
.A2(n_425),
.B1(n_426),
.B2(n_427),
.Y(n_470)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_428),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.Y(n_480)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_462),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_442),
.B(n_462),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.C(n_458),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_443),
.B(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_445),
.B(n_459),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_449),
.C(n_457),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_446),
.B(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_457),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.C(n_454),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_450),
.B(n_454),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_451),
.B(n_515),
.Y(n_514)
);

INVx3_ASAP7_75t_SL g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_456),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_465),
.A2(n_483),
.B(n_565),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_481),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_466),
.B(n_481),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_469),
.C(n_479),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_467),
.B(n_563),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_469),
.B(n_479),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.C(n_472),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_470),
.B(n_471),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_472),
.B(n_509),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_476),
.Y(n_472)
);

AO22x1_ASAP7_75t_L g505 ( 
.A1(n_473),
.A2(n_474),
.B1(n_476),
.B2(n_477),
.Y(n_505)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_484),
.A2(n_560),
.B(n_564),
.Y(n_483)
);

OAI21x1_ASAP7_75t_SL g484 ( 
.A1(n_485),
.A2(n_517),
.B(n_559),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_506),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_486),
.B(n_506),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_499),
.C(n_505),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_487),
.A2(n_488),
.B1(n_555),
.B2(n_557),
.Y(n_554)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_493),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_512),
.C(n_513),
.Y(n_511)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_497),
.Y(n_493)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_494),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_497),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_499),
.A2(n_500),
.B1(n_505),
.B2(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_501),
.B(n_504),
.Y(n_535)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_505),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_507),
.A2(n_508),
.B1(n_510),
.B2(n_516),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_507),
.B(n_511),
.C(n_514),
.Y(n_561)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_510),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_511),
.B(n_514),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_552),
.B(n_558),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_519),
.A2(n_536),
.B(n_551),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_528),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_520),
.B(n_528),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_525),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_521),
.B(n_525),
.Y(n_544)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx8_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_525),
.B(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_535),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_530),
.A2(n_531),
.B1(n_532),
.B2(n_534),
.Y(n_529)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_530),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_534),
.C(n_535),
.Y(n_553)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_545),
.B(n_550),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_544),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_544),
.Y(n_550)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx3_ASAP7_75t_SL g547 ( 
.A(n_548),
.Y(n_547)
);

INVx8_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_554),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_554),
.Y(n_558)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_555),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g560 ( 
.A(n_561),
.B(n_562),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_561),
.B(n_562),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_586),
.Y(n_574)
);

AOI221xp5_ASAP7_75t_L g575 ( 
.A1(n_576),
.A2(n_577),
.B1(n_583),
.B2(n_584),
.C(n_585),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_576),
.A2(n_577),
.B1(n_583),
.B2(n_584),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_577),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_579),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_579),
.B(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_584),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_585),
.B(n_590),
.Y(n_589)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);


endmodule