module fake_netlist_6_809_n_2073 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2073);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2073;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1950;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2052;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_186),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_120),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_106),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_149),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_100),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_58),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_27),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_119),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_195),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_42),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_152),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_161),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_114),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_75),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_39),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_103),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_86),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_40),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_20),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_126),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_144),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_38),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_74),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_32),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_148),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_138),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_45),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_4),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_197),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_25),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_61),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_40),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_88),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_29),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_59),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_110),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_20),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_167),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_1),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_2),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_169),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_166),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_153),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_158),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_140),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_73),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_180),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_11),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_198),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_202),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_13),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_117),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_66),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_123),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_17),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_37),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_89),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_90),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_168),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_189),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_177),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_30),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_124),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_56),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_94),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_83),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_23),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_93),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_101),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_102),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_24),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_75),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_109),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_155),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_62),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_61),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_49),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_52),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_111),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_22),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_97),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_51),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_39),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_108),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_1),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_184),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_7),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_139),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_131),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_42),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_9),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_178),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_57),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_96),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_160),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_2),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_170),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_69),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_6),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_190),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_116),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_78),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_85),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_157),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_58),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_154),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_52),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_71),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_127),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_51),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_162),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_147),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_62),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_19),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_72),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_48),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_44),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_11),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_151),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_23),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_156),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_73),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_57),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_133),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_91),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_9),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_87),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_45),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_71),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_78),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_81),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_163),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_82),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_80),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_193),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_92),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_16),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_142),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_150),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_65),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_192),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_55),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_54),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_74),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_16),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_174),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_159),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_6),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_36),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_60),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_4),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_129),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_104),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_67),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_135),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_5),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_29),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_34),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_79),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_64),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_173),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_5),
.Y(n_373)
);

INVx2_ASAP7_75t_R g374 ( 
.A(n_115),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_65),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_200),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_36),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_31),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_113),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_145),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_165),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_19),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_201),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_26),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_18),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_7),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_176),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_112),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_105),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_76),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_79),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_21),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_181),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_84),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_50),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_48),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_187),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_141),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_31),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_72),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_134),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_118),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_260),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_218),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_218),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_218),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_366),
.B(n_0),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_218),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_203),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_245),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_204),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_205),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_207),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_211),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_212),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_397),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_234),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_380),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_214),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_245),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_366),
.B(n_0),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_218),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_380),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_206),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_215),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_234),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_216),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_250),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_280),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_250),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_337),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_218),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_219),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_221),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_224),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_208),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_294),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_225),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_294),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_368),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_R g443 ( 
.A(n_231),
.B(n_95),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_233),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_236),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_294),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_294),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_294),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_238),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_294),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_241),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_313),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_251),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_313),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_253),
.Y(n_455)
);

INVxp33_ASAP7_75t_SL g456 ( 
.A(n_368),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_254),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_313),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_257),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_259),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_332),
.B(n_3),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_313),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_313),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_264),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_249),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_332),
.B(n_220),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_267),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_313),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_268),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_269),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_280),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_351),
.Y(n_472)
);

BUFx2_ASAP7_75t_SL g473 ( 
.A(n_242),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_222),
.B(n_3),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_220),
.B(n_8),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_270),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_351),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_274),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_337),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_276),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_279),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_281),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_284),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_208),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_285),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_337),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_302),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_242),
.B(n_8),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_351),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_302),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_290),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_351),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_351),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_351),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_222),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_292),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_382),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_319),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_382),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_382),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_382),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_382),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_230),
.B(n_10),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_319),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_295),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_229),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_209),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_297),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_308),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_298),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_311),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_312),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g514 ( 
.A(n_344),
.B(n_10),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_298),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_314),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_329),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_329),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_315),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_410),
.Y(n_520)
);

INVxp33_ASAP7_75t_SL g521 ( 
.A(n_412),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_413),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_430),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_414),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_463),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_415),
.B(n_416),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_463),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_463),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_404),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_404),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_411),
.B(n_328),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_403),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_406),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_406),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_420),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_407),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_407),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_409),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_438),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_426),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_409),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_498),
.B(n_255),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_442),
.A2(n_275),
.B1(n_278),
.B2(n_261),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_423),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_R g546 ( 
.A(n_425),
.B(n_317),
.Y(n_546)
);

NOR2xp67_ASAP7_75t_L g547 ( 
.A(n_433),
.B(n_358),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_433),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_428),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_432),
.B(n_210),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_466),
.B(n_320),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_439),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_439),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_487),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_435),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_441),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_441),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_490),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_446),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_446),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_479),
.B(n_210),
.Y(n_561)
);

CKINVDCx16_ASAP7_75t_R g562 ( 
.A(n_437),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_436),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_447),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_447),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_411),
.B(n_328),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_440),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_405),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_450),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_438),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_450),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_486),
.B(n_322),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_452),
.Y(n_574)
);

CKINVDCx16_ASAP7_75t_R g575 ( 
.A(n_437),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_452),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_430),
.B(n_228),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_444),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_445),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_454),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_454),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_458),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_458),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_430),
.B(n_228),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_462),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_462),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_468),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_468),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_449),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_472),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_472),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_477),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_477),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_489),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_430),
.B(n_471),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_419),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g597 ( 
.A(n_484),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_489),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_417),
.Y(n_599)
);

NAND2x1_ASAP7_75t_L g600 ( 
.A(n_492),
.B(n_246),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_451),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_455),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_492),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_493),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_494),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_505),
.B(n_255),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_494),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_434),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_457),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_497),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_551),
.B(n_464),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_539),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_523),
.Y(n_614)
);

AND2x2_ASAP7_75t_SL g615 ( 
.A(n_562),
.B(n_408),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_550),
.B(n_561),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_595),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_539),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_554),
.B(n_484),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_554),
.B(n_465),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_573),
.A2(n_461),
.B1(n_422),
.B2(n_456),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_541),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_542),
.A2(n_459),
.B1(n_460),
.B2(n_453),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_558),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_550),
.B(n_246),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_539),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_550),
.A2(n_561),
.B1(n_418),
.B2(n_504),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_573),
.A2(n_467),
.B1(n_481),
.B2(n_480),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_523),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_577),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_541),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_544),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_550),
.B(n_469),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_561),
.B(n_470),
.Y(n_634)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_523),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_577),
.Y(n_636)
);

AND2x2_ASAP7_75t_SL g637 ( 
.A(n_562),
.B(n_475),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_577),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_577),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_584),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_544),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_584),
.Y(n_642)
);

INVx6_ASAP7_75t_L g643 ( 
.A(n_584),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_539),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_561),
.B(n_421),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_548),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_584),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_525),
.Y(n_648)
);

BUFx8_ASAP7_75t_SL g649 ( 
.A(n_532),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_607),
.A2(n_325),
.B1(n_384),
.B2(n_213),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_548),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_520),
.B(n_363),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_539),
.Y(n_653)
);

INVx4_ASAP7_75t_SL g654 ( 
.A(n_539),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_525),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_558),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_527),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_527),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_546),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_528),
.Y(n_660)
);

BUFx10_ASAP7_75t_L g661 ( 
.A(n_526),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_548),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_531),
.B(n_363),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_522),
.B(n_476),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_528),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_547),
.B(n_478),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_571),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_571),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_L g669 ( 
.A(n_543),
.B(n_424),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_571),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_547),
.B(n_482),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_529),
.B(n_483),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_531),
.A2(n_427),
.B1(n_374),
.B2(n_429),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_529),
.B(n_485),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_567),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_530),
.Y(n_676)
);

NAND2x1p5_ASAP7_75t_L g677 ( 
.A(n_600),
.B(n_398),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_552),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_521),
.B(n_496),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_567),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_524),
.B(n_506),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_536),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_537),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_535),
.A2(n_491),
.B1(n_510),
.B2(n_509),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_540),
.B(n_512),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_537),
.B(n_421),
.Y(n_686)
);

INVx4_ASAP7_75t_SL g687 ( 
.A(n_571),
.Y(n_687)
);

INVxp67_ASAP7_75t_SL g688 ( 
.A(n_571),
.Y(n_688)
);

AO21x2_ASAP7_75t_L g689 ( 
.A1(n_538),
.A2(n_232),
.B(n_230),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_538),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_553),
.B(n_473),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_549),
.B(n_513),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_575),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_553),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_555),
.B(n_516),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_571),
.B(n_232),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_600),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_533),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_556),
.B(n_519),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_563),
.B(n_568),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_552),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_578),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_552),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_579),
.B(n_248),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_543),
.B(n_508),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_556),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_557),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_589),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_557),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_596),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_559),
.B(n_430),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_559),
.B(n_473),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_575),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_560),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_533),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_560),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_601),
.B(n_248),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_564),
.B(n_471),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_564),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_533),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_602),
.B(n_252),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_566),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_533),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_566),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_569),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_565),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_572),
.B(n_471),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_534),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_610),
.B(n_252),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_565),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_597),
.B(n_431),
.C(n_427),
.Y(n_731)
);

INVx5_ASAP7_75t_L g732 ( 
.A(n_534),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_597),
.B(n_471),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_576),
.A2(n_374),
.B1(n_474),
.B2(n_344),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_580),
.B(n_581),
.Y(n_735)
);

INVx5_ASAP7_75t_L g736 ( 
.A(n_534),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_580),
.B(n_383),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_581),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_534),
.Y(n_739)
);

AND2x2_ASAP7_75t_SL g740 ( 
.A(n_596),
.B(n_262),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_585),
.B(n_495),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_585),
.B(n_499),
.Y(n_742)
);

INVx5_ASAP7_75t_L g743 ( 
.A(n_545),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_565),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_545),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_586),
.B(n_507),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_586),
.B(n_474),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_588),
.B(n_499),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_545),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_591),
.B(n_262),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_591),
.A2(n_514),
.B1(n_488),
.B2(n_223),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_545),
.Y(n_752)
);

AND2x6_ASAP7_75t_L g753 ( 
.A(n_598),
.B(n_271),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_603),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_583),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_606),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_583),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_583),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_606),
.B(n_229),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_570),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_621),
.A2(n_616),
.B1(n_634),
.B2(n_633),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_705),
.A2(n_354),
.B1(n_341),
.B2(n_266),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_639),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_616),
.B(n_608),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_689),
.A2(n_374),
.B1(n_354),
.B2(n_341),
.Y(n_765)
);

OAI221xp5_ASAP7_75t_L g766 ( 
.A1(n_673),
.A2(n_627),
.B1(n_734),
.B2(n_747),
.C(n_759),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_616),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_638),
.B(n_383),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_638),
.B(n_383),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_630),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_622),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_620),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_612),
.B(n_608),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_620),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_675),
.B(n_609),
.Y(n_775)
);

AOI22x1_ASAP7_75t_L g776 ( 
.A1(n_617),
.A2(n_299),
.B1(n_300),
.B2(n_271),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_649),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_675),
.B(n_443),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_636),
.A2(n_300),
.B(n_303),
.C(n_299),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_639),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_680),
.B(n_217),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_622),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_649),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_640),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_631),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_631),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_642),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_645),
.B(n_304),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_632),
.Y(n_789)
);

OR2x6_ASAP7_75t_L g790 ( 
.A(n_713),
.B(n_235),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_647),
.Y(n_791)
);

NOR3xp33_ASAP7_75t_L g792 ( 
.A(n_650),
.B(n_227),
.C(n_226),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_686),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_680),
.B(n_237),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_725),
.Y(n_795)
);

INVx8_ASAP7_75t_L g796 ( 
.A(n_663),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_637),
.A2(n_645),
.B1(n_733),
.B2(n_674),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_672),
.B(n_239),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_714),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_699),
.B(n_240),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_632),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_714),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_759),
.B(n_303),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_756),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_756),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_638),
.B(n_383),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_691),
.B(n_712),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_635),
.A2(n_611),
.B(n_574),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_715),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_676),
.B(n_583),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_715),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_656),
.B(n_304),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_625),
.A2(n_503),
.B(n_502),
.C(n_501),
.Y(n_813)
);

O2A1O1Ixp5_ASAP7_75t_L g814 ( 
.A1(n_750),
.A2(n_605),
.B(n_381),
.C(n_387),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_682),
.B(n_605),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_683),
.B(n_605),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_679),
.B(n_335),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_690),
.B(n_605),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_694),
.B(n_305),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_619),
.B(n_656),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_720),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_643),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_659),
.B(n_304),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_704),
.B(n_243),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_L g825 ( 
.A(n_628),
.B(n_247),
.C(n_244),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_704),
.B(n_256),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_706),
.B(n_305),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_624),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_725),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_740),
.B(n_373),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_638),
.B(n_383),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_720),
.B(n_383),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_707),
.B(n_306),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_709),
.B(n_306),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_716),
.B(n_323),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_719),
.B(n_323),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_759),
.B(n_330),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_629),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_723),
.Y(n_839)
);

BUFx6f_ASAP7_75t_SL g840 ( 
.A(n_702),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_723),
.B(n_383),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_740),
.A2(n_394),
.B1(n_372),
.B2(n_388),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_717),
.B(n_263),
.C(n_258),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_717),
.B(n_265),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_723),
.B(n_383),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_721),
.B(n_272),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_689),
.A2(n_296),
.B1(n_266),
.B2(n_377),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_722),
.B(n_330),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_689),
.A2(n_296),
.B1(n_377),
.B2(n_235),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_721),
.A2(n_357),
.B1(n_364),
.B2(n_376),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_741),
.B(n_373),
.Y(n_851)
);

AND2x6_ASAP7_75t_L g852 ( 
.A(n_697),
.B(n_728),
.Y(n_852)
);

INVx5_ASAP7_75t_L g853 ( 
.A(n_663),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_728),
.Y(n_854)
);

NAND3xp33_ASAP7_75t_L g855 ( 
.A(n_729),
.B(n_652),
.C(n_746),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_724),
.B(n_352),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_729),
.B(n_273),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_619),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_705),
.B(n_277),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_713),
.B(n_373),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_641),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_750),
.A2(n_500),
.B(n_291),
.C(n_327),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_641),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_728),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_693),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_646),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_738),
.B(n_381),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_643),
.A2(n_387),
.B1(n_402),
.B2(n_401),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_754),
.B(n_402),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_749),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_648),
.A2(n_291),
.B(n_327),
.C(n_339),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_753),
.A2(n_378),
.B1(n_355),
.B2(n_339),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_615),
.A2(n_350),
.B1(n_379),
.B2(n_336),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_655),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_657),
.B(n_570),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_666),
.B(n_671),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_664),
.B(n_282),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_658),
.A2(n_378),
.B(n_355),
.C(n_342),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_660),
.B(n_574),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_664),
.B(n_283),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_665),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_646),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_752),
.B(n_643),
.Y(n_883)
);

NOR2xp67_ASAP7_75t_SL g884 ( 
.A(n_643),
.B(n_342),
.Y(n_884)
);

OAI221xp5_ASAP7_75t_L g885 ( 
.A1(n_759),
.A2(n_365),
.B1(n_286),
.B2(n_287),
.C(n_288),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_615),
.A2(n_393),
.B1(n_389),
.B2(n_347),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_684),
.B(n_338),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_661),
.B(n_343),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_751),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_688),
.A2(n_604),
.B(n_574),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_661),
.B(n_346),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_681),
.B(n_289),
.Y(n_892)
);

AO221x1_ASAP7_75t_L g893 ( 
.A1(n_614),
.A2(n_255),
.B1(n_511),
.B2(n_517),
.C(n_515),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_698),
.B(n_255),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_735),
.B(n_604),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_681),
.B(n_293),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_698),
.B(n_582),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_663),
.A2(n_371),
.B1(n_369),
.B2(n_386),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_731),
.B(n_301),
.Y(n_899)
);

NOR2xp67_ASAP7_75t_L g900 ( 
.A(n_623),
.B(n_98),
.Y(n_900)
);

AND2x6_ASAP7_75t_SL g901 ( 
.A(n_669),
.B(n_511),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_702),
.B(n_373),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_753),
.A2(n_391),
.B1(n_395),
.B2(n_396),
.Y(n_903)
);

BUFx6f_ASAP7_75t_SL g904 ( 
.A(n_702),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_739),
.B(n_745),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_711),
.A2(n_590),
.B(n_594),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_883),
.A2(n_668),
.B(n_613),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_774),
.B(n_661),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_767),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_865),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_770),
.Y(n_911)
);

INVx3_ASAP7_75t_SL g912 ( 
.A(n_829),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_772),
.B(n_710),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_853),
.A2(n_667),
.B(n_653),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_763),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_763),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_807),
.B(n_739),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_824),
.B(n_669),
.C(n_685),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_784),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_820),
.B(n_710),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_797),
.B(n_708),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_761),
.B(n_708),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_765),
.A2(n_737),
.B(n_663),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_876),
.A2(n_663),
.B1(n_692),
.B2(n_685),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_828),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_798),
.B(n_800),
.Y(n_926)
);

AND2x2_ASAP7_75t_SL g927 ( 
.A(n_903),
.B(n_708),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_765),
.A2(n_662),
.B(n_651),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_L g929 ( 
.A(n_826),
.B(n_695),
.C(n_700),
.Y(n_929)
);

NAND2xp33_ASAP7_75t_L g930 ( 
.A(n_852),
.B(n_677),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_876),
.B(n_677),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_773),
.B(n_739),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_798),
.B(n_599),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_775),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_787),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_764),
.A2(n_614),
.B(n_618),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_783),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_791),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_800),
.B(n_614),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_809),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_855),
.B(n_763),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_905),
.A2(n_748),
.B(n_742),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_905),
.A2(n_614),
.B(n_618),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_851),
.B(n_375),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_812),
.B(n_375),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_895),
.A2(n_670),
.B(n_626),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_811),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_844),
.A2(n_718),
.B(n_727),
.C(n_670),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_780),
.B(n_755),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_796),
.A2(n_644),
.B(n_732),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_828),
.B(n_755),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_766),
.A2(n_760),
.B(n_662),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_796),
.A2(n_644),
.B(n_732),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_846),
.A2(n_760),
.B(n_730),
.C(n_726),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_796),
.A2(n_644),
.B(n_732),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_780),
.B(n_755),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_822),
.A2(n_736),
.B(n_743),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_842),
.B(n_678),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_874),
.B(n_757),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_822),
.A2(n_736),
.B(n_743),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_847),
.A2(n_390),
.B1(n_309),
.B2(n_310),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_780),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_793),
.B(n_654),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_881),
.B(n_757),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_799),
.B(n_757),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_810),
.A2(n_736),
.B(n_743),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_815),
.A2(n_757),
.B(n_758),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_816),
.A2(n_758),
.B(n_701),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_SL g969 ( 
.A(n_840),
.B(n_375),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_780),
.B(n_758),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_847),
.A2(n_385),
.B1(n_316),
.B2(n_318),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_877),
.B(n_758),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_846),
.A2(n_678),
.B(n_744),
.C(n_726),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_818),
.A2(n_701),
.B(n_703),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_768),
.A2(n_592),
.B(n_587),
.Y(n_975)
);

OAI21xp33_ASAP7_75t_L g976 ( 
.A1(n_857),
.A2(n_367),
.B(n_321),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_830),
.B(n_307),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_849),
.A2(n_753),
.B(n_696),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_802),
.B(n_804),
.Y(n_979)
);

OAI321xp33_ASAP7_75t_L g980 ( 
.A1(n_762),
.A2(n_518),
.A3(n_517),
.B1(n_515),
.B2(n_375),
.C(n_594),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_858),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_805),
.B(n_753),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_821),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_838),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_857),
.A2(n_370),
.B(n_326),
.C(n_331),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_769),
.A2(n_593),
.B(n_587),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_769),
.A2(n_594),
.B(n_590),
.Y(n_987)
);

AND2x6_ASAP7_75t_L g988 ( 
.A(n_803),
.B(n_837),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_806),
.A2(n_593),
.B(n_590),
.Y(n_989)
);

OAI321xp33_ASAP7_75t_L g990 ( 
.A1(n_762),
.A2(n_518),
.A3(n_333),
.B1(n_334),
.B2(n_340),
.C(n_345),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_877),
.A2(n_753),
.B1(n_696),
.B2(n_687),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_788),
.B(n_324),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_790),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_839),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_854),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_864),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_838),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_831),
.A2(n_687),
.B(n_654),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_831),
.A2(n_687),
.B(n_654),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_880),
.B(n_892),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_849),
.A2(n_348),
.B1(n_353),
.B2(n_356),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_880),
.B(n_359),
.Y(n_1002)
);

AND2x6_ASAP7_75t_L g1003 ( 
.A(n_803),
.B(n_696),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_896),
.A2(n_392),
.B(n_400),
.C(n_399),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_795),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_790),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_777),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_859),
.B(n_360),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_781),
.A2(n_362),
.B(n_361),
.C(n_14),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_903),
.A2(n_872),
.B1(n_898),
.B2(n_889),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_870),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_832),
.A2(n_845),
.B(n_841),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_852),
.B(n_99),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_823),
.B(n_12),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_781),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_794),
.B(n_15),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_900),
.B(n_902),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_838),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_832),
.A2(n_199),
.B(n_191),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_794),
.B(n_852),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_897),
.A2(n_879),
.B(n_875),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_808),
.A2(n_183),
.B(n_179),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_838),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_790),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_852),
.B(n_17),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_837),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_894),
.A2(n_172),
.B1(n_171),
.B2(n_164),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_771),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_817),
.B(n_24),
.Y(n_1029)
);

INVxp67_ASAP7_75t_SL g1030 ( 
.A(n_782),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_843),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_819),
.B(n_28),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_890),
.A2(n_146),
.B(n_143),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_873),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_825),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_899),
.B(n_38),
.Y(n_1036)
);

AOI21x1_ASAP7_75t_L g1037 ( 
.A1(n_906),
.A2(n_137),
.B(n_132),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_778),
.A2(n_130),
.B(n_128),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_894),
.A2(n_125),
.B1(n_122),
.B2(n_121),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_901),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_827),
.B(n_833),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_779),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_860),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_785),
.A2(n_107),
.B(n_43),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_814),
.A2(n_41),
.B(n_46),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_786),
.A2(n_46),
.B(n_47),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_789),
.A2(n_47),
.B(n_49),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_801),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_834),
.B(n_50),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_886),
.B(n_53),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_835),
.B(n_53),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_861),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_887),
.B(n_54),
.C(n_55),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_863),
.A2(n_56),
.B(n_59),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_866),
.B(n_60),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_888),
.B(n_63),
.Y(n_1056)
);

NOR3xp33_ASAP7_75t_L g1057 ( 
.A(n_891),
.B(n_63),
.C(n_64),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_850),
.B(n_66),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_882),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_836),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_848),
.A2(n_67),
.B(n_68),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_856),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_1000),
.B(n_926),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_911),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_930),
.A2(n_872),
.B(n_867),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_923),
.A2(n_939),
.B(n_931),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1002),
.B(n_1060),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_934),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_907),
.A2(n_869),
.B(n_813),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_SL g1070 ( 
.A1(n_1019),
.A2(n_862),
.B(n_776),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1062),
.B(n_792),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_977),
.B(n_868),
.Y(n_1072)
);

INVx6_ASAP7_75t_SL g1073 ( 
.A(n_963),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_912),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_915),
.B(n_884),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_968),
.A2(n_893),
.B(n_878),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1041),
.B(n_885),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_932),
.A2(n_871),
.B(n_904),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_R g1079 ( 
.A(n_1040),
.B(n_904),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_952),
.A2(n_840),
.B(n_70),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_918),
.A2(n_83),
.B1(n_70),
.B2(n_76),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_919),
.B(n_935),
.Y(n_1082)
);

AOI221x1_ASAP7_75t_L g1083 ( 
.A1(n_1016),
.A2(n_68),
.B1(n_77),
.B2(n_80),
.C(n_81),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_910),
.Y(n_1084)
);

BUFx4f_ASAP7_75t_L g1085 ( 
.A(n_1026),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_936),
.A2(n_77),
.B(n_1021),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_943),
.A2(n_967),
.B(n_942),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_1050),
.A2(n_1010),
.B(n_1029),
.C(n_1056),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1020),
.A2(n_972),
.B(n_917),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_920),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_1008),
.B(n_925),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_940),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_938),
.B(n_944),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_SL g1094 ( 
.A1(n_1010),
.A2(n_971),
.B1(n_961),
.B2(n_1001),
.C(n_976),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_929),
.A2(n_1014),
.B(n_924),
.C(n_990),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_927),
.A2(n_922),
.B1(n_921),
.B2(n_933),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_992),
.B(n_1043),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_913),
.B(n_908),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_954),
.A2(n_973),
.A3(n_948),
.B(n_1015),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_945),
.B(n_1005),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1026),
.B(n_909),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_928),
.A2(n_1012),
.B(n_914),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1036),
.B(n_979),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_SL g1104 ( 
.A1(n_1019),
.A2(n_1038),
.B(n_1013),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_SL g1105 ( 
.A1(n_978),
.A2(n_1013),
.B(n_991),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_916),
.B(n_962),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_978),
.A2(n_970),
.B(n_949),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_916),
.B(n_962),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_SL g1109 ( 
.A1(n_1025),
.A2(n_1032),
.B(n_1049),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_951),
.B(n_988),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_981),
.Y(n_1111)
);

INVx6_ASAP7_75t_L g1112 ( 
.A(n_984),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_956),
.A2(n_941),
.B(n_982),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1059),
.Y(n_1114)
);

O2A1O1Ixp5_ASAP7_75t_L g1115 ( 
.A1(n_1037),
.A2(n_1022),
.B(n_1045),
.C(n_1051),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_990),
.A2(n_1009),
.B(n_1034),
.C(n_1058),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1028),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_984),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1052),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1030),
.A2(n_959),
.B(n_964),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_958),
.A2(n_998),
.B(n_999),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1053),
.A2(n_1035),
.B(n_1057),
.C(n_980),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_988),
.B(n_997),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_SL g1124 ( 
.A1(n_969),
.A2(n_1001),
.B1(n_971),
.B2(n_961),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_947),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_1031),
.A2(n_1055),
.A3(n_1004),
.B(n_985),
.Y(n_1126)
);

AO21x1_ASAP7_75t_L g1127 ( 
.A1(n_1045),
.A2(n_1017),
.B(n_1055),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_983),
.A2(n_1011),
.B(n_994),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1026),
.B(n_915),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_988),
.B(n_997),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_950),
.A2(n_955),
.B(n_953),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_975),
.A2(n_987),
.B(n_986),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_995),
.A2(n_996),
.B1(n_916),
.B2(n_962),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_988),
.B(n_1018),
.Y(n_1134)
);

NOR2x1_ASAP7_75t_SL g1135 ( 
.A(n_984),
.B(n_1018),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_965),
.A2(n_966),
.B(n_989),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_963),
.A2(n_957),
.B(n_960),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1033),
.A2(n_1023),
.B(n_1018),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_1023),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1023),
.B(n_1048),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1048),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_993),
.B(n_1006),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1048),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1024),
.B(n_1003),
.Y(n_1144)
);

AOI221x1_ASAP7_75t_L g1145 ( 
.A1(n_1061),
.A2(n_1054),
.B1(n_1047),
.B2(n_1046),
.C(n_1044),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1027),
.A2(n_1039),
.B(n_980),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1042),
.A2(n_1003),
.B(n_1007),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1003),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1003),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_937),
.A2(n_907),
.B(n_946),
.Y(n_1150)
);

NAND2x1p5_ASAP7_75t_L g1151 ( 
.A(n_915),
.B(n_916),
.Y(n_1151)
);

OAI22x1_ASAP7_75t_L g1152 ( 
.A1(n_1000),
.A2(n_669),
.B1(n_918),
.B2(n_926),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_926),
.B(n_1000),
.Y(n_1153)
);

AO21x1_ASAP7_75t_L g1154 ( 
.A1(n_1000),
.A2(n_926),
.B(n_1002),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_930),
.A2(n_853),
.B(n_923),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_920),
.Y(n_1156)
);

O2A1O1Ixp5_ASAP7_75t_L g1157 ( 
.A1(n_926),
.A2(n_1000),
.B(n_1002),
.C(n_1016),
.Y(n_1157)
);

NOR2x1_ASAP7_75t_L g1158 ( 
.A(n_929),
.B(n_1017),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_920),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_912),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_907),
.A2(n_946),
.B(n_974),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_930),
.A2(n_853),
.B(n_923),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_911),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_916),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_930),
.A2(n_853),
.B(n_923),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_907),
.A2(n_946),
.B(n_974),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_926),
.B(n_1000),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_907),
.A2(n_946),
.B(n_974),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_920),
.B(n_820),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1000),
.A2(n_926),
.B(n_1050),
.C(n_1002),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_926),
.A2(n_1000),
.B(n_952),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_940),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_945),
.B(n_772),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1000),
.B(n_926),
.C(n_1002),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_945),
.B(n_772),
.Y(n_1175)
);

O2A1O1Ixp5_ASAP7_75t_L g1176 ( 
.A1(n_926),
.A2(n_1000),
.B(n_1002),
.C(n_1016),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_SL g1177 ( 
.A1(n_1019),
.A2(n_1038),
.B(n_1013),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_911),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_926),
.A2(n_1000),
.B(n_952),
.Y(n_1179)
);

AOI221x1_ASAP7_75t_L g1180 ( 
.A1(n_1000),
.A2(n_926),
.B1(n_1002),
.B2(n_1016),
.C(n_931),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1000),
.B(n_926),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1026),
.B(n_911),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_926),
.B(n_1000),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_945),
.B(n_772),
.Y(n_1184)
);

OAI22x1_ASAP7_75t_L g1185 ( 
.A1(n_1000),
.A2(n_669),
.B1(n_918),
.B2(n_926),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_984),
.Y(n_1186)
);

OAI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_926),
.A2(n_1000),
.B(n_1002),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1000),
.A2(n_762),
.B1(n_621),
.B2(n_650),
.C(n_1010),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_926),
.B(n_1000),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_930),
.A2(n_853),
.B(n_923),
.Y(n_1190)
);

AO21x1_ASAP7_75t_L g1191 ( 
.A1(n_1000),
.A2(n_926),
.B(n_1002),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_920),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_926),
.B(n_1000),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_930),
.A2(n_853),
.B(n_923),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_934),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1026),
.B(n_911),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1000),
.B(n_926),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1000),
.B(n_926),
.Y(n_1198)
);

OAI22x1_ASAP7_75t_L g1199 ( 
.A1(n_1000),
.A2(n_669),
.B1(n_918),
.B2(n_926),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_926),
.B(n_1000),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_926),
.B(n_1000),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_945),
.B(n_772),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_981),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_952),
.A2(n_1037),
.B(n_1022),
.Y(n_1204)
);

AOI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_1000),
.A2(n_926),
.B(n_1002),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1092),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1063),
.A2(n_1197),
.B1(n_1198),
.B2(n_1174),
.Y(n_1207)
);

INVx5_ASAP7_75t_L g1208 ( 
.A(n_1118),
.Y(n_1208)
);

AND2x2_ASAP7_75t_SL g1209 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_1085),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1198),
.A2(n_1174),
.B1(n_1187),
.B2(n_1205),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_1074),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1169),
.B(n_1159),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1153),
.B(n_1167),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1183),
.B(n_1189),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1090),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1084),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1125),
.Y(n_1218)
);

OR2x6_ASAP7_75t_L g1219 ( 
.A(n_1090),
.B(n_1129),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1101),
.B(n_1182),
.Y(n_1220)
);

BUFx8_ASAP7_75t_SL g1221 ( 
.A(n_1074),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1192),
.B(n_1193),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1160),
.Y(n_1223)
);

INVx5_ASAP7_75t_L g1224 ( 
.A(n_1118),
.Y(n_1224)
);

CKINVDCx6p67_ASAP7_75t_R g1225 ( 
.A(n_1084),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1068),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1155),
.A2(n_1165),
.B(n_1162),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1118),
.Y(n_1228)
);

NOR2x1_ASAP7_75t_SL g1229 ( 
.A(n_1133),
.B(n_1110),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1101),
.B(n_1182),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1082),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1118),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1160),
.Y(n_1233)
);

INVxp67_ASAP7_75t_SL g1234 ( 
.A(n_1200),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1195),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1201),
.A2(n_1170),
.B1(n_1088),
.B2(n_1171),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1156),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1190),
.A2(n_1194),
.B(n_1066),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1181),
.B(n_1170),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1181),
.B(n_1067),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1088),
.A2(n_1179),
.B1(n_1124),
.B2(n_1188),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1103),
.B(n_1098),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1073),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1203),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1114),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_1100),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1139),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1129),
.B(n_1134),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1157),
.A2(n_1176),
.B(n_1095),
.Y(n_1249)
);

INVx8_ASAP7_75t_L g1250 ( 
.A(n_1139),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1077),
.B(n_1094),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1204),
.A2(n_1115),
.B(n_1086),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1154),
.B(n_1191),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1142),
.Y(n_1254)
);

NAND2x1_ASAP7_75t_L g1255 ( 
.A(n_1186),
.B(n_1129),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1064),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1111),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1180),
.B(n_1096),
.Y(n_1258)
);

BUFx10_ASAP7_75t_L g1259 ( 
.A(n_1098),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1124),
.A2(n_1072),
.B1(n_1122),
.B2(n_1095),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1103),
.B(n_1071),
.Y(n_1261)
);

NAND3xp33_ASAP7_75t_L g1262 ( 
.A(n_1157),
.B(n_1176),
.C(n_1080),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1139),
.Y(n_1263)
);

BUFx5_ASAP7_75t_L g1264 ( 
.A(n_1149),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1146),
.A2(n_1116),
.B(n_1122),
.C(n_1065),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1116),
.A2(n_1097),
.B(n_1093),
.C(n_1091),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1163),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1173),
.B(n_1175),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1184),
.B(n_1202),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1152),
.B(n_1185),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1182),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1105),
.A2(n_1089),
.B(n_1177),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1178),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1081),
.A2(n_1085),
.B1(n_1158),
.B2(n_1128),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1104),
.A2(n_1120),
.B(n_1121),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1112),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1199),
.B(n_1196),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1144),
.B(n_1196),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1073),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1138),
.A2(n_1131),
.B(n_1107),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1131),
.A2(n_1113),
.B(n_1137),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1196),
.B(n_1101),
.Y(n_1282)
);

INVxp67_ASAP7_75t_SL g1283 ( 
.A(n_1164),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1117),
.B(n_1119),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1172),
.B(n_1141),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1073),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1078),
.A2(n_1070),
.B(n_1127),
.C(n_1143),
.Y(n_1287)
);

A2O1A1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1150),
.A2(n_1147),
.B(n_1076),
.C(n_1102),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1139),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1112),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1164),
.A2(n_1148),
.B1(n_1075),
.B2(n_1141),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_SL g1292 ( 
.A1(n_1148),
.A2(n_1130),
.B(n_1123),
.C(n_1140),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_1186),
.B(n_1135),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1112),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1151),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1126),
.B(n_1106),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1106),
.B(n_1108),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1126),
.B(n_1151),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1108),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1075),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1079),
.B(n_1136),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1126),
.B(n_1099),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1161),
.A2(n_1168),
.B(n_1166),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1087),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1109),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1083),
.A2(n_1126),
.B1(n_1109),
.B2(n_1145),
.Y(n_1306)
);

CKINVDCx6p67_ASAP7_75t_R g1307 ( 
.A(n_1099),
.Y(n_1307)
);

BUFx12f_ASAP7_75t_L g1308 ( 
.A(n_1099),
.Y(n_1308)
);

BUFx4f_ASAP7_75t_L g1309 ( 
.A(n_1099),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1069),
.Y(n_1310)
);

OAI321xp33_ASAP7_75t_L g1311 ( 
.A1(n_1132),
.A2(n_1198),
.A3(n_1063),
.B1(n_1197),
.B2(n_1187),
.C(n_1167),
.Y(n_1311)
);

AND2x2_ASAP7_75t_SL g1312 ( 
.A(n_1063),
.B(n_927),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1125),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1073),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_SL g1315 ( 
.A(n_1170),
.B(n_1000),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1317)
);

BUFx12f_ASAP7_75t_L g1318 ( 
.A(n_1074),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1124),
.A2(n_1063),
.B1(n_1198),
.B2(n_1197),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1321)
);

AOI222xp33_ASAP7_75t_L g1322 ( 
.A1(n_1063),
.A2(n_1197),
.B1(n_1198),
.B2(n_1188),
.C1(n_1174),
.C2(n_1187),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1155),
.A2(n_1165),
.B(n_1162),
.Y(n_1323)
);

O2A1O1Ixp5_ASAP7_75t_L g1324 ( 
.A1(n_1205),
.A2(n_926),
.B(n_1000),
.C(n_1170),
.Y(n_1324)
);

INVx6_ASAP7_75t_L g1325 ( 
.A(n_1090),
.Y(n_1325)
);

INVx3_ASAP7_75t_SL g1326 ( 
.A(n_1074),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1084),
.Y(n_1327)
);

CKINVDCx8_ASAP7_75t_R g1328 ( 
.A(n_1074),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1118),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_SL g1330 ( 
.A(n_1170),
.B(n_1000),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1174),
.A2(n_1000),
.B1(n_926),
.B2(n_1205),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1084),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1159),
.Y(n_1333)
);

NAND3xp33_ASAP7_75t_L g1334 ( 
.A(n_1205),
.B(n_1000),
.C(n_926),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1084),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1092),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1159),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1159),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1342)
);

OAI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1063),
.A2(n_1198),
.B(n_1197),
.Y(n_1343)
);

O2A1O1Ixp5_ASAP7_75t_SL g1344 ( 
.A1(n_1205),
.A2(n_1080),
.B(n_1181),
.C(n_1179),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1159),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1205),
.B(n_1000),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1169),
.Y(n_1348)
);

BUFx4_ASAP7_75t_SL g1349 ( 
.A(n_1074),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1063),
.A2(n_1198),
.B1(n_1197),
.B2(n_1167),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1068),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1155),
.A2(n_1165),
.B(n_1162),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1068),
.Y(n_1355)
);

NAND2x1p5_ASAP7_75t_L g1356 ( 
.A(n_1085),
.B(n_915),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1068),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1118),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1063),
.B(n_1197),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1169),
.B(n_1159),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_L g1361 ( 
.A1(n_1205),
.A2(n_926),
.B(n_1000),
.C(n_1170),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1084),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1159),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1298),
.B(n_1309),
.Y(n_1364)
);

NAND2x1p5_ASAP7_75t_L g1365 ( 
.A(n_1309),
.B(n_1310),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1308),
.B(n_1241),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1218),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1319),
.A2(n_1312),
.B1(n_1330),
.B2(n_1315),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1327),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1313),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1332),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1220),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_SL g1373 ( 
.A1(n_1229),
.A2(n_1287),
.B(n_1239),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1283),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1220),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1257),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1207),
.A2(n_1334),
.B1(n_1330),
.B2(n_1315),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1242),
.B(n_1234),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1208),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1226),
.Y(n_1380)
);

INVx6_ASAP7_75t_L g1381 ( 
.A(n_1210),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1322),
.A2(n_1331),
.B1(n_1343),
.B2(n_1241),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1209),
.A2(n_1350),
.B1(n_1260),
.B2(n_1236),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1230),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1245),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1225),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1230),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1322),
.A2(n_1260),
.B1(n_1347),
.B2(n_1236),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1333),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1275),
.A2(n_1281),
.B(n_1272),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1353),
.A2(n_1359),
.B1(n_1335),
.B2(n_1320),
.Y(n_1391)
);

BUFx12f_ASAP7_75t_L g1392 ( 
.A(n_1216),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1350),
.A2(n_1270),
.B1(n_1211),
.B2(n_1274),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1256),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1214),
.B(n_1317),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1267),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1273),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1244),
.Y(n_1398)
);

NOR2x1_ASAP7_75t_R g1399 ( 
.A(n_1233),
.B(n_1212),
.Y(n_1399)
);

INVx4_ASAP7_75t_SL g1400 ( 
.A(n_1300),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1336),
.B(n_1340),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1274),
.A2(n_1277),
.B1(n_1261),
.B2(n_1321),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1208),
.Y(n_1403)
);

CKINVDCx16_ASAP7_75t_R g1404 ( 
.A(n_1223),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1338),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1299),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1316),
.A2(n_1345),
.B1(n_1320),
.B2(n_1351),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1208),
.Y(n_1408)
);

AOI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1306),
.A2(n_1280),
.B(n_1323),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1264),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1208),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1324),
.A2(n_1361),
.B(n_1344),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1261),
.A2(n_1316),
.B1(n_1351),
.B2(n_1335),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1333),
.Y(n_1414)
);

BUFx12f_ASAP7_75t_L g1415 ( 
.A(n_1318),
.Y(n_1415)
);

INVx4_ASAP7_75t_L g1416 ( 
.A(n_1224),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1302),
.B(n_1240),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1321),
.B(n_1342),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1224),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1264),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1345),
.A2(n_1359),
.B1(n_1259),
.B2(n_1262),
.Y(n_1421)
);

BUFx2_ASAP7_75t_R g1422 ( 
.A(n_1221),
.Y(n_1422)
);

AO21x1_ASAP7_75t_SL g1423 ( 
.A1(n_1253),
.A2(n_1296),
.B(n_1258),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1278),
.B(n_1251),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1259),
.A2(n_1215),
.B1(n_1325),
.B2(n_1258),
.Y(n_1425)
);

BUFx2_ASAP7_75t_R g1426 ( 
.A(n_1328),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1284),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1231),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1326),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1224),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1249),
.A2(n_1238),
.B(n_1265),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1285),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1222),
.A2(n_1246),
.B1(n_1268),
.B2(n_1348),
.Y(n_1433)
);

CKINVDCx11_ASAP7_75t_R g1434 ( 
.A(n_1219),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1251),
.A2(n_1266),
.B(n_1253),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1237),
.Y(n_1436)
);

OAI22x1_ASAP7_75t_L g1437 ( 
.A1(n_1305),
.A2(n_1301),
.B1(n_1246),
.B2(n_1296),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1311),
.B(n_1300),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1269),
.A2(n_1307),
.B1(n_1213),
.B2(n_1360),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1289),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1248),
.B(n_1271),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1297),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1248),
.B(n_1282),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1228),
.Y(n_1444)
);

INVx4_ASAP7_75t_L g1445 ( 
.A(n_1224),
.Y(n_1445)
);

OAI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1339),
.A2(n_1363),
.B1(n_1346),
.B2(n_1341),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1247),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1325),
.A2(n_1306),
.B1(n_1363),
.B2(n_1341),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1228),
.Y(n_1449)
);

BUFx4f_ASAP7_75t_L g1450 ( 
.A(n_1356),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1247),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1339),
.B(n_1346),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1349),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1235),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1352),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1232),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1355),
.A2(n_1357),
.B1(n_1254),
.B2(n_1219),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1219),
.A2(n_1248),
.B1(n_1210),
.B2(n_1362),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1358),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1358),
.Y(n_1460)
);

OR2x6_ASAP7_75t_L g1461 ( 
.A(n_1227),
.B(n_1354),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1217),
.A2(n_1337),
.B1(n_1314),
.B2(n_1243),
.Y(n_1462)
);

CKINVDCx11_ASAP7_75t_R g1463 ( 
.A(n_1279),
.Y(n_1463)
);

CKINVDCx11_ASAP7_75t_R g1464 ( 
.A(n_1286),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1250),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1232),
.Y(n_1466)
);

OAI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1311),
.A2(n_1255),
.B1(n_1291),
.B2(n_1294),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1263),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1288),
.B(n_1252),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1295),
.A2(n_1293),
.B1(n_1304),
.B2(n_1276),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1247),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1304),
.B(n_1247),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1304),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1290),
.B(n_1292),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1329),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1250),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1329),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1329),
.Y(n_1478)
);

AO21x1_ASAP7_75t_SL g1479 ( 
.A1(n_1253),
.A2(n_1080),
.B(n_1239),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1220),
.B(n_1230),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1333),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1283),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1242),
.B(n_1063),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1319),
.A2(n_1000),
.B1(n_926),
.B2(n_1063),
.Y(n_1484)
);

BUFx12f_ASAP7_75t_L g1485 ( 
.A(n_1216),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1208),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1303),
.A2(n_1086),
.B(n_1087),
.Y(n_1487)
);

BUFx4f_ASAP7_75t_SL g1488 ( 
.A(n_1212),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1218),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1333),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1242),
.B(n_1063),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1319),
.A2(n_1000),
.B1(n_927),
.B2(n_1063),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1218),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1208),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1319),
.A2(n_1000),
.B1(n_927),
.B2(n_1063),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1206),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1206),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1333),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1333),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1218),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1322),
.B(n_1239),
.Y(n_1501)
);

BUFx2_ASAP7_75t_R g1502 ( 
.A(n_1221),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1220),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1298),
.B(n_1309),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1303),
.A2(n_1086),
.B(n_1087),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1218),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1218),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1218),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1218),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1208),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1333),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1319),
.A2(n_1000),
.B1(n_926),
.B2(n_1174),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1206),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1218),
.Y(n_1514)
);

INVx6_ASAP7_75t_L g1515 ( 
.A(n_1210),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1412),
.A2(n_1390),
.B(n_1409),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1417),
.B(n_1418),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1410),
.B(n_1420),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1389),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1481),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1490),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1498),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1469),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_L g1524 ( 
.A(n_1377),
.B(n_1407),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1499),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1469),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1420),
.Y(n_1527)
);

AOI21xp33_ASAP7_75t_L g1528 ( 
.A1(n_1484),
.A2(n_1512),
.B(n_1382),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1472),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1378),
.B(n_1413),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_1414),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1435),
.A2(n_1505),
.B(n_1487),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1431),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1483),
.B(n_1491),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1455),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1431),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1431),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1369),
.Y(n_1538)
);

BUFx12f_ASAP7_75t_L g1539 ( 
.A(n_1453),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1366),
.B(n_1365),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1424),
.B(n_1364),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1367),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1364),
.B(n_1504),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1364),
.B(n_1504),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1373),
.A2(n_1438),
.B(n_1467),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1492),
.A2(n_1495),
.B(n_1388),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1370),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1406),
.Y(n_1548)
);

INVxp67_ASAP7_75t_SL g1549 ( 
.A(n_1482),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1374),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1504),
.B(n_1437),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1473),
.B(n_1443),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1383),
.B(n_1501),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1385),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1406),
.Y(n_1555)
);

OR2x6_ASAP7_75t_L g1556 ( 
.A(n_1366),
.B(n_1461),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1437),
.B(n_1393),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1438),
.A2(n_1402),
.B(n_1421),
.Y(n_1558)
);

NAND2x1p5_ASAP7_75t_L g1559 ( 
.A(n_1374),
.B(n_1416),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1511),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1455),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1423),
.B(n_1366),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1366),
.B(n_1443),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1489),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1493),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1479),
.B(n_1368),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1500),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_SL g1568 ( 
.A(n_1386),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1506),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1454),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1507),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1433),
.B(n_1439),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1508),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1391),
.B(n_1461),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1441),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1509),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1514),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1394),
.Y(n_1578)
);

NOR2xp67_ASAP7_75t_SL g1579 ( 
.A(n_1392),
.B(n_1485),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1396),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1397),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1496),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1515),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1497),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1442),
.A2(n_1474),
.B(n_1513),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1497),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1395),
.B(n_1401),
.Y(n_1587)
);

INVx8_ASAP7_75t_L g1588 ( 
.A(n_1379),
.Y(n_1588)
);

AO21x2_ASAP7_75t_L g1589 ( 
.A1(n_1428),
.A2(n_1432),
.B(n_1405),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1479),
.B(n_1372),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1381),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1440),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1436),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1475),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1369),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1376),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1447),
.A2(n_1471),
.B(n_1458),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1427),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1478),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1404),
.B(n_1376),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_L g1601 ( 
.A(n_1448),
.B(n_1425),
.C(n_1457),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1478),
.Y(n_1602)
);

INVxp33_ASAP7_75t_L g1603 ( 
.A(n_1452),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1446),
.B(n_1452),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1470),
.A2(n_1449),
.B(n_1459),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1372),
.B(n_1387),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1372),
.B(n_1387),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1375),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1375),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1375),
.Y(n_1610)
);

CKINVDCx6p67_ASAP7_75t_R g1611 ( 
.A(n_1392),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1380),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1400),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1450),
.A2(n_1445),
.B(n_1419),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1462),
.A2(n_1450),
.B(n_1468),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1380),
.B(n_1503),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1400),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1384),
.B(n_1503),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1384),
.B(n_1503),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1398),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1400),
.Y(n_1621)
);

INVx4_ASAP7_75t_L g1622 ( 
.A(n_1540),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1550),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1556),
.B(n_1590),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1550),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1523),
.B(n_1456),
.Y(n_1626)
);

INVx5_ASAP7_75t_L g1627 ( 
.A(n_1556),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1523),
.B(n_1460),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1526),
.B(n_1444),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1518),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1589),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1517),
.B(n_1480),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1530),
.B(n_1534),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1542),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1589),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1517),
.B(n_1480),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1574),
.B(n_1466),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1548),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1587),
.B(n_1480),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1548),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1541),
.B(n_1434),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1552),
.B(n_1434),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1519),
.B(n_1398),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1528),
.A2(n_1386),
.B1(n_1371),
.B2(n_1450),
.C(n_1453),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1555),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1590),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1574),
.B(n_1371),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1533),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1589),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1555),
.Y(n_1650)
);

NOR2x1_ASAP7_75t_SL g1651 ( 
.A(n_1556),
.B(n_1451),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1540),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1520),
.B(n_1381),
.Y(n_1653)
);

OAI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1546),
.A2(n_1515),
.B1(n_1381),
.B2(n_1476),
.C(n_1465),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1547),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1521),
.B(n_1381),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1547),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1551),
.B(n_1486),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1522),
.B(n_1515),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1570),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1525),
.B(n_1515),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1556),
.B(n_1486),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1551),
.B(n_1476),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1563),
.B(n_1451),
.Y(n_1664)
);

INVxp67_ASAP7_75t_L g1665 ( 
.A(n_1535),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1524),
.A2(n_1463),
.B1(n_1464),
.B2(n_1485),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1536),
.B(n_1537),
.Y(n_1667)
);

BUFx12f_ASAP7_75t_L g1668 ( 
.A(n_1539),
.Y(n_1668)
);

AND2x4_ASAP7_75t_SL g1669 ( 
.A(n_1540),
.B(n_1430),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1575),
.B(n_1543),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1554),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1604),
.B(n_1510),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1553),
.B(n_1549),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1559),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1553),
.B(n_1464),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1518),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1603),
.A2(n_1494),
.B1(n_1403),
.B2(n_1408),
.C(n_1411),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1544),
.B(n_1403),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1564),
.B(n_1494),
.Y(n_1679)
);

INVxp67_ASAP7_75t_SL g1680 ( 
.A(n_1559),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1565),
.B(n_1494),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1524),
.A2(n_1463),
.B1(n_1429),
.B2(n_1415),
.Y(n_1682)
);

BUFx3_ASAP7_75t_L g1683 ( 
.A(n_1559),
.Y(n_1683)
);

INVx3_ASAP7_75t_L g1684 ( 
.A(n_1518),
.Y(n_1684)
);

OAI221xp5_ASAP7_75t_SL g1685 ( 
.A1(n_1666),
.A2(n_1557),
.B1(n_1682),
.B2(n_1572),
.C(n_1644),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1668),
.A2(n_1601),
.B1(n_1600),
.B2(n_1557),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1654),
.A2(n_1566),
.B1(n_1540),
.B2(n_1642),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1633),
.B(n_1604),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1673),
.B(n_1561),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1660),
.B(n_1593),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1675),
.A2(n_1566),
.B(n_1572),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1665),
.B(n_1593),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1638),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1677),
.B(n_1558),
.C(n_1615),
.Y(n_1694)
);

OAI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1653),
.A2(n_1585),
.B(n_1558),
.Y(n_1695)
);

NAND4xp25_ASAP7_75t_SL g1696 ( 
.A(n_1641),
.B(n_1620),
.C(n_1639),
.D(n_1642),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1664),
.B(n_1612),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1640),
.B(n_1592),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1645),
.B(n_1592),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1672),
.B(n_1558),
.C(n_1618),
.Y(n_1700)
);

AOI211xp5_ASAP7_75t_L g1701 ( 
.A1(n_1647),
.A2(n_1596),
.B(n_1616),
.C(n_1562),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1672),
.A2(n_1558),
.B1(n_1611),
.B2(n_1612),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1627),
.B(n_1606),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1624),
.B(n_1562),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1664),
.B(n_1538),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1627),
.B(n_1606),
.Y(n_1706)
);

OAI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1643),
.A2(n_1579),
.B1(n_1656),
.B2(n_1659),
.C(n_1661),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1670),
.B(n_1545),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1641),
.A2(n_1611),
.B1(n_1568),
.B2(n_1595),
.Y(n_1709)
);

OAI21xp33_ASAP7_75t_L g1710 ( 
.A1(n_1637),
.A2(n_1598),
.B(n_1560),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1663),
.A2(n_1568),
.B1(n_1531),
.B2(n_1616),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1651),
.A2(n_1545),
.B1(n_1652),
.B2(n_1622),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1650),
.B(n_1567),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1663),
.A2(n_1568),
.B1(n_1426),
.B2(n_1614),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1662),
.A2(n_1579),
.B(n_1617),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1650),
.B(n_1567),
.Y(n_1716)
);

OAI221xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1658),
.A2(n_1637),
.B1(n_1680),
.B2(n_1626),
.C(n_1628),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1627),
.B(n_1607),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1627),
.B(n_1607),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1658),
.A2(n_1585),
.B(n_1597),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1662),
.A2(n_1621),
.B(n_1613),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1632),
.B(n_1569),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1632),
.B(n_1569),
.Y(n_1723)
);

OAI221xp5_ASAP7_75t_SL g1724 ( 
.A1(n_1626),
.A2(n_1573),
.B1(n_1576),
.B2(n_1577),
.C(n_1578),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1655),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1669),
.A2(n_1583),
.B1(n_1591),
.B2(n_1613),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1636),
.B(n_1571),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1636),
.B(n_1571),
.Y(n_1728)
);

OAI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1674),
.A2(n_1583),
.B1(n_1591),
.B2(n_1581),
.C(n_1577),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1655),
.A2(n_1578),
.B1(n_1580),
.B2(n_1581),
.C(n_1671),
.Y(n_1730)
);

NOR3xp33_ASAP7_75t_L g1731 ( 
.A(n_1622),
.B(n_1597),
.C(n_1529),
.Y(n_1731)
);

AND2x2_ASAP7_75t_SL g1732 ( 
.A(n_1622),
.B(n_1516),
.Y(n_1732)
);

NAND3xp33_ASAP7_75t_L g1733 ( 
.A(n_1631),
.B(n_1605),
.C(n_1599),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_SL g1734 ( 
.A(n_1668),
.B(n_1422),
.Y(n_1734)
);

NAND3xp33_ASAP7_75t_L g1735 ( 
.A(n_1631),
.B(n_1605),
.C(n_1599),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1657),
.A2(n_1602),
.B1(n_1594),
.B2(n_1584),
.C(n_1586),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1630),
.B(n_1605),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1629),
.B(n_1602),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1679),
.B(n_1527),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1635),
.B(n_1608),
.C(n_1609),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1676),
.B(n_1516),
.Y(n_1741)
);

AND2x2_ASAP7_75t_SL g1742 ( 
.A(n_1622),
.B(n_1532),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_L g1743 ( 
.A(n_1635),
.B(n_1609),
.C(n_1608),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1678),
.B(n_1619),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1657),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1627),
.B(n_1610),
.Y(n_1746)
);

NAND4xp25_ASAP7_75t_L g1747 ( 
.A(n_1679),
.B(n_1594),
.C(n_1582),
.D(n_1584),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1627),
.B(n_1610),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1662),
.A2(n_1669),
.B(n_1624),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1720),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1693),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1725),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1700),
.B(n_1733),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1704),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1708),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1741),
.B(n_1704),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1688),
.B(n_1649),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1745),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1688),
.B(n_1649),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1742),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1704),
.Y(n_1761)
);

AND2x4_ASAP7_75t_SL g1762 ( 
.A(n_1731),
.B(n_1652),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1737),
.Y(n_1763)
);

HB1xp67_ASAP7_75t_L g1764 ( 
.A(n_1737),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1738),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1713),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1716),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1732),
.B(n_1684),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1732),
.B(n_1646),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1739),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1698),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1699),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1746),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1744),
.B(n_1695),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1735),
.B(n_1667),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1740),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1703),
.B(n_1624),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1729),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1703),
.B(n_1648),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1706),
.B(n_1648),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1743),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1747),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1697),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1692),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1690),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1746),
.Y(n_1787)
);

INVx4_ASAP7_75t_L g1788 ( 
.A(n_1705),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1701),
.B(n_1683),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1730),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1689),
.B(n_1634),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1748),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1722),
.Y(n_1793)
);

NAND2x1_ASAP7_75t_L g1794 ( 
.A(n_1694),
.B(n_1652),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1723),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1724),
.Y(n_1796)
);

INVxp67_ASAP7_75t_SL g1797 ( 
.A(n_1717),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1758),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1797),
.A2(n_1691),
.B(n_1685),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1782),
.B(n_1727),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1758),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1780),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1782),
.B(n_1728),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1782),
.B(n_1702),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1776),
.B(n_1623),
.Y(n_1805)
);

INVxp67_ASAP7_75t_SL g1806 ( 
.A(n_1777),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1780),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1752),
.Y(n_1808)
);

AND2x4_ASAP7_75t_SL g1809 ( 
.A(n_1788),
.B(n_1652),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1752),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1754),
.B(n_1718),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1770),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1752),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1761),
.B(n_1712),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1761),
.B(n_1749),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1767),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1785),
.B(n_1710),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1785),
.B(n_1711),
.Y(n_1818)
);

INVx3_ASAP7_75t_L g1819 ( 
.A(n_1756),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1776),
.B(n_1623),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1796),
.B(n_1681),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1796),
.B(n_1681),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1780),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1797),
.B(n_1707),
.Y(n_1824)
);

INVxp67_ASAP7_75t_SL g1825 ( 
.A(n_1777),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1781),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1751),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1767),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1786),
.B(n_1772),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1786),
.B(n_1715),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1767),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1751),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1776),
.B(n_1623),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1781),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1789),
.A2(n_1686),
.B(n_1714),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1768),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1772),
.B(n_1625),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1757),
.B(n_1625),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1773),
.B(n_1625),
.Y(n_1839)
);

NAND5xp2_ASAP7_75t_L g1840 ( 
.A(n_1779),
.B(n_1734),
.C(n_1687),
.D(n_1750),
.E(n_1790),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_SL g1841 ( 
.A(n_1788),
.B(n_1502),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1793),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1784),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1773),
.B(n_1736),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1768),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1783),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1768),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1789),
.A2(n_1696),
.B1(n_1662),
.B2(n_1709),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1771),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1781),
.Y(n_1850)
);

AOI211xp5_ASAP7_75t_L g1851 ( 
.A1(n_1753),
.A2(n_1721),
.B(n_1718),
.C(n_1719),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1827),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1812),
.B(n_1760),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1835),
.A2(n_1753),
.B(n_1779),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1812),
.B(n_1760),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1821),
.B(n_1790),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1815),
.B(n_1762),
.Y(n_1857)
);

HB1xp67_ASAP7_75t_L g1858 ( 
.A(n_1832),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1806),
.B(n_1753),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1808),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1808),
.Y(n_1861)
);

NOR2x1p5_ASAP7_75t_SL g1862 ( 
.A(n_1804),
.B(n_1760),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1815),
.B(n_1760),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1810),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1822),
.B(n_1790),
.Y(n_1865)
);

AOI21xp33_ASAP7_75t_L g1866 ( 
.A1(n_1799),
.A2(n_1794),
.B(n_1750),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1810),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1824),
.B(n_1783),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1827),
.Y(n_1869)
);

AOI221xp5_ASAP7_75t_L g1870 ( 
.A1(n_1825),
.A2(n_1750),
.B1(n_1783),
.B2(n_1794),
.C(n_1757),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1844),
.B(n_1759),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1813),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1830),
.B(n_1800),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1804),
.B(n_1759),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1800),
.B(n_1793),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1813),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_SL g1877 ( 
.A(n_1841),
.B(n_1788),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1798),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1814),
.B(n_1766),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1842),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1803),
.B(n_1775),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1814),
.B(n_1766),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1803),
.B(n_1775),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1798),
.Y(n_1884)
);

INVx3_ASAP7_75t_L g1885 ( 
.A(n_1819),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1811),
.B(n_1766),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1801),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1818),
.B(n_1775),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1811),
.B(n_1766),
.Y(n_1889)
);

NOR4xp25_ASAP7_75t_L g1890 ( 
.A(n_1846),
.B(n_1774),
.C(n_1787),
.D(n_1792),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1802),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1811),
.B(n_1778),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1817),
.B(n_1851),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1801),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1819),
.B(n_1843),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1816),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1809),
.B(n_1819),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1829),
.B(n_1795),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1837),
.B(n_1795),
.Y(n_1899)
);

NAND2x1p5_ASAP7_75t_L g1900 ( 
.A(n_1805),
.B(n_1794),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1805),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1802),
.B(n_1763),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1807),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1816),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1848),
.A2(n_1761),
.B1(n_1788),
.B2(n_1770),
.Y(n_1905)
);

NAND2x1p5_ASAP7_75t_L g1906 ( 
.A(n_1820),
.B(n_1719),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1860),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1859),
.B(n_1874),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1906),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1857),
.B(n_1762),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1860),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1863),
.B(n_1807),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1859),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1852),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1906),
.Y(n_1915)
);

INVxp67_ASAP7_75t_SL g1916 ( 
.A(n_1880),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1857),
.B(n_1762),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1861),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1863),
.B(n_1823),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1861),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1874),
.B(n_1823),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1875),
.B(n_1826),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1897),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1892),
.B(n_1826),
.Y(n_1924)
);

OR2x6_ASAP7_75t_L g1925 ( 
.A(n_1854),
.B(n_1852),
.Y(n_1925)
);

INVx1_ASAP7_75t_SL g1926 ( 
.A(n_1869),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1857),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1881),
.B(n_1834),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1892),
.B(n_1834),
.Y(n_1929)
);

INVx1_ASAP7_75t_SL g1930 ( 
.A(n_1869),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1856),
.B(n_1763),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1906),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1858),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1883),
.B(n_1850),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1873),
.B(n_1850),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1886),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1865),
.B(n_1764),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1900),
.Y(n_1938)
);

CKINVDCx14_ASAP7_75t_R g1939 ( 
.A(n_1905),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1868),
.B(n_1764),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1871),
.B(n_1893),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1901),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1884),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1879),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1879),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1882),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1888),
.B(n_1795),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1864),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1882),
.B(n_1809),
.Y(n_1949)
);

INVx3_ASAP7_75t_L g1950 ( 
.A(n_1910),
.Y(n_1950)
);

OAI21xp33_ASAP7_75t_L g1951 ( 
.A1(n_1925),
.A2(n_1840),
.B(n_1866),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1927),
.Y(n_1952)
);

AOI32xp33_ASAP7_75t_L g1953 ( 
.A1(n_1941),
.A2(n_1870),
.A3(n_1853),
.B1(n_1855),
.B2(n_1889),
.Y(n_1953)
);

OAI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1925),
.A2(n_1939),
.B(n_1890),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1933),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1943),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1943),
.Y(n_1957)
);

NOR3xp33_ASAP7_75t_SL g1958 ( 
.A(n_1916),
.B(n_1887),
.C(n_1884),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1945),
.B(n_1899),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1925),
.A2(n_1877),
.B1(n_1855),
.B2(n_1853),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1927),
.Y(n_1961)
);

INVxp67_ASAP7_75t_SL g1962 ( 
.A(n_1908),
.Y(n_1962)
);

NAND3xp33_ASAP7_75t_SL g1963 ( 
.A(n_1942),
.B(n_1900),
.C(n_1895),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1943),
.Y(n_1964)
);

AOI32xp33_ASAP7_75t_L g1965 ( 
.A1(n_1942),
.A2(n_1913),
.A3(n_1946),
.B1(n_1944),
.B2(n_1926),
.Y(n_1965)
);

AOI221xp5_ASAP7_75t_L g1966 ( 
.A1(n_1914),
.A2(n_1878),
.B1(n_1887),
.B2(n_1894),
.C(n_1900),
.Y(n_1966)
);

NOR2x1_ASAP7_75t_L g1967 ( 
.A(n_1925),
.B(n_1894),
.Y(n_1967)
);

AOI211xp5_ASAP7_75t_L g1968 ( 
.A1(n_1930),
.A2(n_1889),
.B(n_1886),
.C(n_1895),
.Y(n_1968)
);

INVxp33_ASAP7_75t_L g1969 ( 
.A(n_1949),
.Y(n_1969)
);

AOI222xp33_ASAP7_75t_L g1970 ( 
.A1(n_1944),
.A2(n_1862),
.B1(n_1946),
.B2(n_1940),
.C1(n_1931),
.C2(n_1937),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1907),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1908),
.B(n_1936),
.Y(n_1972)
);

AOI32xp33_ASAP7_75t_L g1973 ( 
.A1(n_1949),
.A2(n_1897),
.A3(n_1762),
.B1(n_1770),
.B2(n_1778),
.Y(n_1973)
);

INVx2_ASAP7_75t_SL g1974 ( 
.A(n_1923),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1907),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1910),
.B(n_1897),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1936),
.B(n_1898),
.Y(n_1977)
);

INVxp67_ASAP7_75t_SL g1978 ( 
.A(n_1938),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1911),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1962),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1969),
.B(n_1925),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1976),
.B(n_1923),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1951),
.B(n_1539),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1952),
.B(n_1862),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1961),
.B(n_1924),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1967),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1955),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1950),
.B(n_1415),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1950),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_1978),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1974),
.B(n_1924),
.Y(n_1991)
);

INVxp67_ASAP7_75t_L g1992 ( 
.A(n_1956),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1972),
.B(n_1935),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1958),
.B(n_1910),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1957),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1972),
.B(n_1935),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1960),
.B(n_1910),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1971),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1975),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1968),
.B(n_1917),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1963),
.B(n_1917),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1959),
.B(n_1922),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1954),
.B(n_1917),
.Y(n_2003)
);

OAI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_2001),
.A2(n_1954),
.B1(n_1965),
.B2(n_1953),
.Y(n_2004)
);

AOI221xp5_ASAP7_75t_L g2005 ( 
.A1(n_1990),
.A2(n_1966),
.B1(n_1964),
.B2(n_1979),
.C(n_1973),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1985),
.B(n_1977),
.Y(n_2006)
);

AOI21xp33_ASAP7_75t_SL g2007 ( 
.A1(n_1981),
.A2(n_1970),
.B(n_1917),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1984),
.B(n_1970),
.Y(n_2008)
);

OAI211xp5_ASAP7_75t_L g2009 ( 
.A1(n_1986),
.A2(n_1938),
.B(n_1909),
.C(n_1932),
.Y(n_2009)
);

AOI221xp5_ASAP7_75t_L g2010 ( 
.A1(n_1987),
.A2(n_1909),
.B1(n_1915),
.B2(n_1932),
.C(n_1948),
.Y(n_2010)
);

AOI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1986),
.A2(n_1915),
.B(n_1947),
.Y(n_2011)
);

NAND3xp33_ASAP7_75t_L g2012 ( 
.A(n_1980),
.B(n_1918),
.C(n_1911),
.Y(n_2012)
);

NAND4xp25_ASAP7_75t_L g2013 ( 
.A(n_1983),
.B(n_1928),
.C(n_1934),
.D(n_1922),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1988),
.B(n_1429),
.Y(n_2014)
);

AOI222xp33_ASAP7_75t_L g2015 ( 
.A1(n_1994),
.A2(n_1948),
.B1(n_1920),
.B2(n_1918),
.C1(n_1929),
.C2(n_1919),
.Y(n_2015)
);

O2A1O1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1980),
.A2(n_1920),
.B(n_1921),
.C(n_1928),
.Y(n_2016)
);

AOI32xp33_ASAP7_75t_L g2017 ( 
.A1(n_1994),
.A2(n_1929),
.A3(n_1919),
.B1(n_1912),
.B2(n_1934),
.Y(n_2017)
);

NAND4xp25_ASAP7_75t_L g2018 ( 
.A(n_1997),
.B(n_1921),
.C(n_1912),
.D(n_1885),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1982),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_2004),
.A2(n_1989),
.B1(n_1991),
.B2(n_2002),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_2008),
.A2(n_1982),
.B1(n_2000),
.B2(n_1997),
.Y(n_2021)
);

NOR3xp33_ASAP7_75t_L g2022 ( 
.A(n_2007),
.B(n_1992),
.C(n_2003),
.Y(n_2022)
);

NOR3x1_ASAP7_75t_L g2023 ( 
.A(n_2009),
.B(n_1999),
.C(n_1998),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2019),
.Y(n_2024)
);

NOR3xp33_ASAP7_75t_L g2025 ( 
.A(n_2005),
.B(n_2003),
.C(n_1995),
.Y(n_2025)
);

NAND4xp75_ASAP7_75t_L g2026 ( 
.A(n_2010),
.B(n_2000),
.C(n_1999),
.D(n_1998),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_2014),
.B(n_1993),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_2017),
.B(n_1993),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_2006),
.B(n_1996),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_2015),
.B(n_2002),
.Y(n_2030)
);

AND3x1_ASAP7_75t_L g2031 ( 
.A(n_2016),
.B(n_1885),
.C(n_1891),
.Y(n_2031)
);

NAND3xp33_ASAP7_75t_SL g2032 ( 
.A(n_2025),
.B(n_2011),
.C(n_1996),
.Y(n_2032)
);

NOR4xp25_ASAP7_75t_L g2033 ( 
.A(n_2030),
.B(n_2012),
.C(n_2018),
.D(n_2013),
.Y(n_2033)
);

NAND3xp33_ASAP7_75t_SL g2034 ( 
.A(n_2022),
.B(n_1902),
.C(n_1833),
.Y(n_2034)
);

OAI311xp33_ASAP7_75t_L g2035 ( 
.A1(n_2021),
.A2(n_1902),
.A3(n_1885),
.B1(n_1820),
.C1(n_1833),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2020),
.B(n_1891),
.Y(n_2036)
);

AOI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_2028),
.A2(n_1399),
.B(n_1896),
.Y(n_2037)
);

OAI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_2031),
.A2(n_1903),
.B1(n_1904),
.B2(n_1896),
.C(n_1864),
.Y(n_2038)
);

AOI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_2026),
.A2(n_1904),
.B1(n_1903),
.B2(n_1876),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2024),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2036),
.Y(n_2041)
);

NOR2x1p5_ASAP7_75t_L g2042 ( 
.A(n_2034),
.B(n_2023),
.Y(n_2042)
);

NOR2x1_ASAP7_75t_L g2043 ( 
.A(n_2032),
.B(n_2029),
.Y(n_2043)
);

AND3x4_ASAP7_75t_L g2044 ( 
.A(n_2033),
.B(n_2027),
.C(n_1488),
.Y(n_2044)
);

INVxp67_ASAP7_75t_L g2045 ( 
.A(n_2040),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2039),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2038),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2037),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_2035),
.B(n_1867),
.Y(n_2049)
);

NAND3xp33_ASAP7_75t_SL g2050 ( 
.A(n_2044),
.B(n_1872),
.C(n_1867),
.Y(n_2050)
);

XOR2xp5_ASAP7_75t_L g2051 ( 
.A(n_2043),
.B(n_1726),
.Y(n_2051)
);

BUFx6f_ASAP7_75t_L g2052 ( 
.A(n_2048),
.Y(n_2052)
);

NAND4xp75_ASAP7_75t_L g2053 ( 
.A(n_2046),
.B(n_1876),
.C(n_1872),
.D(n_1778),
.Y(n_2053)
);

NOR4xp75_ASAP7_75t_L g2054 ( 
.A(n_2042),
.B(n_1839),
.C(n_1769),
.D(n_1791),
.Y(n_2054)
);

NAND4xp75_ASAP7_75t_L g2055 ( 
.A(n_2041),
.B(n_1792),
.C(n_1787),
.D(n_1774),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_2049),
.A2(n_2047),
.B(n_2045),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_2053),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2051),
.Y(n_2058)
);

NOR3xp33_ASAP7_75t_L g2059 ( 
.A(n_2056),
.B(n_2049),
.C(n_1788),
.Y(n_2059)
);

XNOR2xp5_ASAP7_75t_L g2060 ( 
.A(n_2054),
.B(n_1769),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_2058),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2059),
.A2(n_2052),
.B1(n_2050),
.B2(n_2055),
.Y(n_2062)
);

XNOR2xp5_ASAP7_75t_L g2063 ( 
.A(n_2062),
.B(n_2061),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_2063),
.A2(n_2057),
.B1(n_2060),
.B2(n_1828),
.Y(n_2064)
);

AOI221x1_ASAP7_75t_L g2065 ( 
.A1(n_2063),
.A2(n_1831),
.B1(n_1847),
.B2(n_1845),
.C(n_1836),
.Y(n_2065)
);

OAI22xp33_ASAP7_75t_SL g2066 ( 
.A1(n_2064),
.A2(n_1828),
.B1(n_1847),
.B2(n_1845),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_2065),
.A2(n_1836),
.B(n_1831),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_2067),
.A2(n_1849),
.B1(n_1838),
.B2(n_1774),
.Y(n_2068)
);

AOI21xp33_ASAP7_75t_SL g2069 ( 
.A1(n_2066),
.A2(n_1838),
.B(n_1588),
.Y(n_2069)
);

OAI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_2069),
.A2(n_2068),
.B(n_1849),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_2070),
.A2(n_1792),
.B1(n_1787),
.B2(n_1774),
.Y(n_2071)
);

AOI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_2071),
.A2(n_1792),
.B1(n_1787),
.B2(n_1765),
.C(n_1755),
.Y(n_2072)
);

AOI211xp5_ASAP7_75t_L g2073 ( 
.A1(n_2072),
.A2(n_1408),
.B(n_1411),
.C(n_1477),
.Y(n_2073)
);


endmodule