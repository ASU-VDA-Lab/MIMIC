module fake_jpeg_3488_n_476 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_54),
.Y(n_146)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_30),
.Y(n_55)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_57),
.Y(n_175)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_58),
.Y(n_190)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_61),
.B(n_108),
.Y(n_122)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_62),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_63),
.B(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_26),
.B(n_8),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_8),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_83),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_72),
.Y(n_178)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_51),
.Y(n_74)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_76),
.Y(n_183)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_79),
.A2(n_21),
.B1(n_25),
.B2(n_6),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g188 ( 
.A(n_81),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_82),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_26),
.B(n_7),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_87),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_88),
.Y(n_120)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_90),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_18),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_91),
.B(n_113),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_92),
.Y(n_197)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_106),
.Y(n_159)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_99),
.Y(n_199)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_37),
.B(n_11),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_107),
.Y(n_132)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_23),
.B(n_11),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g109 ( 
.A(n_51),
.Y(n_109)
);

BUFx2_ASAP7_75t_R g193 ( 
.A(n_109),
.Y(n_193)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_21),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_111),
.B(n_112),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_29),
.B(n_1),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_37),
.B(n_13),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_61),
.Y(n_127)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_89),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_19),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_32),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g203 ( 
.A(n_118),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_127),
.B(n_172),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_34),
.B1(n_52),
.B2(n_48),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_129),
.A2(n_134),
.B1(n_139),
.B2(n_145),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_54),
.A2(n_29),
.B1(n_52),
.B2(n_48),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_135),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_137),
.B(n_142),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_46),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_138),
.B(n_160),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_46),
.B1(n_43),
.B2(n_33),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_43),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_100),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_144),
.B(n_165),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_47),
.B1(n_31),
.B2(n_41),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_78),
.B1(n_76),
.B2(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_148),
.A2(n_162),
.B1(n_167),
.B2(n_177),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_79),
.A2(n_33),
.B1(n_44),
.B2(n_38),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_150),
.A2(n_154),
.B1(n_157),
.B2(n_6),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_60),
.A2(n_53),
.B1(n_44),
.B2(n_38),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_71),
.A2(n_53),
.B1(n_41),
.B2(n_32),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_19),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_161),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_73),
.A2(n_31),
.B1(n_47),
.B2(n_25),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_82),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_87),
.B(n_16),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_166),
.B(n_169),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_92),
.A2(n_25),
.B1(n_39),
.B2(n_16),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_65),
.B(n_16),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_93),
.B(n_17),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_88),
.B(n_39),
.C(n_25),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_174),
.B(n_180),
.C(n_159),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_106),
.A2(n_25),
.B1(n_21),
.B2(n_6),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_68),
.B(n_14),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_181),
.B(n_187),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_74),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_120),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_177),
.B(n_198),
.Y(n_218)
);

OR2x2_ASAP7_75t_SL g186 ( 
.A(n_107),
.B(n_25),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_186),
.B(n_201),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_68),
.B(n_14),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_55),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_194),
.B1(n_192),
.B2(n_153),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_114),
.B(n_14),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_204),
.A2(n_209),
.B1(n_224),
.B2(n_227),
.Y(n_310)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_205),
.Y(n_314)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_207),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_146),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_208),
.B(n_221),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_157),
.A2(n_200),
.B1(n_154),
.B2(n_161),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_213),
.Y(n_307)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_214),
.Y(n_321)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_215),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_218),
.A2(n_228),
.B1(n_270),
.B2(n_272),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_126),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g293 ( 
.A(n_219),
.B(n_238),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_148),
.A2(n_145),
.B1(n_133),
.B2(n_143),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_220),
.A2(n_262),
.B1(n_273),
.B2(n_226),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_146),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_223),
.Y(n_297)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_225),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_190),
.A2(n_185),
.B1(n_130),
.B2(n_136),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_185),
.A2(n_130),
.B1(n_128),
.B2(n_159),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_171),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_229),
.B(n_232),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_230),
.Y(n_324)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_231),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_131),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_147),
.Y(n_234)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_125),
.Y(n_235)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_235),
.Y(n_318)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_237),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_124),
.B(n_191),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_240),
.B(n_242),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_132),
.B(n_122),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_241),
.B(n_244),
.Y(n_320)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_123),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_175),
.B(n_163),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_139),
.B(n_189),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_248),
.Y(n_282)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_252),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_152),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_134),
.B(n_180),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_250),
.Y(n_309)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_178),
.B(n_179),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_251),
.B(n_253),
.Y(n_322)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_125),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_152),
.B(n_170),
.Y(n_253)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_170),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_178),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_255),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_183),
.A2(n_140),
.B1(n_162),
.B2(n_119),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_256),
.A2(n_265),
.B1(n_267),
.B2(n_266),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_131),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_257),
.Y(n_299)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_179),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_261),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_125),
.A2(n_155),
.B(n_173),
.C(n_149),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_266),
.B(n_265),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_119),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_176),
.A2(n_197),
.B1(n_195),
.B2(n_183),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_264),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_195),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_197),
.A2(n_149),
.B1(n_151),
.B2(n_199),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_203),
.A2(n_149),
.B(n_151),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_155),
.A2(n_121),
.B1(n_199),
.B2(n_151),
.Y(n_267)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_199),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_274),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_203),
.B(n_173),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_219),
.C(n_238),
.Y(n_304)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_173),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_168),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_305),
.B1(n_316),
.B2(n_287),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_287),
.A2(n_310),
.B1(n_281),
.B2(n_311),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_220),
.A2(n_204),
.B1(n_209),
.B2(n_256),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_296),
.A2(n_298),
.B1(n_306),
.B2(n_317),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_239),
.A2(n_243),
.B1(n_262),
.B2(n_240),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_217),
.B(n_222),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_302),
.C(n_311),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_243),
.B(n_268),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_260),
.A2(n_216),
.B(n_238),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g346 ( 
.A1(n_303),
.A2(n_293),
.B(n_279),
.Y(n_346)
);

OAI21xp33_ASAP7_75t_L g361 ( 
.A1(n_304),
.A2(n_301),
.B(n_321),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_236),
.A2(n_263),
.B1(n_219),
.B2(n_211),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_214),
.A2(n_274),
.B1(n_231),
.B2(n_246),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_SL g311 ( 
.A(n_233),
.B(n_271),
.C(n_259),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_254),
.A2(n_247),
.B1(n_242),
.B2(n_237),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_225),
.A2(n_252),
.B1(n_272),
.B2(n_210),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_206),
.A2(n_213),
.B1(n_270),
.B2(n_205),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_319),
.A2(n_323),
.B1(n_286),
.B2(n_276),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_271),
.A2(n_220),
.B1(n_226),
.B2(n_273),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_325),
.Y(n_363)
);

OR2x2_ASAP7_75t_SL g326 ( 
.A(n_304),
.B(n_235),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_326),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_300),
.B(n_269),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_327),
.B(n_329),
.Y(n_369)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_328),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_295),
.A2(n_309),
.B(n_282),
.C(n_303),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_330),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_302),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_357),
.C(n_306),
.Y(n_364)
);

INVx13_ASAP7_75t_L g333 ( 
.A(n_314),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_291),
.B(n_320),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_334),
.B(n_346),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_335),
.A2(n_350),
.B1(n_349),
.B2(n_332),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_324),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_336),
.B(n_338),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_295),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_348),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_279),
.B(n_289),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_341),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_323),
.A2(n_296),
.B1(n_281),
.B2(n_298),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_340),
.A2(n_285),
.B1(n_301),
.B2(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_284),
.Y(n_342)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_275),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_356),
.Y(n_366)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_345),
.B(n_347),
.Y(n_382)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

O2A1O1Ixp33_ASAP7_75t_L g348 ( 
.A1(n_293),
.A2(n_318),
.B(n_292),
.C(n_289),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_305),
.A2(n_280),
.B1(n_316),
.B2(n_285),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_288),
.B(n_292),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_351),
.B(n_352),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_278),
.B(n_294),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_297),
.B(n_313),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_354),
.Y(n_372)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_313),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_278),
.B(n_294),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_293),
.B(n_297),
.C(n_312),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_308),
.A2(n_318),
.B(n_312),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_361),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_308),
.B(n_277),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_360),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_308),
.B(n_277),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_362),
.A2(n_385),
.B1(n_350),
.B2(n_332),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_343),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_353),
.Y(n_370)
);

BUFx24_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_359),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_376),
.Y(n_395)
);

AND2x6_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_307),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_381),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_331),
.B(n_283),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_326),
.C(n_329),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_339),
.A2(n_307),
.B1(n_341),
.B2(n_325),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_379),
.A2(n_349),
.B1(n_330),
.B2(n_342),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_334),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_327),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_345),
.B(n_347),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_357),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_368),
.A2(n_332),
.B(n_348),
.Y(n_389)
);

AO21x1_ASAP7_75t_L g421 ( 
.A1(n_389),
.A2(n_397),
.B(n_408),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_378),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_404),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_366),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_391),
.B(n_393),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_407),
.C(n_411),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_384),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_368),
.A2(n_335),
.B1(n_340),
.B2(n_328),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_372),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_403),
.Y(n_425)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_399),
.Y(n_418)
);

OAI22x1_ASAP7_75t_L g414 ( 
.A1(n_400),
.A2(n_371),
.B1(n_362),
.B2(n_363),
.Y(n_414)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_401),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_380),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_369),
.B(n_346),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_386),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_410),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_379),
.A2(n_346),
.B1(n_360),
.B2(n_354),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_367),
.A2(n_358),
.B1(n_355),
.B2(n_333),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_409),
.A2(n_371),
.B1(n_363),
.B2(n_374),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_386),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_365),
.B(n_373),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_382),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_412),
.B(n_370),
.Y(n_413)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_413),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_414),
.A2(n_419),
.B1(n_418),
.B2(n_422),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_373),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_406),
.Y(n_445)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_387),
.C(n_375),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_417),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_402),
.B(n_387),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_399),
.B(n_375),
.Y(n_422)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_422),
.Y(n_442)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_400),
.Y(n_426)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_426),
.Y(n_444)
);

OAI21xp33_ASAP7_75t_L g428 ( 
.A1(n_407),
.A2(n_388),
.B(n_374),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_428),
.A2(n_395),
.B1(n_397),
.B2(n_394),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_389),
.A2(n_367),
.B(n_376),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_431),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_408),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_390),
.C(n_365),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_435),
.C(n_439),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_401),
.C(n_411),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_421),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_426),
.A2(n_367),
.B1(n_409),
.B2(n_396),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_437),
.A2(n_423),
.B1(n_414),
.B2(n_419),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_429),
.C(n_432),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_377),
.C(n_406),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_440),
.B(n_421),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_443),
.B(n_430),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_446),
.B(n_443),
.Y(n_455)
);

BUFx24_ASAP7_75t_SL g447 ( 
.A(n_438),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_453),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_448),
.B(n_434),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_449),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_413),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_451),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_421),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_452),
.B(n_440),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_424),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_457),
.Y(n_466)
);

AO221x1_ASAP7_75t_L g457 ( 
.A1(n_451),
.A2(n_406),
.B1(n_417),
.B2(n_425),
.C(n_442),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_458),
.B(n_460),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_459),
.B(n_454),
.C(n_439),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_463),
.B(n_464),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_454),
.C(n_461),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_460),
.A2(n_427),
.B(n_456),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_465),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_455),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_467),
.B(n_466),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g472 ( 
.A1(n_470),
.A2(n_471),
.B(n_468),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_469),
.B(n_463),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_472),
.B(n_467),
.Y(n_473)
);

AOI211xp5_ASAP7_75t_SL g474 ( 
.A1(n_473),
.A2(n_445),
.B(n_418),
.C(n_431),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_437),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_444),
.Y(n_476)
);


endmodule