module real_jpeg_5393_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_0),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_0),
.Y(n_355)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_2),
.Y(n_110)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_2),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_3),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_3),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_3),
.B(n_83),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_3),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_3),
.B(n_112),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_3),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_3),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_3),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_4),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_4),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_4),
.B(n_301),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_4),
.B(n_357),
.Y(n_356)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_6),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_6),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_6),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_7),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_7),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_7),
.B(n_345),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_8),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_8),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_8),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_8),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_8),
.B(n_116),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_8),
.B(n_387),
.Y(n_386)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_9),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_9),
.Y(n_329)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_11),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_11),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_11),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_11),
.B(n_102),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_11),
.B(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_11),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_11),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_12),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_12),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_12),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_12),
.B(n_301),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_13),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_13),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_13),
.B(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_13),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_13),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_13),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_14),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_14),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_14),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_14),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_14),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_14),
.B(n_60),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g240 ( 
.A(n_15),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_15),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_15),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_15),
.B(n_401),
.Y(n_400)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_16),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_16),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_16),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_17),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_17),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_17),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_17),
.B(n_83),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_17),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_17),
.B(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_364),
.Y(n_18)
);

AOI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_319),
.B(n_363),
.Y(n_19)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_272),
.B(n_318),
.Y(n_20)
);

AOI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_230),
.B(n_271),
.Y(n_21)
);

AO21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_148),
.B(n_229),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_133),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_24),
.B(n_133),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_70),
.B2(n_132),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_25),
.B(n_71),
.C(n_113),
.Y(n_270)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_46),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_27),
.B(n_47),
.C(n_69),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_40),
.C(n_44),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_28),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_29),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_138)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_33),
.Y(n_155)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_33),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_33),
.Y(n_335)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_39),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_40),
.B(n_44),
.Y(n_147)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_42),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_42),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_43),
.Y(n_289)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_45),
.Y(n_299)
);

INVx3_ASAP7_75t_SL g396 ( 
.A(n_45),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_56),
.B1(n_68),
.B2(n_69),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_55),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_51),
.Y(n_55)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_55),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_55),
.B(n_235),
.C(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_57),
.B(n_62),
.C(n_66),
.Y(n_269)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_65),
.Y(n_296)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_65),
.Y(n_343)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_113),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_89),
.C(n_105),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_85),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_80),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_80),
.C(n_85),
.Y(n_131)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_77),
.Y(n_301)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_79),
.Y(n_203)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_84),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_86),
.Y(n_401)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_89),
.A2(n_90),
.B1(n_105),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_100),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_91),
.A2(n_92),
.B1(n_100),
.B2(n_101),
.Y(n_222)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_94),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_95),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_98),
.Y(n_257)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_107),
.B(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g308 ( 
.A(n_110),
.Y(n_308)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

XOR2x1_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_129),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_114),
.B(n_130),
.C(n_131),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_115),
.B(n_123),
.C(n_127),
.Y(n_248)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_123),
.B1(n_127),
.B2(n_128),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_122),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_123),
.Y(n_128)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_126),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_146),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_134),
.B(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_137),
.B(n_146),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.C(n_140),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_138),
.B(n_139),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_140),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_144),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_224),
.B(n_228),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_209),
.B(n_223),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_189),
.B(n_208),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_176),
.B(n_188),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_170),
.B2(n_171),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_166),
.C(n_170),
.Y(n_207)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_165),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_175),
.Y(n_193)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_183),
.B(n_187),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_179),
.Y(n_187)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_207),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_207),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_193),
.C(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_204),
.C(n_206),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_212),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_219),
.C(n_220),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_270),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_270),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_250),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_234),
.C(n_250),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_247),
.B2(n_249),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_253),
.C(n_263),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_259),
.C(n_260),
.Y(n_303)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_269),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_267),
.C(n_269),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_274),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_275),
.B(n_292),
.C(n_316),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_292),
.B1(n_316),
.B2(n_317),
.Y(n_276)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_277),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_291),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_284),
.B(n_287),
.C(n_290),
.Y(n_351)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx6_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_302),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_293),
.B(n_303),
.C(n_304),
.Y(n_349)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_293),
.Y(n_406)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_297),
.CI(n_300),
.CON(n_293),
.SN(n_293)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_294),
.B(n_297),
.C(n_300),
.Y(n_360)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_313),
.B2(n_314),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_306)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_312),
.C(n_313),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_309),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_309),
.A2(n_312),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_312),
.B(n_326),
.C(n_332),
.Y(n_378)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_362),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_320),
.B(n_362),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_321),
.B(n_323),
.C(n_347),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_347),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_336),
.B2(n_346),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_337),
.C(n_338),
.Y(n_372)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_331),
.A2(n_332),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_336),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_344),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_340),
.B(n_341),
.C(n_344),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.B1(n_350),
.B2(n_361),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_351),
.C(n_352),
.Y(n_368)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_350),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_360),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_356),
.B1(n_358),
.B2(n_359),
.Y(n_353)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_354),
.Y(n_358)
);

INVx8_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_356),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_358),
.C(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_359),
.B1(n_380),
.B2(n_383),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_360),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_404),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_403),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_403),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_384),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_377),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_380),
.Y(n_383)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_392),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_389),
.Y(n_385)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_397),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_399),
.B1(n_400),
.B2(n_402),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_398),
.Y(n_402)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);


endmodule