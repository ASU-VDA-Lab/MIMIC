module real_jpeg_26065_n_19 (n_17, n_123, n_8, n_116, n_0, n_2, n_10, n_114, n_9, n_12, n_124, n_6, n_121, n_11, n_14, n_7, n_117, n_18, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_16, n_15, n_13, n_120, n_19);

input n_17;
input n_123;
input n_8;
input n_116;
input n_0;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_124;
input n_6;
input n_121;
input n_11;
input n_14;
input n_7;
input n_117;
input n_18;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_16;
input n_15;
input n_13;
input n_120;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_0),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_1),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_3),
.B(n_98),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_4),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_33),
.C(n_111),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_6),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_6),
.B(n_35),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_7),
.B(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_8),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_8),
.B(n_95),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_9),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_10),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_11),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_13),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_13),
.B(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_15),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_15),
.B(n_64),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_18),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_28),
.B(n_46),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_28),
.B(n_107),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_29),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B(n_110),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_104),
.B(n_109),
.Y(n_38)
);

OAI321xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_94),
.A3(n_97),
.B1(n_102),
.B2(n_103),
.C(n_114),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_88),
.B(n_93),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_83),
.B(n_87),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_75),
.B(n_82),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B(n_74),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_67),
.B(n_73),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_63),
.B(n_66),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_55),
.B(n_62),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_69),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_77),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_96),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_90),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_108),
.Y(n_109)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_115),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_116),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_117),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_118),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_119),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_120),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_121),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_122),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_123),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_124),
.Y(n_101)
);


endmodule