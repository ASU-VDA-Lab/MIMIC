module fake_jpeg_15307_n_346 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_32),
.Y(n_62)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_16),
.B1(n_19),
.B2(n_26),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_36),
.B1(n_35),
.B2(n_27),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_54),
.B(n_58),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_26),
.B(n_22),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_30),
.B(n_18),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_19),
.B1(n_16),
.B2(n_27),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_65),
.A2(n_20),
.B1(n_32),
.B2(n_28),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_30),
.Y(n_114)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_37),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_19),
.B1(n_16),
.B2(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_102),
.B1(n_67),
.B2(n_74),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_86),
.A2(n_99),
.B1(n_113),
.B2(n_66),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_87),
.B(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_90),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_39),
.C(n_30),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_29),
.C(n_34),
.Y(n_126)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_97),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_30),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_47),
.B1(n_44),
.B2(n_24),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_17),
.B1(n_23),
.B2(n_20),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_10),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_55),
.A2(n_23),
.B(n_17),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_107),
.A2(n_111),
.B(n_32),
.Y(n_121)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_32),
.B1(n_28),
.B2(n_11),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_115),
.B(n_127),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_140),
.B1(n_112),
.B2(n_100),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g160 ( 
.A(n_121),
.B(n_144),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_99),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_77),
.Y(n_127)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_137),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_89),
.A2(n_68),
.B1(n_66),
.B2(n_61),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_85),
.B1(n_113),
.B2(n_109),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_78),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_21),
.C(n_29),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_25),
.C(n_34),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_21),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_87),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_146),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_85),
.B(n_80),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_137),
.B(n_132),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_149),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_135),
.B1(n_133),
.B2(n_125),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_91),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_151),
.B(n_159),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_153),
.A2(n_168),
.B1(n_105),
.B2(n_123),
.Y(n_200)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g157 ( 
.A(n_122),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_157),
.B(n_167),
.Y(n_212)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_93),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_174),
.C(n_29),
.Y(n_193)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_79),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_178),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_115),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_108),
.B1(n_61),
.B2(n_101),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_169),
.B(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_171),
.B(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_92),
.C(n_104),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_175),
.Y(n_180)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_133),
.Y(n_190)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_63),
.B(n_96),
.C(n_81),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_139),
.A3(n_144),
.B1(n_136),
.B2(n_119),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_181),
.B(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_185),
.B(n_148),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_187),
.A2(n_206),
.B1(n_149),
.B2(n_116),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_159),
.B(n_124),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_188),
.B(n_178),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_131),
.B1(n_125),
.B2(n_135),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_189),
.A2(n_198),
.B1(n_157),
.B2(n_155),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_166),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_195),
.B(n_148),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_199),
.C(n_207),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_200),
.B1(n_203),
.B2(n_1),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_0),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_82),
.B1(n_103),
.B2(n_123),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_104),
.C(n_34),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_149),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_116),
.B1(n_9),
.B2(n_10),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_25),
.C(n_21),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_25),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_213),
.Y(n_214)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_158),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_219),
.C(n_222),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_204),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_216),
.B(n_226),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_232),
.B1(n_239),
.B2(n_240),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_156),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_230),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_194),
.A2(n_208),
.B1(n_209),
.B2(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_175),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_173),
.B(n_163),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_224),
.B(n_231),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_197),
.Y(n_226)
);

INVxp33_ASAP7_75t_SL g228 ( 
.A(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_165),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_241),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_182),
.B(n_162),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_235),
.B(n_211),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_180),
.Y(n_250)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_208),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_186),
.B1(n_195),
.B2(n_196),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_1),
.B(n_2),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_8),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_229),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_214),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_185),
.B1(n_184),
.B2(n_238),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_222),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_257),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_181),
.B1(n_195),
.B2(n_187),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_254),
.A2(n_256),
.B1(n_230),
.B2(n_234),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_199),
.B1(n_189),
.B2(n_186),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_220),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_210),
.C(n_207),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_257),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_191),
.Y(n_261)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_275),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_227),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_271),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_SL g270 ( 
.A(n_265),
.B(n_212),
.C(n_219),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_227),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_221),
.B(n_241),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_277),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_217),
.B1(n_223),
.B2(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_184),
.B(n_8),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_255),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_7),
.B(n_13),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_284),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_248),
.A2(n_7),
.B(n_12),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_252),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_247),
.CI(n_253),
.CON(n_287),
.SN(n_287)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_258),
.C(n_247),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_299),
.C(n_300),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_259),
.C(n_243),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_259),
.C(n_242),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_269),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_260),
.C(n_3),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_14),
.C(n_3),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_306),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_275),
.B1(n_273),
.B2(n_272),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_291),
.B1(n_298),
.B2(n_303),
.Y(n_322)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_310),
.C(n_293),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_285),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_295),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_315),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_286),
.B1(n_277),
.B2(n_284),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_313),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_274),
.B1(n_282),
.B2(n_281),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_290),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_299),
.B(n_12),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_297),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_297),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_319),
.B(n_321),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_325),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_326),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_293),
.C(n_287),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_314),
.C(n_305),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_287),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_330),
.Y(n_335)
);

INVx11_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_327),
.A2(n_304),
.B1(n_307),
.B2(n_326),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_333),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_318),
.B(n_314),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_334),
.B(n_323),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_337),
.B(n_338),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_331),
.B(n_324),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_335),
.A2(n_332),
.B(n_328),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_339),
.A2(n_340),
.B(n_329),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_336),
.B(n_328),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_333),
.B(n_330),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_317),
.Y(n_346)
);


endmodule