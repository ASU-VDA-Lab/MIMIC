module fake_netlist_6_1453_n_2040 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2040);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2040;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1828;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx3_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_194),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_15),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_117),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_101),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_202),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_17),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_96),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_12),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_108),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_125),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_63),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_91),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_132),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_133),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_82),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_94),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_107),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_43),
.Y(n_231)
);

BUFx2_ASAP7_75t_SL g232 ( 
.A(n_10),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_113),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_29),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_148),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_169),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_11),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_157),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_119),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_49),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_189),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_87),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_188),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_167),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_32),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_8),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_121),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_25),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_43),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_147),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_111),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_21),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_19),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_49),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_80),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_61),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_23),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_155),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_154),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_65),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_128),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_142),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_162),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_110),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_196),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_165),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_13),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_57),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_67),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_105),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_59),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_86),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_6),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_152),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_124),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_38),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_122),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_6),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_32),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_47),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_71),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_71),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_173),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_176),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_90),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_114),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_30),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_14),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_68),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_186),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_67),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_140),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_53),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_183),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_34),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_103),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_134),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_143),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_33),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_93),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_127),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_38),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_52),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_136),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_52),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_14),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_68),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_131),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_77),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_184),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_47),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_198),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_60),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_89),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_16),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_145),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_179),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_95),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_37),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_54),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_168),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_56),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_208),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_109),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_149),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_88),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_164),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_37),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_78),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_175),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_17),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_156),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_72),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_181),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_69),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_115),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_178),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_160),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_100),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_27),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_104),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_3),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_54),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_63),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_150),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_44),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_126),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_29),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_61),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_83),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_62),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_19),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_75),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_33),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_123),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_191),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_3),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_0),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_57),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_177),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_166),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_48),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_51),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_65),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_182),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_135),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_144),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_130),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_159),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_75),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_11),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_60),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_45),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_73),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_139),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_102),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_197),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_97),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_201),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_79),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_15),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_204),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_27),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_116),
.Y(n_389)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_35),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_31),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_1),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_56),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_174),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_171),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_58),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_35),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_141),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_84),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_163),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_39),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_4),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_18),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_5),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_58),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_7),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_205),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_1),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_69),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_13),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_76),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_25),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_23),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_210),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_212),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_325),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_325),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_390),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_390),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_213),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_0),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_215),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_219),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_324),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_225),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_249),
.B(n_2),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g429 ( 
.A(n_378),
.B(n_2),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_226),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_390),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_390),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_383),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_233),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_228),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_390),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_229),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_383),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_390),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_324),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_324),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_324),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_240),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_279),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_289),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_230),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_334),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_324),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_324),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_221),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_227),
.B(n_5),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_221),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_209),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_236),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_237),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_243),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_356),
.B(n_9),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_244),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_251),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_268),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_251),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_245),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_268),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_248),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_255),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_255),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_263),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_263),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_252),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_295),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_295),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_336),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_261),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_336),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_313),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_209),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_313),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_265),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_267),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_376),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_222),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_350),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_365),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_376),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_235),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_235),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_269),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_238),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_238),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_254),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_214),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_254),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_211),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_274),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_256),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_276),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_256),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_270),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_270),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_227),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_271),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_287),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_271),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_209),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_302),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_303),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_305),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_314),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_242),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_239),
.B(n_9),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_319),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_272),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_232),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_272),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_283),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_283),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_285),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_415),
.Y(n_519)
);

XNOR2x2_ASAP7_75t_L g520 ( 
.A(n_452),
.B(n_333),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_461),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_434),
.A2(n_296),
.B1(n_316),
.B2(n_280),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_415),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_441),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_494),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g526 ( 
.A1(n_441),
.A2(n_286),
.B(n_285),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_442),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_454),
.B(n_260),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_442),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_419),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_449),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_419),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_449),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

BUFx8_ASAP7_75t_L g535 ( 
.A(n_477),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_450),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_450),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_440),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_426),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_420),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_438),
.B(n_214),
.Y(n_541)
);

CKINVDCx11_ASAP7_75t_R g542 ( 
.A(n_464),
.Y(n_542)
);

INVxp33_ASAP7_75t_L g543 ( 
.A(n_417),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_424),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_424),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_426),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_431),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_426),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_476),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_440),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_432),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_436),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_511),
.B(n_239),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_436),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_439),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_439),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_492),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_492),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_451),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_514),
.B(n_399),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_451),
.Y(n_563)
);

BUFx8_ASAP7_75t_L g564 ( 
.A(n_477),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_477),
.B(n_399),
.Y(n_565)
);

OA21x2_ASAP7_75t_L g566 ( 
.A1(n_422),
.A2(n_298),
.B(n_286),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_468),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_468),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_505),
.B(n_260),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_433),
.B(n_327),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_418),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_458),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_481),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_481),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_SL g575 ( 
.A(n_482),
.B(n_356),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_SL g576 ( 
.A(n_483),
.B(n_351),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_477),
.B(n_220),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_453),
.Y(n_578)
);

AND2x2_ASAP7_75t_SL g579 ( 
.A(n_484),
.B(n_220),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_453),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_460),
.Y(n_581)
);

OA21x2_ASAP7_75t_L g582 ( 
.A1(n_460),
.A2(n_300),
.B(n_298),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_501),
.B(n_438),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_477),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_462),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_462),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_414),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_466),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_466),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_467),
.B(n_327),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_467),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_SL g592 ( 
.A(n_445),
.B(n_377),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_469),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_469),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_471),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_471),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_472),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_472),
.B(n_473),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_473),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_475),
.B(n_354),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_475),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_577),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_555),
.A2(n_429),
.B1(n_408),
.B2(n_354),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_532),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_519),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_519),
.Y(n_606)
);

BUFx10_ASAP7_75t_L g607 ( 
.A(n_583),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_577),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_542),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_577),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_577),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_579),
.B(n_478),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_577),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_519),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_577),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_535),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_555),
.A2(n_409),
.B1(n_428),
.B2(n_224),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_579),
.B(n_416),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_532),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_520),
.A2(n_408),
.B1(n_300),
.B2(n_308),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_579),
.B(n_421),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_572),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_592),
.A2(n_231),
.B1(n_241),
.B2(n_216),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_519),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_579),
.B(n_510),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_535),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_541),
.B(n_485),
.Y(n_627)
);

AND3x2_ASAP7_75t_L g628 ( 
.A(n_572),
.B(n_395),
.C(n_297),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_535),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_583),
.B(n_484),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_523),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_520),
.A2(n_307),
.B1(n_310),
.B2(n_308),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_523),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_525),
.B(n_423),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_582),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_542),
.Y(n_636)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_576),
.Y(n_637)
);

AND3x2_ASAP7_75t_L g638 ( 
.A(n_587),
.B(n_297),
.C(n_223),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_582),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_541),
.B(n_485),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_528),
.B(n_425),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_525),
.B(n_427),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_582),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_523),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_541),
.B(n_486),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_528),
.B(n_430),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_571),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_523),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_582),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_582),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_532),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_535),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_532),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_530),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_530),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_532),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_541),
.B(n_486),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_570),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_530),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_582),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_582),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_571),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_528),
.B(n_435),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_532),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_569),
.B(n_437),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_569),
.B(n_232),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_569),
.B(n_447),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_551),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_551),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_587),
.B(n_455),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_570),
.B(n_456),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_532),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_570),
.B(n_487),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_532),
.Y(n_674)
);

INVx4_ASAP7_75t_SL g675 ( 
.A(n_532),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_534),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_530),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_551),
.B(n_457),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_587),
.B(n_218),
.Y(n_679)
);

HB1xp67_ASAP7_75t_SL g680 ( 
.A(n_521),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_566),
.B(n_218),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_521),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_562),
.A2(n_495),
.B1(n_508),
.B2(n_488),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_551),
.B(n_459),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_534),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_521),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_535),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_551),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_551),
.Y(n_689)
);

AO22x2_ASAP7_75t_L g690 ( 
.A1(n_520),
.A2(n_310),
.B1(n_311),
.B2(n_307),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_543),
.A2(n_247),
.B1(n_258),
.B2(n_246),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_566),
.B(n_234),
.C(n_223),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_534),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_540),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_562),
.B(n_463),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_540),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_540),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_584),
.B(n_465),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_540),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_543),
.B(n_470),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_534),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_544),
.Y(n_702)
);

AND2x6_ASAP7_75t_L g703 ( 
.A(n_544),
.B(n_234),
.Y(n_703)
);

CKINVDCx11_ASAP7_75t_R g704 ( 
.A(n_549),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_520),
.A2(n_273),
.B1(n_275),
.B2(n_259),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_584),
.B(n_474),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_584),
.B(n_479),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_534),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_592),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_575),
.A2(n_357),
.B1(n_362),
.B2(n_363),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_544),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_566),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_565),
.B(n_480),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_575),
.B(n_497),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_544),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_566),
.A2(n_512),
.B1(n_509),
.B2(n_503),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_552),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_552),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_535),
.B(n_506),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_564),
.B(n_507),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_576),
.Y(n_721)
);

AND2x6_ASAP7_75t_L g722 ( 
.A(n_552),
.B(n_250),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_586),
.B(n_501),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_552),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_598),
.B(n_487),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_584),
.B(n_501),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_549),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_556),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_556),
.B(n_558),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_564),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_598),
.B(n_489),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_534),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_564),
.B(n_501),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_564),
.Y(n_734)
);

NOR3xp33_ASAP7_75t_L g735 ( 
.A(n_522),
.B(n_549),
.C(n_299),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_534),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_564),
.B(n_242),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_556),
.B(n_217),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_534),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_556),
.B(n_315),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_534),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_564),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_558),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_586),
.B(n_443),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_586),
.B(n_444),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_545),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_545),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_558),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_558),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_561),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_561),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_L g752 ( 
.A1(n_566),
.A2(n_282),
.B1(n_284),
.B2(n_277),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_566),
.A2(n_311),
.B1(n_412),
.B2(n_403),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_565),
.B(n_343),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_658),
.B(n_590),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_622),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_622),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_602),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_656),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_750),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_641),
.B(n_566),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_632),
.A2(n_526),
.B1(n_349),
.B2(n_359),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_602),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_658),
.B(n_545),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_618),
.B(n_545),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_754),
.B(n_545),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_680),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_608),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_621),
.B(n_545),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_673),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_751),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_666),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_678),
.B(n_545),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_610),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_611),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_612),
.A2(n_446),
.B1(n_448),
.B2(n_352),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_611),
.B(n_545),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_613),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_684),
.B(n_545),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_613),
.B(n_547),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_615),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_654),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_673),
.B(n_547),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_646),
.B(n_291),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_615),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_627),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_712),
.B(n_663),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_725),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_L g789 ( 
.A(n_683),
.B(n_578),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_625),
.A2(n_326),
.B1(n_329),
.B2(n_322),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_712),
.B(n_547),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_665),
.B(n_547),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_667),
.B(n_547),
.Y(n_793)
);

BUFx5_ASAP7_75t_L g794 ( 
.A(n_616),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_671),
.B(n_547),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_713),
.B(n_547),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_713),
.B(n_547),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_634),
.B(n_292),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_723),
.B(n_547),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_627),
.Y(n_800)
);

NAND2x1_ASAP7_75t_L g801 ( 
.A(n_635),
.B(n_526),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_647),
.B(n_590),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_727),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_635),
.B(n_553),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_639),
.B(n_553),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_654),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_725),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_695),
.B(n_666),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_647),
.B(n_590),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_731),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_666),
.B(n_293),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_639),
.B(n_553),
.Y(n_812)
);

XOR2xp5_ASAP7_75t_L g813 ( 
.A(n_637),
.B(n_522),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_643),
.B(n_553),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_643),
.B(n_553),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_640),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_649),
.B(n_553),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_649),
.B(n_650),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_716),
.A2(n_331),
.B1(n_337),
.B2(n_330),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_650),
.B(n_660),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_656),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_660),
.B(n_553),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_661),
.B(n_553),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_654),
.Y(n_824)
);

BUFx6f_ASAP7_75t_SL g825 ( 
.A(n_607),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_731),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_661),
.B(n_553),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_666),
.A2(n_341),
.B1(n_342),
.B2(n_339),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_666),
.B(n_304),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_752),
.B(n_554),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_617),
.B(n_312),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_655),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_655),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_692),
.B(n_616),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_744),
.A2(n_355),
.B1(n_361),
.B2(n_346),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_745),
.A2(n_366),
.B1(n_371),
.B2(n_373),
.Y(n_836)
);

INVx5_ASAP7_75t_L g837 ( 
.A(n_681),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_655),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_659),
.Y(n_839)
);

NOR2xp67_ASAP7_75t_L g840 ( 
.A(n_692),
.B(n_578),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_659),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_656),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_738),
.B(n_554),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_740),
.B(n_554),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_616),
.B(n_626),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_640),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_662),
.B(n_522),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_645),
.B(n_554),
.Y(n_848)
);

NAND3xp33_ASAP7_75t_L g849 ( 
.A(n_620),
.B(n_603),
.C(n_623),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_626),
.B(n_554),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_645),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_657),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_626),
.B(n_554),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_657),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_668),
.B(n_669),
.Y(n_855)
);

OAI21xp33_ASAP7_75t_L g856 ( 
.A1(n_623),
.A2(n_600),
.B(n_349),
.Y(n_856)
);

AND2x6_ASAP7_75t_L g857 ( 
.A(n_629),
.B(n_250),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_668),
.B(n_554),
.Y(n_858)
);

BUFx6f_ASAP7_75t_SL g859 ( 
.A(n_607),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_669),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_659),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_688),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_642),
.B(n_318),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_677),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_688),
.B(n_554),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_689),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_677),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_677),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_679),
.A2(n_407),
.B1(n_380),
.B2(n_389),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_711),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_630),
.B(n_320),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_656),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_711),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_727),
.B(n_600),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_629),
.B(n_652),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_607),
.B(n_700),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_753),
.B(n_554),
.Y(n_877)
);

BUFx5_ASAP7_75t_L g878 ( 
.A(n_629),
.Y(n_878)
);

AOI221xp5_ASAP7_75t_L g879 ( 
.A1(n_705),
.A2(n_369),
.B1(n_364),
.B2(n_340),
.C(n_359),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_681),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_711),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_681),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_681),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_681),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_696),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_698),
.B(n_557),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_696),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_652),
.B(n_557),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_706),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_656),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_743),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_L g892 ( 
.A(n_707),
.B(n_737),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_682),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_652),
.B(n_557),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_679),
.A2(n_374),
.B1(n_382),
.B2(n_384),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_709),
.B(n_262),
.C(n_253),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_679),
.A2(n_400),
.B1(n_398),
.B2(n_387),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_743),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_679),
.A2(n_385),
.B1(n_526),
.B2(n_262),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_709),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_607),
.B(n_338),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_686),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_651),
.B(n_557),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_691),
.B(n_670),
.Y(n_904)
);

NAND2xp33_ASAP7_75t_SL g905 ( 
.A(n_714),
.B(n_345),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_702),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_743),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_679),
.B(n_347),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_L g909 ( 
.A(n_735),
.B(n_353),
.C(n_348),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_702),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_L g911 ( 
.A(n_726),
.B(n_253),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_715),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_704),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_719),
.A2(n_526),
.B1(n_332),
.B2(n_328),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_651),
.B(n_557),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_651),
.B(n_557),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_721),
.B(n_358),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_651),
.B(n_557),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_637),
.B(n_266),
.C(n_264),
.Y(n_919)
);

AO21x1_ASAP7_75t_L g920 ( 
.A1(n_830),
.A2(n_733),
.B(n_720),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_758),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_763),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_818),
.A2(n_730),
.B(n_687),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_798),
.B(n_710),
.Y(n_924)
);

NOR2x1_ASAP7_75t_R g925 ( 
.A(n_767),
.B(n_367),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_820),
.A2(n_730),
.B(n_687),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_787),
.A2(n_729),
.B(n_749),
.C(n_718),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_802),
.B(n_710),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_808),
.A2(n_904),
.B1(n_798),
.B2(n_761),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_796),
.A2(n_730),
.B(n_687),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_808),
.A2(n_690),
.B1(n_664),
.B2(n_672),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_797),
.A2(n_742),
.B(n_734),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_770),
.B(n_734),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_759),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_768),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_852),
.B(n_653),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_900),
.B(n_756),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_761),
.A2(n_749),
.B(n_718),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_809),
.B(n_690),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_852),
.B(n_653),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_787),
.A2(n_748),
.B(n_715),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_904),
.A2(n_266),
.B(n_278),
.C(n_264),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_876),
.B(n_755),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_886),
.A2(n_742),
.B(n_734),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_791),
.A2(n_742),
.B(n_619),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_889),
.B(n_653),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_759),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_774),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_791),
.A2(n_619),
.B(n_604),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_889),
.B(n_653),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_837),
.A2(n_690),
.B1(n_281),
.B2(n_288),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_876),
.B(n_656),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_784),
.B(n_664),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_784),
.B(n_664),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_837),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_880),
.A2(n_690),
.B1(n_672),
.B2(n_685),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_R g957 ( 
.A(n_905),
.B(n_609),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_759),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_786),
.B(n_664),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_851),
.B(n_600),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_800),
.B(n_816),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_792),
.A2(n_619),
.B(n_604),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_775),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_SL g964 ( 
.A(n_893),
.B(n_902),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_803),
.Y(n_965)
);

BUFx12f_ASAP7_75t_L g966 ( 
.A(n_913),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_759),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_821),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_773),
.A2(n_619),
.B(n_604),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_917),
.B(n_636),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_788),
.B(n_672),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_778),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_779),
.A2(n_674),
.B(n_604),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_917),
.B(n_628),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_807),
.B(n_672),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_849),
.A2(n_278),
.B(n_281),
.C(n_288),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_877),
.A2(n_697),
.B(n_694),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_810),
.B(n_685),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_826),
.B(n_685),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_783),
.A2(n_697),
.B(n_694),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_781),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_831),
.A2(n_748),
.B(n_699),
.C(n_717),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_831),
.A2(n_699),
.B(n_717),
.C(n_724),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_837),
.B(n_526),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_785),
.B(n_685),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_848),
.A2(n_795),
.B(n_793),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_793),
.A2(n_728),
.B(n_724),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_795),
.A2(n_728),
.B(n_674),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_896),
.A2(n_703),
.B1(n_722),
.B2(n_290),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_801),
.A2(n_606),
.B(n_605),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_854),
.A2(n_394),
.B(n_294),
.C(n_301),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_846),
.B(n_701),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_874),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_804),
.A2(n_614),
.B(n_606),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_766),
.A2(n_736),
.B(n_674),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_900),
.B(n_638),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_789),
.B(n_586),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_756),
.B(n_757),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_762),
.B(n_701),
.Y(n_999)
);

AO21x1_ASAP7_75t_L g1000 ( 
.A1(n_830),
.A2(n_294),
.B(n_290),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_843),
.A2(n_736),
.B(n_674),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_757),
.B(n_736),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_L g1003 ( 
.A(n_835),
.B(n_489),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_860),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_762),
.B(n_764),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_805),
.A2(n_624),
.B(n_614),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_862),
.Y(n_1007)
);

AOI21x1_ASAP7_75t_L g1008 ( 
.A1(n_765),
.A2(n_631),
.B(n_624),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_901),
.B(n_701),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_812),
.A2(n_633),
.B(n_631),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_844),
.A2(n_736),
.B(n_644),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_856),
.A2(n_323),
.B(n_394),
.C(n_381),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_821),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_814),
.A2(n_644),
.B(n_633),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_901),
.B(n_701),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_866),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_815),
.A2(n_648),
.B(n_708),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_817),
.A2(n_648),
.B(n_708),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_840),
.B(n_708),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_765),
.A2(n_527),
.B(n_524),
.Y(n_1020)
);

AND2x6_ASAP7_75t_L g1021 ( 
.A(n_882),
.B(n_883),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_822),
.A2(n_732),
.B(n_708),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_896),
.B(n_732),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_776),
.B(n_732),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_837),
.B(n_242),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_823),
.B(n_732),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_L g1027 ( 
.A(n_794),
.B(n_703),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_863),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_827),
.A2(n_741),
.B(n_739),
.Y(n_1029)
);

CKINVDCx10_ASAP7_75t_R g1030 ( 
.A(n_825),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_871),
.B(n_739),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_769),
.A2(n_741),
.B(n_739),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_871),
.B(n_739),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_855),
.B(n_741),
.Y(n_1034)
);

AO21x1_ASAP7_75t_L g1035 ( 
.A1(n_769),
.A2(n_892),
.B(n_834),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_772),
.B(n_598),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_885),
.B(n_741),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_887),
.B(n_746),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_906),
.B(n_746),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_821),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_884),
.A2(n_323),
.B1(n_309),
.B2(n_381),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_834),
.A2(n_747),
.B(n_746),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_777),
.A2(n_747),
.B(n_746),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_777),
.A2(n_747),
.B(n_722),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_910),
.B(n_747),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_912),
.B(n_703),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_863),
.B(n_703),
.Y(n_1047)
);

BUFx4f_ASAP7_75t_L g1048 ( 
.A(n_847),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_811),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_760),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_879),
.A2(n_370),
.B(n_332),
.C(n_328),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_908),
.B(n_598),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_799),
.B(n_703),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_908),
.B(n_703),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_780),
.A2(n_722),
.B(n_703),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_811),
.B(n_722),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_780),
.A2(n_693),
.B(n_676),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_821),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_858),
.A2(n_693),
.B(n_676),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_865),
.A2(n_915),
.B(n_903),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_850),
.A2(n_370),
.B(n_309),
.C(n_306),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_842),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_829),
.B(n_722),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_829),
.A2(n_772),
.B1(n_911),
.B2(n_819),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_916),
.A2(n_722),
.B(n_526),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_842),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_918),
.A2(n_693),
.B(n_676),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_SL g1068 ( 
.A(n_825),
.B(n_242),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_850),
.A2(n_693),
.B(n_676),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_853),
.A2(n_693),
.B(n_676),
.Y(n_1070)
);

BUFx4f_ASAP7_75t_L g1071 ( 
.A(n_857),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_919),
.B(n_490),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_842),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_909),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_853),
.A2(n_693),
.B(n_676),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_914),
.B(n_722),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_888),
.A2(n_557),
.B(n_559),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_782),
.B(n_526),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_888),
.A2(n_557),
.B(n_559),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_842),
.Y(n_1080)
);

INVx11_ASAP7_75t_L g1081 ( 
.A(n_857),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_806),
.B(n_675),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_894),
.A2(n_560),
.B(n_559),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_919),
.B(n_490),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_794),
.B(n_257),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_899),
.A2(n_301),
.B(n_344),
.C(n_306),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_L g1087 ( 
.A(n_794),
.B(n_317),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_894),
.A2(n_875),
.B(n_845),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_869),
.A2(n_317),
.B1(n_321),
.B2(n_335),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_824),
.B(n_675),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_832),
.A2(n_546),
.B(n_539),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_833),
.B(n_675),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_771),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_845),
.A2(n_546),
.B(n_539),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_794),
.B(n_257),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_838),
.B(n_675),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_839),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_828),
.A2(n_360),
.B(n_344),
.C(n_321),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_L g1099 ( 
.A(n_836),
.B(n_375),
.C(n_368),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_841),
.B(n_675),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_890),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_861),
.A2(n_539),
.B(n_546),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_895),
.A2(n_548),
.B1(n_560),
.B2(n_533),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_864),
.B(n_585),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_867),
.A2(n_548),
.B(n_527),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_875),
.A2(n_560),
.B(n_537),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_993),
.B(n_965),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_924),
.A2(n_897),
.B1(n_859),
.B2(n_790),
.Y(n_1108)
);

BUFx12f_ASAP7_75t_L g1109 ( 
.A(n_966),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1048),
.Y(n_1110)
);

BUFx4f_ASAP7_75t_L g1111 ( 
.A(n_1021),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_921),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1028),
.A2(n_859),
.B1(n_813),
.B2(n_857),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_952),
.A2(n_1015),
.B(n_1009),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_929),
.A2(n_872),
.B1(n_890),
.B2(n_340),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_922),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1027),
.A2(n_890),
.B(n_878),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1024),
.A2(n_907),
.B(n_898),
.C(n_891),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1005),
.B(n_872),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1087),
.A2(n_890),
.B(n_878),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1048),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1052),
.B(n_868),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_930),
.A2(n_873),
.B(n_870),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_928),
.A2(n_857),
.B1(n_881),
.B2(n_257),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1049),
.B(n_794),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_1088),
.A2(n_1064),
.B(n_943),
.C(n_1074),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_986),
.A2(n_857),
.B(n_536),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1099),
.A2(n_878),
.B1(n_794),
.B2(n_372),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_953),
.A2(n_878),
.B(n_561),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_935),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_930),
.A2(n_529),
.B(n_524),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_972),
.B(n_960),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_970),
.B(n_491),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_936),
.B(n_878),
.Y(n_1134)
);

NOR3xp33_ASAP7_75t_SL g1135 ( 
.A(n_937),
.B(n_413),
.C(n_411),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_948),
.B(n_878),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_SL g1137 ( 
.A(n_1068),
.B(n_410),
.C(n_379),
.Y(n_1137)
);

NAND2xp33_ASAP7_75t_SL g1138 ( 
.A(n_957),
.B(n_364),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1036),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_939),
.B(n_491),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_SL g1141 ( 
.A(n_964),
.B(n_257),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_R g1142 ( 
.A(n_1030),
.B(n_974),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1088),
.A2(n_369),
.B(n_386),
.C(n_412),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_996),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_R g1145 ( 
.A(n_1036),
.B(n_1054),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1072),
.B(n_493),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_961),
.B(n_372),
.Y(n_1147)
);

NOR2xp67_ASAP7_75t_SL g1148 ( 
.A(n_955),
.B(n_386),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_954),
.A2(n_561),
.B(n_563),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_963),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_981),
.B(n_1084),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_958),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1002),
.B(n_578),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_998),
.B(n_388),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1003),
.B(n_493),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_955),
.B(n_372),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1004),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_962),
.A2(n_563),
.B(n_568),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_925),
.B(n_391),
.Y(n_1159)
);

INVx3_ASAP7_75t_SL g1160 ( 
.A(n_1025),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1021),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1007),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1008),
.A2(n_585),
.B(n_597),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1016),
.B(n_372),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_956),
.B(n_396),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_940),
.B(n_580),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1031),
.A2(n_563),
.B(n_568),
.Y(n_1167)
);

BUFx12f_ASAP7_75t_L g1168 ( 
.A(n_1021),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1033),
.A2(n_563),
.B(n_568),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_969),
.A2(n_568),
.B(n_537),
.Y(n_1170)
);

BUFx12f_ASAP7_75t_L g1171 ( 
.A(n_1021),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_R g1172 ( 
.A(n_934),
.B(n_402),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1021),
.B(n_1093),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1089),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1097),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_931),
.B(n_585),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1047),
.A2(n_392),
.B(n_397),
.C(n_401),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_971),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_958),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_999),
.B(n_585),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_SL g1181 ( 
.A1(n_920),
.A2(n_392),
.B(n_397),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_951),
.A2(n_404),
.B1(n_405),
.B2(n_406),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_946),
.B(n_401),
.Y(n_1183)
);

BUFx12f_ASAP7_75t_L g1184 ( 
.A(n_958),
.Y(n_1184)
);

BUFx8_ASAP7_75t_L g1185 ( 
.A(n_1050),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_942),
.A2(n_403),
.B(n_496),
.C(n_498),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_L g1187 ( 
.A(n_1056),
.B(n_1063),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_967),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_973),
.A2(n_537),
.B(n_536),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_950),
.B(n_585),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_975),
.B(n_585),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_L g1192 ( 
.A(n_1051),
.B(n_1098),
.C(n_1041),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_976),
.A2(n_496),
.B(n_498),
.C(n_499),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_978),
.B(n_597),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_967),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_SL g1196 ( 
.A1(n_989),
.A2(n_517),
.B1(n_500),
.B2(n_502),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1026),
.A2(n_531),
.B(n_536),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_986),
.A2(n_524),
.B(n_527),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_959),
.B(n_10),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_979),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1086),
.A2(n_1071),
.B1(n_1023),
.B2(n_1076),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_992),
.B(n_597),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1034),
.B(n_597),
.Y(n_1203)
);

AOI33xp33_ASAP7_75t_L g1204 ( 
.A1(n_1012),
.A2(n_499),
.A3(n_500),
.B1(n_502),
.B2(n_504),
.B3(n_513),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_938),
.A2(n_529),
.B(n_531),
.Y(n_1205)
);

NOR3xp33_ASAP7_75t_SL g1206 ( 
.A(n_991),
.B(n_504),
.C(n_513),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1042),
.A2(n_597),
.B(n_533),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_997),
.B(n_12),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_995),
.A2(n_533),
.B(n_531),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_995),
.A2(n_529),
.B(n_538),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_967),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1035),
.B(n_597),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_933),
.B(n_16),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1001),
.A2(n_945),
.B(n_949),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1078),
.B(n_581),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1042),
.A2(n_550),
.B(n_580),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1060),
.B(n_581),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_968),
.B(n_580),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_982),
.A2(n_601),
.B(n_588),
.C(n_596),
.Y(n_1219)
);

INVx4_ASAP7_75t_L g1220 ( 
.A(n_968),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_968),
.B(n_515),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_934),
.B(n_581),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_947),
.B(n_581),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1085),
.A2(n_516),
.B(n_517),
.C(n_518),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_947),
.B(n_593),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1104),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1013),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1095),
.A2(n_516),
.B(n_518),
.C(n_596),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1058),
.B(n_593),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1013),
.B(n_1040),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_983),
.A2(n_601),
.B(n_588),
.C(n_596),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1013),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1058),
.B(n_593),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1073),
.B(n_593),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1017),
.A2(n_550),
.B(n_588),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1040),
.B(n_1062),
.Y(n_1236)
);

NAND3xp33_ASAP7_75t_SL g1237 ( 
.A(n_1000),
.B(n_601),
.C(n_591),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1001),
.A2(n_538),
.B(n_574),
.Y(n_1238)
);

OAI21xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1018),
.A2(n_595),
.B(n_594),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1046),
.A2(n_595),
.B(n_594),
.C(n_591),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1053),
.A2(n_538),
.B(n_574),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1037),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1038),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_985),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1039),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1019),
.B(n_18),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1045),
.B(n_20),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1073),
.B(n_21),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_984),
.B(n_1040),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1020),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1017),
.B(n_1014),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_984),
.B(n_22),
.Y(n_1252)
);

INVx5_ASAP7_75t_L g1253 ( 
.A(n_1062),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1103),
.Y(n_1254)
);

CKINVDCx8_ASAP7_75t_R g1255 ( 
.A(n_1062),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1066),
.B(n_22),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1066),
.B(n_24),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1071),
.A2(n_595),
.B1(n_594),
.B2(n_591),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1066),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_R g1260 ( 
.A(n_1080),
.B(n_85),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1080),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_944),
.A2(n_932),
.B(n_1011),
.Y(n_1262)
);

NAND2x1p5_ASAP7_75t_L g1263 ( 
.A(n_1080),
.B(n_574),
.Y(n_1263)
);

INVx5_ASAP7_75t_L g1264 ( 
.A(n_1101),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1262),
.A2(n_932),
.A3(n_923),
.B(n_926),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1163),
.A2(n_987),
.B(n_1014),
.Y(n_1266)
);

OR2x6_ASAP7_75t_L g1267 ( 
.A(n_1168),
.B(n_1101),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1216),
.A2(n_987),
.B(n_980),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1214),
.A2(n_926),
.B(n_923),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1126),
.A2(n_980),
.B(n_977),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1133),
.B(n_1106),
.Y(n_1271)
);

AOI221x1_ASAP7_75t_L g1272 ( 
.A1(n_1181),
.A2(n_1106),
.B1(n_1011),
.B2(n_1032),
.C(n_941),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1235),
.A2(n_977),
.B(n_1029),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1109),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1184),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1146),
.B(n_1029),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1154),
.B(n_1101),
.Y(n_1277)
);

AO32x2_ASAP7_75t_L g1278 ( 
.A1(n_1115),
.A2(n_1061),
.A3(n_927),
.B1(n_1065),
.B2(n_1010),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1173),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1110),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1187),
.A2(n_1022),
.B(n_1032),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1116),
.Y(n_1282)
);

INVx3_ASAP7_75t_SL g1283 ( 
.A(n_1107),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1201),
.A2(n_988),
.B(n_1083),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1251),
.A2(n_988),
.A3(n_1094),
.B(n_1079),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_SL g1286 ( 
.A1(n_1176),
.A2(n_1055),
.B(n_1094),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1134),
.A2(n_1117),
.B(n_1251),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1108),
.A2(n_1081),
.B1(n_1090),
.B2(n_1100),
.Y(n_1288)
);

AOI221x1_ASAP7_75t_L g1289 ( 
.A1(n_1201),
.A2(n_1077),
.B1(n_1006),
.B2(n_994),
.C(n_1105),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1121),
.B(n_1044),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1185),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1151),
.B(n_1043),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1134),
.A2(n_990),
.B(n_1102),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1120),
.A2(n_1091),
.B(n_1043),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1129),
.A2(n_1096),
.B(n_1092),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1132),
.B(n_567),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1255),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1140),
.B(n_1082),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1130),
.Y(n_1299)
);

AOI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1131),
.A2(n_1059),
.B(n_1067),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1192),
.A2(n_1069),
.B(n_1059),
.C(n_1075),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1123),
.A2(n_1067),
.B(n_1069),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1147),
.A2(n_573),
.B(n_567),
.C(n_599),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1207),
.A2(n_1070),
.B(n_1057),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1158),
.A2(n_1057),
.B(n_550),
.Y(n_1305)
);

AO21x1_ASAP7_75t_L g1306 ( 
.A1(n_1115),
.A2(n_573),
.B(n_567),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1165),
.A2(n_599),
.B(n_573),
.C(n_538),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1238),
.A2(n_599),
.B(n_538),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1246),
.A2(n_599),
.B(n_589),
.C(n_28),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1254),
.A2(n_589),
.B(n_26),
.C(n_28),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1174),
.B(n_24),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1127),
.A2(n_589),
.B(n_206),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1127),
.A2(n_589),
.B(n_195),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1185),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1239),
.A2(n_589),
.B(n_192),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1183),
.B(n_589),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1150),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1171),
.B(n_589),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1217),
.A2(n_589),
.B(n_190),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1157),
.Y(n_1320)
);

INVx4_ASAP7_75t_L g1321 ( 
.A(n_1253),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1139),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1144),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1217),
.A2(n_589),
.B(n_187),
.Y(n_1324)
);

OAI22x1_ASAP7_75t_L g1325 ( 
.A1(n_1113),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_1325)
);

AOI221x1_ASAP7_75t_L g1326 ( 
.A1(n_1143),
.A2(n_1177),
.B1(n_1252),
.B2(n_1247),
.C(n_1199),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1208),
.A2(n_34),
.B1(n_36),
.B2(n_39),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1119),
.A2(n_1153),
.B(n_1166),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1162),
.Y(n_1329)
);

NOR4xp25_ASAP7_75t_L g1330 ( 
.A(n_1186),
.B(n_40),
.C(n_41),
.D(n_42),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1210),
.A2(n_185),
.B(n_180),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1119),
.A2(n_1215),
.B(n_1136),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1170),
.A2(n_170),
.B(n_161),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1215),
.A2(n_158),
.B(n_151),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1142),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1152),
.Y(n_1336)
);

NOR4xp25_ASAP7_75t_L g1337 ( 
.A(n_1137),
.B(n_40),
.C(n_41),
.D(n_42),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1155),
.B(n_44),
.Y(n_1338)
);

INVx8_ASAP7_75t_L g1339 ( 
.A(n_1253),
.Y(n_1339)
);

AOI221xp5_ASAP7_75t_L g1340 ( 
.A1(n_1138),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.C(n_50),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1141),
.B(n_46),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1203),
.A2(n_146),
.B(n_138),
.Y(n_1342)
);

A2O1A1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1213),
.A2(n_50),
.B(n_51),
.C(n_53),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1128),
.A2(n_55),
.B(n_59),
.C(n_62),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1175),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_1221),
.B(n_92),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1206),
.A2(n_55),
.B(n_64),
.C(n_66),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1160),
.B(n_64),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1182),
.B(n_70),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1164),
.B(n_73),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1167),
.A2(n_106),
.B(n_129),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1161),
.B(n_137),
.Y(n_1352)
);

AOI221x1_ASAP7_75t_L g1353 ( 
.A1(n_1248),
.A2(n_74),
.B1(n_76),
.B2(n_81),
.C(n_98),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1172),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1212),
.A2(n_74),
.A3(n_99),
.B(n_112),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1169),
.A2(n_118),
.B(n_120),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1250),
.A2(n_1219),
.A3(n_1209),
.B(n_1118),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1149),
.A2(n_1189),
.B(n_1198),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1135),
.Y(n_1359)
);

AO22x2_ASAP7_75t_L g1360 ( 
.A1(n_1176),
.A2(n_1178),
.B1(n_1200),
.B2(n_1156),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1203),
.A2(n_1125),
.B(n_1122),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1244),
.B(n_1242),
.Y(n_1362)
);

AO21x1_ASAP7_75t_L g1363 ( 
.A1(n_1180),
.A2(n_1198),
.B(n_1145),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1224),
.Y(n_1364)
);

OA22x2_ASAP7_75t_L g1365 ( 
.A1(n_1221),
.A2(n_1259),
.B1(n_1236),
.B2(n_1230),
.Y(n_1365)
);

NOR2xp67_ASAP7_75t_SL g1366 ( 
.A(n_1253),
.B(n_1264),
.Y(n_1366)
);

A2O1A1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1124),
.A2(n_1111),
.B(n_1204),
.C(n_1258),
.Y(n_1367)
);

AO32x2_ASAP7_75t_L g1368 ( 
.A1(n_1196),
.A2(n_1220),
.A3(n_1211),
.B1(n_1114),
.B2(n_1205),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1256),
.A2(n_1257),
.B1(n_1243),
.B2(n_1245),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1195),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1241),
.A2(n_1190),
.B(n_1180),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1111),
.A2(n_1240),
.B(n_1226),
.C(n_1228),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1231),
.A2(n_1173),
.B(n_1249),
.C(n_1193),
.Y(n_1373)
);

AO32x2_ASAP7_75t_L g1374 ( 
.A1(n_1211),
.A2(n_1220),
.A3(n_1205),
.B1(n_1237),
.B2(n_1148),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1227),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1152),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1190),
.A2(n_1202),
.B(n_1194),
.Y(n_1377)
);

AOI31xp67_ASAP7_75t_L g1378 ( 
.A1(n_1191),
.A2(n_1202),
.A3(n_1194),
.B(n_1223),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1159),
.A2(n_1260),
.B1(n_1264),
.B2(n_1188),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1218),
.A2(n_1191),
.B1(n_1229),
.B2(n_1234),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1152),
.B(n_1179),
.Y(n_1381)
);

AOI21x1_ASAP7_75t_SL g1382 ( 
.A1(n_1222),
.A2(n_1234),
.B(n_1223),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1179),
.B(n_1188),
.Y(n_1383)
);

OAI21xp33_ASAP7_75t_L g1384 ( 
.A1(n_1222),
.A2(n_1233),
.B(n_1225),
.Y(n_1384)
);

AO21x1_ASAP7_75t_L g1385 ( 
.A1(n_1197),
.A2(n_1263),
.B(n_1225),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_SL g1386 ( 
.A1(n_1229),
.A2(n_1233),
.B(n_1263),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1264),
.A2(n_1179),
.B(n_1188),
.Y(n_1387)
);

AO31x2_ASAP7_75t_L g1388 ( 
.A1(n_1264),
.A2(n_1232),
.A3(n_1261),
.B(n_920),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1232),
.B(n_1261),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1232),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1261),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_SL g1392 ( 
.A(n_1141),
.B(n_924),
.C(n_798),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1163),
.A2(n_1216),
.B(n_1235),
.Y(n_1393)
);

NAND2x1_ASAP7_75t_L g1394 ( 
.A(n_1211),
.B(n_955),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1108),
.A2(n_924),
.B1(n_929),
.B2(n_1028),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1141),
.A2(n_924),
.B1(n_1048),
.B2(n_1174),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_SL g1397 ( 
.A1(n_1126),
.A2(n_924),
.B(n_976),
.C(n_942),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1214),
.A2(n_626),
.B(n_616),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1214),
.A2(n_626),
.B(n_616),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1126),
.A2(n_929),
.B(n_924),
.Y(n_1400)
);

NOR4xp25_ASAP7_75t_L g1401 ( 
.A(n_1126),
.B(n_924),
.C(n_942),
.D(n_1012),
.Y(n_1401)
);

NOR2xp67_ASAP7_75t_L g1402 ( 
.A(n_1151),
.B(n_1074),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1126),
.A2(n_929),
.B(n_924),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1112),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1146),
.B(n_924),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1163),
.A2(n_1216),
.B(n_1235),
.Y(n_1406)
);

AO22x1_ASAP7_75t_SL g1407 ( 
.A1(n_1254),
.A2(n_356),
.B1(n_238),
.B2(n_254),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1262),
.A2(n_1251),
.B(n_1198),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1214),
.A2(n_626),
.B(n_616),
.Y(n_1409)
);

OAI222xp33_ASAP7_75t_L g1410 ( 
.A1(n_1174),
.A2(n_924),
.B1(n_929),
.B2(n_617),
.C1(n_819),
.C2(n_632),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1146),
.B(n_924),
.Y(n_1411)
);

O2A1O1Ixp5_ASAP7_75t_SL g1412 ( 
.A1(n_1147),
.A2(n_737),
.B(n_952),
.C(n_630),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1110),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1108),
.A2(n_924),
.B(n_929),
.C(n_904),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1146),
.B(n_924),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1112),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1108),
.A2(n_924),
.B(n_929),
.C(n_904),
.Y(n_1417)
);

OAI21xp33_ASAP7_75t_L g1418 ( 
.A1(n_1154),
.A2(n_924),
.B(n_798),
.Y(n_1418)
);

AO31x2_ASAP7_75t_L g1419 ( 
.A1(n_1262),
.A2(n_920),
.A3(n_1000),
.B(n_1035),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1214),
.A2(n_626),
.B(n_616),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1126),
.A2(n_929),
.B(n_924),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1126),
.A2(n_929),
.B(n_924),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1110),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1107),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1335),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1418),
.A2(n_1414),
.B1(n_1417),
.B2(n_1396),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1339),
.Y(n_1427)
);

OAI22x1_ASAP7_75t_L g1428 ( 
.A1(n_1327),
.A2(n_1369),
.B1(n_1311),
.B2(n_1350),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1283),
.Y(n_1429)
);

OAI22x1_ASAP7_75t_L g1430 ( 
.A1(n_1327),
.A2(n_1369),
.B1(n_1341),
.B2(n_1277),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1404),
.Y(n_1431)
);

BUFx12f_ASAP7_75t_L g1432 ( 
.A(n_1274),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1418),
.A2(n_1392),
.B1(n_1395),
.B2(n_1415),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_L g1434 ( 
.A(n_1275),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1400),
.A2(n_1403),
.B1(n_1422),
.B2(n_1421),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1416),
.Y(n_1436)
);

BUFx2_ASAP7_75t_SL g1437 ( 
.A(n_1297),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1400),
.A2(n_1421),
.B1(n_1403),
.B2(n_1422),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1326),
.A2(n_1411),
.B(n_1405),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1349),
.A2(n_1313),
.B1(n_1312),
.B2(n_1346),
.Y(n_1440)
);

BUFx12f_ASAP7_75t_L g1441 ( 
.A(n_1275),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1340),
.A2(n_1325),
.B1(n_1313),
.B2(n_1312),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1402),
.A2(n_1271),
.B1(n_1348),
.B2(n_1346),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1362),
.B(n_1329),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1346),
.A2(n_1410),
.B1(n_1315),
.B2(n_1359),
.Y(n_1445)
);

BUFx12f_ASAP7_75t_L g1446 ( 
.A(n_1275),
.Y(n_1446)
);

INVx11_ASAP7_75t_L g1447 ( 
.A(n_1297),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1315),
.A2(n_1338),
.B1(n_1276),
.B2(n_1363),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1424),
.Y(n_1449)
);

BUFx4f_ASAP7_75t_SL g1450 ( 
.A(n_1291),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1317),
.A2(n_1320),
.B1(n_1345),
.B2(n_1360),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1339),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1360),
.A2(n_1292),
.B1(n_1364),
.B2(n_1299),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1354),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1365),
.A2(n_1423),
.B1(n_1413),
.B2(n_1280),
.Y(n_1455)
);

OAI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1353),
.A2(n_1298),
.B1(n_1296),
.B2(n_1314),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1370),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1379),
.A2(n_1323),
.B1(n_1375),
.B2(n_1372),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1352),
.A2(n_1290),
.B1(n_1322),
.B2(n_1284),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1366),
.B(n_1321),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1321),
.B(n_1279),
.Y(n_1461)
);

BUFx8_ASAP7_75t_L g1462 ( 
.A(n_1381),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1336),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1336),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1388),
.Y(n_1465)
);

INVx6_ASAP7_75t_L g1466 ( 
.A(n_1376),
.Y(n_1466)
);

BUFx8_ASAP7_75t_L g1467 ( 
.A(n_1376),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1380),
.A2(n_1267),
.B1(n_1289),
.B2(n_1328),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1376),
.Y(n_1469)
);

BUFx4f_ASAP7_75t_SL g1470 ( 
.A(n_1390),
.Y(n_1470)
);

AOI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1284),
.A2(n_1309),
.B(n_1286),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1367),
.A2(n_1373),
.B1(n_1267),
.B2(n_1380),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1397),
.B(n_1352),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1408),
.A2(n_1384),
.B1(n_1270),
.B2(n_1306),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1389),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1343),
.B(n_1337),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1408),
.A2(n_1384),
.B1(n_1270),
.B2(n_1337),
.Y(n_1477)
);

BUFx8_ASAP7_75t_SL g1478 ( 
.A(n_1390),
.Y(n_1478)
);

NAND2x1p5_ASAP7_75t_L g1479 ( 
.A(n_1394),
.B(n_1391),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1401),
.B(n_1347),
.Y(n_1480)
);

INVx6_ASAP7_75t_L g1481 ( 
.A(n_1390),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1288),
.A2(n_1334),
.B1(n_1342),
.B2(n_1407),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1285),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1391),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1383),
.Y(n_1485)
);

BUFx8_ASAP7_75t_SL g1486 ( 
.A(n_1318),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1419),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1355),
.Y(n_1488)
);

BUFx2_ASAP7_75t_SL g1489 ( 
.A(n_1387),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1318),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1344),
.A2(n_1316),
.B1(n_1310),
.B2(n_1301),
.Y(n_1491)
);

CKINVDCx11_ASAP7_75t_R g1492 ( 
.A(n_1318),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1407),
.A2(n_1401),
.B1(n_1333),
.B2(n_1386),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1293),
.A2(n_1361),
.B1(n_1287),
.B2(n_1332),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1377),
.A2(n_1330),
.B1(n_1385),
.B2(n_1281),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1355),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1319),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1331),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1355),
.Y(n_1499)
);

CKINVDCx11_ASAP7_75t_R g1500 ( 
.A(n_1412),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1330),
.A2(n_1281),
.B1(n_1324),
.B2(n_1371),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1272),
.A2(n_1294),
.B1(n_1269),
.B2(n_1295),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1307),
.A2(n_1420),
.B1(n_1409),
.B2(n_1399),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1368),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1398),
.A2(n_1300),
.B1(n_1303),
.B2(n_1382),
.Y(n_1505)
);

BUFx8_ASAP7_75t_L g1506 ( 
.A(n_1368),
.Y(n_1506)
);

CKINVDCx11_ASAP7_75t_R g1507 ( 
.A(n_1368),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_SL g1508 ( 
.A1(n_1278),
.A2(n_1374),
.B(n_1351),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1356),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1358),
.A2(n_1273),
.B1(n_1268),
.B2(n_1278),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1378),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1266),
.A2(n_1302),
.B1(n_1308),
.B2(n_1305),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1278),
.A2(n_1304),
.B1(n_1393),
.B2(n_1406),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1265),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1419),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1374),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1374),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1419),
.B(n_1357),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1357),
.A2(n_1418),
.B1(n_924),
.B2(n_1395),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1357),
.A2(n_924),
.B(n_1418),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1265),
.A2(n_1418),
.B1(n_924),
.B2(n_1417),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1265),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1418),
.A2(n_924),
.B(n_1414),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1524)
);

INVx6_ASAP7_75t_L g1525 ( 
.A(n_1297),
.Y(n_1525)
);

BUFx12f_ASAP7_75t_L g1526 ( 
.A(n_1274),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1417),
.B2(n_1414),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1395),
.A2(n_924),
.B1(n_1141),
.B2(n_831),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1283),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1417),
.B2(n_1414),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1283),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1392),
.B2(n_1396),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1325),
.A2(n_924),
.B1(n_1311),
.B2(n_1395),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1297),
.Y(n_1535)
);

CKINVDCx11_ASAP7_75t_R g1536 ( 
.A(n_1283),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1327),
.A2(n_1403),
.B1(n_1421),
.B2(n_1400),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1283),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1335),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1339),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1282),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1392),
.B2(n_1396),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_SL g1545 ( 
.A1(n_1395),
.A2(n_924),
.B1(n_1141),
.B2(n_831),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1282),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1282),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1417),
.B2(n_1414),
.Y(n_1550)
);

BUFx2_ASAP7_75t_R g1551 ( 
.A(n_1274),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1335),
.Y(n_1552)
);

CKINVDCx11_ASAP7_75t_R g1553 ( 
.A(n_1283),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1335),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1297),
.Y(n_1556)
);

INVx6_ASAP7_75t_SL g1557 ( 
.A(n_1267),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1395),
.A2(n_924),
.B1(n_1141),
.B2(n_831),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1335),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1392),
.B2(n_1396),
.Y(n_1560)
);

CKINVDCx11_ASAP7_75t_R g1561 ( 
.A(n_1283),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1395),
.A2(n_924),
.B1(n_1141),
.B2(n_831),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1339),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1418),
.A2(n_924),
.B1(n_1395),
.B2(n_1392),
.Y(n_1567)
);

BUFx8_ASAP7_75t_L g1568 ( 
.A(n_1297),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1274),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1297),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1282),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1483),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1532),
.A2(n_1543),
.B1(n_1560),
.B2(n_1428),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1508),
.A2(n_1495),
.B(n_1477),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1435),
.B(n_1438),
.Y(n_1575)
);

NAND2x1p5_ASAP7_75t_L g1576 ( 
.A(n_1498),
.B(n_1509),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1465),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1462),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1494),
.B(n_1520),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1528),
.A2(n_1562),
.B1(n_1558),
.B2(n_1545),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1495),
.A2(n_1477),
.B(n_1501),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1435),
.B(n_1438),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1488),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1485),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1511),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1496),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1522),
.B(n_1518),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1462),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1499),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1514),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1490),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1498),
.B(n_1509),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1445),
.A2(n_1550),
.B1(n_1527),
.B2(n_1530),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1523),
.A2(n_1533),
.B(n_1524),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_L g1595 ( 
.A(n_1524),
.B(n_1539),
.C(n_1533),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1519),
.B(n_1476),
.Y(n_1596)
);

AOI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1505),
.A2(n_1521),
.B(n_1503),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1487),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1515),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1475),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1515),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1519),
.B(n_1453),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1453),
.B(n_1507),
.Y(n_1603)
);

CKINVDCx6p67_ASAP7_75t_R g1604 ( 
.A(n_1434),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1516),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1490),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1449),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1517),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1504),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1504),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1451),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1451),
.B(n_1433),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1431),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1449),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1490),
.B(n_1427),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1571),
.Y(n_1616)
);

O2A1O1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1426),
.A2(n_1537),
.B(n_1544),
.C(n_1546),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1440),
.A2(n_1563),
.B1(n_1567),
.B2(n_1546),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1436),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1448),
.B(n_1539),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1448),
.B(n_1544),
.Y(n_1621)
);

OR2x6_ASAP7_75t_L g1622 ( 
.A(n_1472),
.B(n_1489),
.Y(n_1622)
);

CKINVDCx9p33_ASAP7_75t_R g1623 ( 
.A(n_1429),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1549),
.B(n_1555),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1529),
.B(n_1538),
.Y(n_1625)
);

INVx6_ASAP7_75t_L g1626 ( 
.A(n_1568),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1452),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1542),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1549),
.B(n_1555),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1547),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1563),
.B(n_1565),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1548),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1506),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1537),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1534),
.A2(n_1473),
.B1(n_1480),
.B2(n_1506),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1467),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1444),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1468),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1468),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1512),
.A2(n_1474),
.B(n_1501),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1502),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1565),
.B(n_1566),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1566),
.B(n_1567),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1502),
.Y(n_1644)
);

CKINVDCx16_ASAP7_75t_R g1645 ( 
.A(n_1437),
.Y(n_1645)
);

AOI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1491),
.A2(n_1430),
.B(n_1439),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1461),
.Y(n_1647)
);

BUFx2_ASAP7_75t_L g1648 ( 
.A(n_1557),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1474),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1557),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1442),
.A2(n_1443),
.B1(n_1455),
.B2(n_1459),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1500),
.Y(n_1652)
);

AOI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1442),
.A2(n_1497),
.B(n_1456),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1461),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1510),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1473),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1479),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1479),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1531),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1467),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1443),
.B(n_1458),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1513),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1456),
.B(n_1457),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1493),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1471),
.A2(n_1512),
.B(n_1482),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1460),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1460),
.A2(n_1541),
.B(n_1564),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1484),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1463),
.B(n_1464),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1525),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1452),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1469),
.A2(n_1570),
.B(n_1556),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1535),
.Y(n_1673)
);

AO21x1_ASAP7_75t_SL g1674 ( 
.A1(n_1557),
.A2(n_1492),
.B(n_1486),
.Y(n_1674)
);

OA21x2_ASAP7_75t_L g1675 ( 
.A1(n_1466),
.A2(n_1481),
.B(n_1470),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1525),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1525),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1470),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1579),
.A2(n_1622),
.B(n_1617),
.Y(n_1679)
);

AOI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1653),
.A2(n_1573),
.B(n_1651),
.C(n_1595),
.Y(n_1680)
);

INVx6_ASAP7_75t_L g1681 ( 
.A(n_1645),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1596),
.B(n_1536),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1596),
.B(n_1561),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1591),
.B(n_1425),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1659),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1637),
.B(n_1553),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1633),
.B(n_1551),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1591),
.B(n_1552),
.Y(n_1688)
);

O2A1O1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1594),
.A2(n_1540),
.B(n_1568),
.C(n_1447),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1633),
.B(n_1441),
.Y(n_1690)
);

OA21x2_ASAP7_75t_L g1691 ( 
.A1(n_1640),
.A2(n_1454),
.B(n_1559),
.Y(n_1691)
);

NOR2x1_ASAP7_75t_SL g1692 ( 
.A(n_1622),
.B(n_1446),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1585),
.B(n_1554),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1580),
.A2(n_1593),
.B(n_1618),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1585),
.B(n_1569),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1603),
.B(n_1432),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1579),
.B(n_1526),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1595),
.A2(n_1450),
.B(n_1478),
.C(n_1620),
.Y(n_1698)
);

OA21x2_ASAP7_75t_L g1699 ( 
.A1(n_1640),
.A2(n_1597),
.B(n_1638),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1663),
.B(n_1661),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1634),
.B(n_1450),
.Y(n_1701)
);

AO32x2_ASAP7_75t_L g1702 ( 
.A1(n_1607),
.A2(n_1614),
.A3(n_1610),
.B1(n_1609),
.B2(n_1676),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1635),
.A2(n_1629),
.B1(n_1642),
.B2(n_1584),
.Y(n_1703)
);

BUFx4f_ASAP7_75t_L g1704 ( 
.A(n_1626),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1600),
.B(n_1612),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_SL g1706 ( 
.A1(n_1622),
.A2(n_1675),
.B(n_1588),
.Y(n_1706)
);

NAND4xp25_ASAP7_75t_L g1707 ( 
.A(n_1638),
.B(n_1639),
.C(n_1643),
.D(n_1631),
.Y(n_1707)
);

AOI211xp5_ASAP7_75t_L g1708 ( 
.A1(n_1620),
.A2(n_1621),
.B(n_1652),
.C(n_1643),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_SL g1709 ( 
.A(n_1622),
.B(n_1579),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_SL g1710 ( 
.A(n_1622),
.B(n_1579),
.Y(n_1710)
);

NAND4xp25_ASAP7_75t_L g1711 ( 
.A(n_1639),
.B(n_1631),
.C(n_1624),
.D(n_1621),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1628),
.B(n_1632),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1624),
.A2(n_1582),
.B1(n_1575),
.B2(n_1602),
.C(n_1641),
.Y(n_1713)
);

OAI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1646),
.A2(n_1582),
.B(n_1575),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1598),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1626),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1602),
.A2(n_1644),
.B1(n_1611),
.B2(n_1664),
.C(n_1649),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1645),
.A2(n_1652),
.B1(n_1664),
.B2(n_1626),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1656),
.B(n_1646),
.Y(n_1719)
);

OAI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1625),
.A2(n_1579),
.B1(n_1611),
.B2(n_1614),
.C(n_1607),
.Y(n_1720)
);

OR2x6_ASAP7_75t_L g1721 ( 
.A(n_1576),
.B(n_1592),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1648),
.A2(n_1650),
.B1(n_1626),
.B2(n_1666),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1666),
.B(n_1677),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1669),
.B(n_1668),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1587),
.B(n_1608),
.Y(n_1725)
);

CKINVDCx20_ASAP7_75t_R g1726 ( 
.A(n_1623),
.Y(n_1726)
);

AOI21xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1578),
.A2(n_1588),
.B(n_1636),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1677),
.B(n_1655),
.Y(n_1728)
);

OA21x2_ASAP7_75t_L g1729 ( 
.A1(n_1583),
.A2(n_1589),
.B(n_1586),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1587),
.B(n_1608),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1613),
.B(n_1609),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_1604),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1669),
.B(n_1668),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1613),
.Y(n_1734)
);

AO32x2_ASAP7_75t_L g1735 ( 
.A1(n_1610),
.A2(n_1670),
.A3(n_1676),
.B1(n_1574),
.B2(n_1605),
.Y(n_1735)
);

A2O1A1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1649),
.A2(n_1655),
.B(n_1662),
.C(n_1660),
.Y(n_1736)
);

AND2x2_ASAP7_75t_SL g1737 ( 
.A(n_1581),
.B(n_1574),
.Y(n_1737)
);

NOR2xp67_ASAP7_75t_L g1738 ( 
.A(n_1578),
.B(n_1647),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1660),
.Y(n_1739)
);

AO32x2_ASAP7_75t_L g1740 ( 
.A1(n_1670),
.A2(n_1574),
.A3(n_1605),
.B1(n_1581),
.B2(n_1601),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1630),
.B(n_1616),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1665),
.A2(n_1581),
.B(n_1574),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1662),
.A2(n_1660),
.B(n_1667),
.C(n_1581),
.Y(n_1743)
);

O2A1O1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1665),
.A2(n_1673),
.B(n_1678),
.C(n_1672),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1700),
.A2(n_1665),
.B1(n_1648),
.B2(n_1650),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1729),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1681),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1700),
.A2(n_1703),
.B1(n_1697),
.B2(n_1711),
.Y(n_1748)
);

NAND3xp33_ASAP7_75t_L g1749 ( 
.A(n_1680),
.B(n_1654),
.C(n_1657),
.Y(n_1749)
);

OAI22xp33_ASAP7_75t_SL g1750 ( 
.A1(n_1697),
.A2(n_1671),
.B1(n_1619),
.B2(n_1616),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1725),
.B(n_1599),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1697),
.A2(n_1654),
.B1(n_1647),
.B2(n_1592),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1693),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1729),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1715),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1730),
.B(n_1599),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_SL g1757 ( 
.A1(n_1679),
.A2(n_1675),
.B1(n_1647),
.B2(n_1606),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1737),
.B(n_1724),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1726),
.Y(n_1759)
);

BUFx2_ASAP7_75t_SL g1760 ( 
.A(n_1726),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1721),
.B(n_1592),
.Y(n_1761)
);

BUFx4f_ASAP7_75t_SL g1762 ( 
.A(n_1684),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1737),
.B(n_1590),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1721),
.B(n_1592),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1721),
.B(n_1577),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1733),
.B(n_1590),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_SL g1767 ( 
.A1(n_1679),
.A2(n_1675),
.B1(n_1647),
.B2(n_1606),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1694),
.B(n_1657),
.C(n_1658),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1731),
.B(n_1601),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1705),
.B(n_1572),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1699),
.B(n_1572),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1686),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1708),
.B(n_1627),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1699),
.B(n_1572),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1713),
.A2(n_1615),
.B1(n_1674),
.B2(n_1658),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1713),
.A2(n_1615),
.B1(n_1674),
.B2(n_1671),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1741),
.Y(n_1777)
);

INVxp67_ASAP7_75t_L g1778 ( 
.A(n_1723),
.Y(n_1778)
);

INVxp33_ASAP7_75t_SL g1779 ( 
.A(n_1732),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1684),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1685),
.B(n_1667),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1712),
.Y(n_1782)
);

NOR2xp67_ASAP7_75t_L g1783 ( 
.A(n_1746),
.B(n_1742),
.Y(n_1783)
);

NOR2x1_ASAP7_75t_L g1784 ( 
.A(n_1747),
.B(n_1706),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1761),
.B(n_1709),
.Y(n_1785)
);

AOI211xp5_ASAP7_75t_L g1786 ( 
.A1(n_1749),
.A2(n_1698),
.B(n_1744),
.C(n_1689),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1778),
.B(n_1714),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1754),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1755),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1782),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_L g1791 ( 
.A1(n_1746),
.A2(n_1742),
.B(n_1744),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1758),
.B(n_1735),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1758),
.B(n_1735),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1763),
.B(n_1735),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1755),
.Y(n_1795)
);

AOI221xp5_ASAP7_75t_L g1796 ( 
.A1(n_1748),
.A2(n_1717),
.B1(n_1707),
.B2(n_1736),
.C(n_1719),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1763),
.B(n_1735),
.Y(n_1797)
);

OR2x6_ASAP7_75t_SL g1798 ( 
.A(n_1768),
.B(n_1718),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1770),
.B(n_1743),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1751),
.B(n_1743),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1777),
.B(n_1728),
.Y(n_1801)
);

NOR2x1_ASAP7_75t_L g1802 ( 
.A(n_1747),
.B(n_1719),
.Y(n_1802)
);

INVx5_ASAP7_75t_L g1803 ( 
.A(n_1781),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1773),
.A2(n_1692),
.B(n_1710),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1761),
.B(n_1702),
.Y(n_1805)
);

AND2x2_ASAP7_75t_SL g1806 ( 
.A(n_1745),
.B(n_1691),
.Y(n_1806)
);

BUFx3_ASAP7_75t_L g1807 ( 
.A(n_1781),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1751),
.B(n_1734),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1761),
.B(n_1702),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1764),
.B(n_1740),
.Y(n_1810)
);

INVxp67_ASAP7_75t_L g1811 ( 
.A(n_1760),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1756),
.B(n_1691),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1769),
.B(n_1691),
.Y(n_1813)
);

BUFx2_ASAP7_75t_L g1814 ( 
.A(n_1781),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1764),
.B(n_1740),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1750),
.B(n_1716),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_SL g1817 ( 
.A1(n_1760),
.A2(n_1683),
.B1(n_1682),
.B2(n_1681),
.Y(n_1817)
);

OAI31xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1780),
.A2(n_1720),
.A3(n_1717),
.B(n_1696),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1810),
.B(n_1815),
.Y(n_1819)
);

NAND2xp33_ASAP7_75t_R g1820 ( 
.A(n_1798),
.B(n_1779),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1788),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1788),
.Y(n_1822)
);

AND2x4_ASAP7_75t_SL g1823 ( 
.A(n_1785),
.B(n_1764),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1792),
.B(n_1793),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1793),
.B(n_1794),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1803),
.B(n_1765),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1794),
.B(n_1757),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1797),
.B(n_1767),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1797),
.B(n_1805),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1789),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1813),
.B(n_1771),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1809),
.B(n_1766),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1809),
.B(n_1766),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1789),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1812),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1812),
.B(n_1771),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1814),
.B(n_1765),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1795),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1799),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1786),
.B(n_1818),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1803),
.B(n_1774),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1798),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1783),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1842),
.B(n_1787),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1830),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1840),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1821),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1830),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_SL g1849 ( 
.A(n_1842),
.B(n_1779),
.Y(n_1849)
);

OR2x6_ASAP7_75t_L g1850 ( 
.A(n_1840),
.B(n_1804),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1839),
.B(n_1829),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1821),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1839),
.B(n_1799),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1839),
.B(n_1796),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1823),
.B(n_1807),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1830),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1821),
.Y(n_1857)
);

NAND2x1_ASAP7_75t_L g1858 ( 
.A(n_1826),
.B(n_1804),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1834),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1821),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1823),
.B(n_1785),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1823),
.B(n_1785),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1822),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1822),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1823),
.B(n_1785),
.Y(n_1865)
);

INVxp67_ASAP7_75t_SL g1866 ( 
.A(n_1820),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1834),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1837),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1839),
.B(n_1790),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1829),
.B(n_1800),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1829),
.B(n_1800),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1834),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1827),
.B(n_1828),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1838),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1827),
.B(n_1803),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1822),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1838),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1827),
.B(n_1801),
.Y(n_1878)
);

INVxp67_ASAP7_75t_SL g1879 ( 
.A(n_1820),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1822),
.Y(n_1880)
);

INVxp67_ASAP7_75t_SL g1881 ( 
.A(n_1843),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1827),
.B(n_1802),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_L g1883 ( 
.A(n_1826),
.B(n_1784),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1826),
.B(n_1803),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1828),
.B(n_1802),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1838),
.Y(n_1886)
);

OAI21xp33_ASAP7_75t_L g1887 ( 
.A1(n_1828),
.A2(n_1806),
.B(n_1786),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1829),
.B(n_1808),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1828),
.B(n_1803),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_SL g1890 ( 
.A(n_1826),
.B(n_1784),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1870),
.B(n_1831),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1846),
.B(n_1832),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1875),
.B(n_1819),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1887),
.A2(n_1850),
.B1(n_1879),
.B2(n_1866),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1851),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1854),
.B(n_1844),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1870),
.B(n_1831),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1871),
.B(n_1831),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1849),
.B(n_1759),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1871),
.B(n_1836),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1851),
.B(n_1836),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1875),
.B(n_1819),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1845),
.Y(n_1903)
);

INVx1_ASAP7_75t_SL g1904 ( 
.A(n_1850),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1889),
.B(n_1819),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1889),
.B(n_1825),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1845),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1873),
.B(n_1836),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1883),
.B(n_1826),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1848),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1861),
.B(n_1825),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1850),
.A2(n_1817),
.B1(n_1811),
.B2(n_1806),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1861),
.B(n_1825),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1883),
.B(n_1826),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1848),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1878),
.B(n_1832),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1856),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1887),
.B(n_1832),
.Y(n_1918)
);

NAND2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1858),
.B(n_1816),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1856),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1881),
.B(n_1833),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1862),
.B(n_1865),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1859),
.Y(n_1923)
);

OR3x2_ASAP7_75t_L g1924 ( 
.A(n_1850),
.B(n_1678),
.C(n_1689),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1850),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1862),
.B(n_1825),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1865),
.B(n_1824),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1894),
.B(n_1882),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1893),
.B(n_1868),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1918),
.B(n_1853),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1924),
.A2(n_1890),
.B1(n_1885),
.B2(n_1806),
.Y(n_1931)
);

HB1xp67_ASAP7_75t_L g1932 ( 
.A(n_1906),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1912),
.A2(n_1884),
.B1(n_1853),
.B2(n_1868),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1893),
.B(n_1855),
.Y(n_1934)
);

OAI211xp5_ASAP7_75t_SL g1935 ( 
.A1(n_1896),
.A2(n_1869),
.B(n_1772),
.C(n_1698),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1903),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1906),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1907),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1902),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1925),
.B(n_1824),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1910),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1915),
.Y(n_1942)
);

INVxp67_ASAP7_75t_L g1943 ( 
.A(n_1899),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1904),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1919),
.A2(n_1858),
.B(n_1884),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1902),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1905),
.B(n_1884),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1905),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1892),
.B(n_1753),
.Y(n_1949)
);

OAI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1919),
.A2(n_1888),
.B1(n_1803),
.B2(n_1722),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1908),
.B(n_1727),
.Y(n_1951)
);

XNOR2xp5_ASAP7_75t_L g1952 ( 
.A(n_1924),
.B(n_1687),
.Y(n_1952)
);

INVxp67_ASAP7_75t_L g1953 ( 
.A(n_1921),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1927),
.B(n_1911),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1946),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1947),
.Y(n_1956)
);

AOI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1952),
.A2(n_1922),
.B1(n_1914),
.B2(n_1909),
.Y(n_1957)
);

AOI21xp5_ASAP7_75t_SL g1958 ( 
.A1(n_1952),
.A2(n_1914),
.B(n_1909),
.Y(n_1958)
);

AOI21xp33_ASAP7_75t_L g1959 ( 
.A1(n_1943),
.A2(n_1908),
.B(n_1895),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1934),
.B(n_1922),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1944),
.B(n_1927),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1940),
.B(n_1916),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1948),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1932),
.Y(n_1964)
);

OAI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1931),
.A2(n_1895),
.B1(n_1897),
.B2(n_1898),
.C(n_1891),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1928),
.B(n_1911),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1934),
.B(n_1929),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1947),
.Y(n_1968)
);

OAI21xp33_ASAP7_75t_L g1969 ( 
.A1(n_1933),
.A2(n_1926),
.B(n_1913),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1937),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1929),
.B(n_1913),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1953),
.B(n_1926),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1936),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1936),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1938),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1960),
.Y(n_1976)
);

AOI222xp33_ASAP7_75t_L g1977 ( 
.A1(n_1965),
.A2(n_1935),
.B1(n_1938),
.B2(n_1942),
.C1(n_1941),
.C2(n_1950),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1967),
.B(n_1947),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1957),
.A2(n_1954),
.B1(n_1939),
.B2(n_1930),
.Y(n_1979)
);

O2A1O1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1955),
.A2(n_1941),
.B(n_1942),
.C(n_1951),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1960),
.B(n_1945),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1961),
.B(n_1909),
.Y(n_1982)
);

OAI31xp33_ASAP7_75t_L g1983 ( 
.A1(n_1969),
.A2(n_1930),
.A3(n_1914),
.B(n_1939),
.Y(n_1983)
);

O2A1O1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1963),
.A2(n_1923),
.B(n_1920),
.C(n_1917),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1966),
.B(n_1891),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1958),
.A2(n_1949),
.B(n_1884),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1967),
.B(n_1897),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1964),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1976),
.B(n_1968),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1978),
.B(n_1956),
.Y(n_1990)
);

NOR2x1_ASAP7_75t_L g1991 ( 
.A(n_1981),
.B(n_1958),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1987),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1988),
.B(n_1959),
.Y(n_1993)
);

NAND4xp25_ASAP7_75t_L g1994 ( 
.A(n_1977),
.B(n_1970),
.C(n_1972),
.D(n_1956),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1977),
.B(n_1971),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1983),
.B(n_1971),
.Y(n_1996)
);

BUFx3_ASAP7_75t_L g1997 ( 
.A(n_1985),
.Y(n_1997)
);

NAND2xp33_ASAP7_75t_SL g1998 ( 
.A(n_1982),
.B(n_1962),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_SL g1999 ( 
.A(n_1986),
.B(n_1973),
.Y(n_1999)
);

NAND3xp33_ASAP7_75t_L g2000 ( 
.A(n_1980),
.B(n_1974),
.C(n_1975),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1984),
.Y(n_2001)
);

NAND3xp33_ASAP7_75t_L g2002 ( 
.A(n_1999),
.B(n_1979),
.C(n_1975),
.Y(n_2002)
);

OAI221xp5_ASAP7_75t_L g2003 ( 
.A1(n_1991),
.A2(n_1962),
.B1(n_1900),
.B2(n_1898),
.C(n_1901),
.Y(n_2003)
);

OAI321xp33_ASAP7_75t_L g2004 ( 
.A1(n_1995),
.A2(n_1900),
.A3(n_1901),
.B1(n_1855),
.B2(n_1636),
.C(n_1776),
.Y(n_2004)
);

NAND4xp25_ASAP7_75t_SL g2005 ( 
.A(n_1996),
.B(n_1695),
.C(n_1888),
.D(n_1690),
.Y(n_2005)
);

OAI221xp5_ASAP7_75t_L g2006 ( 
.A1(n_1994),
.A2(n_1843),
.B1(n_1681),
.B2(n_1835),
.C(n_1739),
.Y(n_2006)
);

OAI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1994),
.A2(n_1835),
.B1(n_1886),
.B2(n_1877),
.C(n_1859),
.Y(n_2007)
);

OAI211xp5_ASAP7_75t_SL g2008 ( 
.A1(n_1993),
.A2(n_1852),
.B(n_1880),
.C(n_1860),
.Y(n_2008)
);

AOI221x1_ASAP7_75t_L g2009 ( 
.A1(n_2000),
.A2(n_1886),
.B1(n_1867),
.B2(n_1877),
.C(n_1872),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_2002),
.A2(n_2001),
.B1(n_1997),
.B2(n_1992),
.Y(n_2010)
);

AOI211xp5_ASAP7_75t_L g2011 ( 
.A1(n_2003),
.A2(n_1990),
.B(n_1989),
.C(n_1998),
.Y(n_2011)
);

NAND5xp2_ASAP7_75t_L g2012 ( 
.A(n_2004),
.B(n_1775),
.C(n_1701),
.D(n_1752),
.E(n_1736),
.Y(n_2012)
);

XNOR2x1_ASAP7_75t_SL g2013 ( 
.A(n_2005),
.B(n_1837),
.Y(n_2013)
);

A2O1A1Ixp33_ASAP7_75t_L g2014 ( 
.A1(n_2006),
.A2(n_1791),
.B(n_1704),
.C(n_1841),
.Y(n_2014)
);

AOI211xp5_ASAP7_75t_SL g2015 ( 
.A1(n_2007),
.A2(n_1762),
.B(n_1738),
.C(n_1872),
.Y(n_2015)
);

NOR3xp33_ASAP7_75t_L g2016 ( 
.A(n_2008),
.B(n_1688),
.C(n_1852),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_2009),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2010),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_2017),
.B(n_1867),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2013),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_2015),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2011),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_2016),
.B(n_1824),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2020),
.Y(n_2024)
);

OAI221xp5_ASAP7_75t_L g2025 ( 
.A1(n_2022),
.A2(n_2014),
.B1(n_2012),
.B2(n_1880),
.C(n_1876),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_2018),
.Y(n_2026)
);

OAI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_2024),
.A2(n_2021),
.B1(n_2023),
.B2(n_2019),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2027),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2028),
.Y(n_2029)
);

INVx3_ASAP7_75t_SL g2030 ( 
.A(n_2028),
.Y(n_2030)
);

OAI22x1_ASAP7_75t_L g2031 ( 
.A1(n_2030),
.A2(n_2026),
.B1(n_2021),
.B2(n_2019),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_SL g2032 ( 
.A1(n_2029),
.A2(n_2025),
.B1(n_1688),
.B2(n_1876),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2031),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_2032),
.A2(n_1880),
.B1(n_1876),
.B2(n_1852),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_2033),
.A2(n_1860),
.B1(n_1864),
.B2(n_1863),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_2034),
.A2(n_1860),
.B(n_1857),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_2035),
.A2(n_1864),
.B1(n_1863),
.B2(n_1857),
.Y(n_2037)
);

CKINVDCx20_ASAP7_75t_R g2038 ( 
.A(n_2037),
.Y(n_2038)
);

OAI221xp5_ASAP7_75t_R g2039 ( 
.A1(n_2038),
.A2(n_2036),
.B1(n_1847),
.B2(n_1874),
.C(n_1835),
.Y(n_2039)
);

AOI211xp5_ASAP7_75t_L g2040 ( 
.A1(n_2039),
.A2(n_1847),
.B(n_1874),
.C(n_1835),
.Y(n_2040)
);


endmodule