module fake_netlist_1_10825_n_42 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_42);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_42;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_30;
wire n_16;
wire n_26;
wire n_33;
wire n_25;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_8), .B(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_0), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_2), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_10), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_3), .Y(n_21) );
NAND2xp5_ASAP7_75t_SL g22 ( .A(n_14), .B(n_0), .Y(n_22) );
AND3x1_ASAP7_75t_L g23 ( .A(n_17), .B(n_1), .C(n_3), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
BUFx2_ASAP7_75t_R g25 ( .A(n_22), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_19), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_26), .B(n_21), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_26), .B(n_23), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
INVx1_ASAP7_75t_SL g30 ( .A(n_27), .Y(n_30) );
AOI221xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_18), .B1(n_17), .B2(n_19), .C(n_20), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
AOI211xp5_ASAP7_75t_SL g33 ( .A1(n_31), .A2(n_18), .B(n_15), .C(n_16), .Y(n_33) );
AOI21xp33_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_30), .B(n_15), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
NOR3x2_ASAP7_75t_L g36 ( .A(n_33), .B(n_25), .C(n_4), .Y(n_36) );
XNOR2x1_ASAP7_75t_L g37 ( .A(n_35), .B(n_1), .Y(n_37) );
NOR4xp75_ASAP7_75t_L g38 ( .A(n_34), .B(n_4), .C(n_15), .D(n_14), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_37), .B(n_35), .Y(n_39) );
OAI22xp5_ASAP7_75t_L g40 ( .A1(n_37), .A2(n_6), .B1(n_7), .B2(n_9), .Y(n_40) );
NAND2xp5_ASAP7_75t_L g41 ( .A(n_39), .B(n_36), .Y(n_41) );
AOI22x1_ASAP7_75t_L g42 ( .A1(n_41), .A2(n_38), .B1(n_40), .B2(n_12), .Y(n_42) );
endmodule