module fake_jpeg_10437_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_2),
.B(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_62),
.Y(n_80)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_67),
.Y(n_86)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_1),
.CON(n_64),
.SN(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_56),
.B(n_12),
.C(n_13),
.Y(n_82)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_40),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_4),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_28),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_74),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_48),
.B1(n_54),
.B2(n_51),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_50),
.B1(n_42),
.B2(n_57),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_40),
.B1(n_47),
.B2(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_77),
.B1(n_83),
.B2(n_84),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_87),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_85),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_11),
.B1(n_15),
.B2(n_16),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_39),
.B1(n_32),
.B2(n_34),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_98),
.B1(n_99),
.B2(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

AOI321xp33_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_103),
.A3(n_95),
.B1(n_97),
.B2(n_101),
.C(n_85),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_80),
.C(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_89),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_93),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_79),
.C(n_86),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_92),
.B(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_31),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_37),
.Y(n_116)
);


endmodule