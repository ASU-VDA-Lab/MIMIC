module fake_jpeg_28684_n_451 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_451);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_451;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_8),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_51),
.B(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_25),
.B(n_9),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_56),
.B(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_9),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_58),
.B(n_66),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_24),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_9),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_27),
.B(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_73),
.Y(n_126)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_6),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_81),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_28),
.B(n_6),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_30),
.B(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_87),
.Y(n_140)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_89),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_30),
.B(n_5),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_36),
.A2(n_5),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_47),
.B1(n_42),
.B2(n_40),
.Y(n_98)
);

BUFx2_ASAP7_75t_R g91 ( 
.A(n_29),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_97),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_98),
.A2(n_100),
.B1(n_118),
.B2(n_128),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_44),
.B1(n_21),
.B2(n_33),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_114),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_44),
.B1(n_46),
.B2(n_35),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_102),
.A2(n_122),
.B1(n_143),
.B2(n_38),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_58),
.A2(n_47),
.B1(n_42),
.B2(n_40),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_113),
.A2(n_135),
.B1(n_84),
.B2(n_61),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_51),
.B(n_39),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_55),
.A2(n_39),
.B1(n_19),
.B2(n_33),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_31),
.C(n_20),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_139),
.C(n_78),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_65),
.A2(n_46),
.B1(n_38),
.B2(n_35),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_31),
.B1(n_20),
.B2(n_21),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_32),
.B1(n_19),
.B2(n_35),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_11),
.B(n_2),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_72),
.A2(n_32),
.B1(n_46),
.B2(n_38),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_57),
.B(n_46),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_88),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_76),
.B(n_38),
.C(n_1),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_93),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_150),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_73),
.C(n_67),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_151),
.B(n_166),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_63),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_156),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_107),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_153),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_119),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_100),
.A2(n_87),
.B(n_88),
.C(n_85),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_170),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_85),
.B(n_60),
.C(n_66),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_159),
.A2(n_120),
.B(n_110),
.C(n_123),
.Y(n_235)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_48),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_161),
.B(n_171),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_59),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_167),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVx6_ASAP7_75t_SL g234 ( 
.A(n_168),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_50),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_169),
.B(n_130),
.Y(n_217)
);

OR2x4_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_92),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_86),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_179),
.B1(n_109),
.B2(n_145),
.Y(n_200)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_184),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_129),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_177),
.B(n_186),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_98),
.A2(n_79),
.B1(n_83),
.B2(n_71),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

INVx4_ASAP7_75t_SL g181 ( 
.A(n_121),
.Y(n_181)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_94),
.B(n_144),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_187),
.A2(n_62),
.B1(n_109),
.B2(n_131),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_112),
.A2(n_49),
.B1(n_64),
.B2(n_61),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_190),
.B(n_105),
.Y(n_218)
);

CKINVDCx12_ASAP7_75t_R g191 ( 
.A(n_137),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_141),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_120),
.Y(n_219)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_84),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_123),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_149),
.A2(n_121),
.B1(n_130),
.B2(n_103),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_200),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_170),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_202),
.B(n_209),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_181),
.B1(n_153),
.B2(n_167),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_178),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_230),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_218),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_165),
.Y(n_249)
);

AO22x2_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_131),
.B1(n_106),
.B2(n_111),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_220),
.B(n_235),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_149),
.A2(n_95),
.B1(n_115),
.B2(n_134),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_226),
.A2(n_236),
.B1(n_181),
.B2(n_167),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_134),
.Y(n_228)
);

NOR2x1_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_166),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_169),
.A2(n_95),
.B1(n_111),
.B2(n_110),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_148),
.B(n_0),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_166),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_151),
.C(n_152),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_265),
.C(n_206),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_239),
.A2(n_250),
.B1(n_207),
.B2(n_225),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_189),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_240),
.B(n_243),
.Y(n_277)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_242),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_201),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_200),
.B1(n_236),
.B2(n_208),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_177),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_246),
.B(n_247),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_195),
.B(n_168),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_255),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_253),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_196),
.B1(n_206),
.B2(n_230),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_195),
.B(n_157),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_203),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_222),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_150),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_262),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_257),
.Y(n_279)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_204),
.B(n_147),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_204),
.B(n_173),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_272),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_208),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_233),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_159),
.C(n_190),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_172),
.B(n_158),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_266),
.A2(n_270),
.B(n_273),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_214),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_269),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_186),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_224),
.A2(n_183),
.B1(n_174),
.B2(n_175),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_271),
.A2(n_233),
.B1(n_227),
.B2(n_203),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_182),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_185),
.B(n_154),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_180),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_220),
.B(n_160),
.Y(n_275)
);

AOI221xp5_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_202),
.B1(n_232),
.B2(n_235),
.C(n_217),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_L g328 ( 
.A1(n_276),
.A2(n_278),
.B(n_242),
.C(n_259),
.D(n_261),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_220),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_303),
.C(n_265),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_281),
.A2(n_310),
.B1(n_244),
.B2(n_274),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_247),
.A2(n_234),
.B1(n_225),
.B2(n_216),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_282),
.A2(n_298),
.B(n_267),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_223),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_269),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_284),
.A2(n_291),
.B1(n_300),
.B2(n_239),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_242),
.Y(n_326)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_252),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_299),
.Y(n_327)
);

AOI32xp33_ASAP7_75t_L g298 ( 
.A1(n_260),
.A2(n_266),
.A3(n_263),
.B1(n_262),
.B2(n_250),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_260),
.A2(n_199),
.B1(n_227),
.B2(n_234),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_199),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_304),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_215),
.C(n_216),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_215),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_273),
.A2(n_231),
.B(n_153),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_297),
.B(n_310),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_267),
.A2(n_155),
.B1(n_176),
.B2(n_205),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_311),
.A2(n_317),
.B1(n_336),
.B2(n_284),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_314),
.C(n_315),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_270),
.C(n_254),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_270),
.C(n_272),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_275),
.C(n_264),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_322),
.C(n_297),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_301),
.A2(n_267),
.B1(n_259),
.B2(n_271),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_318),
.A2(n_324),
.B(n_330),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_277),
.B(n_308),
.Y(n_320)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_321),
.A2(n_283),
.B1(n_290),
.B2(n_307),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_243),
.C(n_240),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_309),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_323),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_325),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_326),
.B(n_337),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_329),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_304),
.B(n_258),
.Y(n_331)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_331),
.Y(n_346)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_251),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_333),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_251),
.Y(n_334)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_334),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_287),
.B(n_257),
.Y(n_335)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_335),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_281),
.A2(n_294),
.B1(n_306),
.B2(n_285),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_293),
.B(n_255),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_288),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_338),
.A2(n_295),
.B1(n_292),
.B2(n_288),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_305),
.A2(n_255),
.B(n_231),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_339),
.A2(n_290),
.B(n_292),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_342),
.B(n_365),
.Y(n_369)
);

FAx1_ASAP7_75t_SL g386 ( 
.A(n_344),
.B(n_213),
.CI(n_146),
.CON(n_386),
.SN(n_386)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_347),
.A2(n_351),
.B1(n_361),
.B2(n_334),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_338),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_289),
.C(n_293),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_352),
.C(n_353),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_311),
.A2(n_336),
.B1(n_317),
.B2(n_318),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_315),
.C(n_316),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_294),
.C(n_306),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_300),
.C(n_296),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_324),
.C(n_327),
.Y(n_375)
);

AO22x1_ASAP7_75t_L g379 ( 
.A1(n_359),
.A2(n_333),
.B1(n_332),
.B2(n_329),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_360),
.A2(n_362),
.B1(n_164),
.B2(n_210),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_339),
.A2(n_291),
.B1(n_279),
.B2(n_309),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_321),
.A2(n_279),
.B1(n_309),
.B2(n_163),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_312),
.B(n_178),
.Y(n_365)
);

INVx13_ASAP7_75t_L g366 ( 
.A(n_363),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_366),
.B(n_370),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_367),
.A2(n_379),
.B1(n_362),
.B2(n_358),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_358),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_368),
.Y(n_387)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_371),
.B(n_374),
.Y(n_390)
);

AOI322xp5_ASAP7_75t_SL g372 ( 
.A1(n_343),
.A2(n_320),
.A3(n_328),
.B1(n_344),
.B2(n_360),
.C1(n_356),
.C2(n_353),
.Y(n_372)
);

BUFx24_ASAP7_75t_SL g400 ( 
.A(n_372),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_331),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_386),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_327),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_376),
.B(n_380),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_342),
.B(n_312),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_382),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_337),
.C(n_319),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_357),
.C(n_348),
.Y(n_394)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_341),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_364),
.B(n_319),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_381),
.A2(n_384),
.B1(n_385),
.B2(n_361),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_178),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_347),
.A2(n_323),
.B1(n_163),
.B2(n_210),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_383),
.A2(n_355),
.B1(n_345),
.B2(n_354),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_213),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_401),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_340),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_399),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_394),
.B(n_396),
.Y(n_413)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_395),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_375),
.A2(n_356),
.B(n_345),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_378),
.C(n_377),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_398),
.C(n_403),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_365),
.C(n_348),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_351),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_382),
.B(n_359),
.C(n_354),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_408),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_367),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_412),
.Y(n_421)
);

BUFx4f_ASAP7_75t_SL g408 ( 
.A(n_402),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_394),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_409),
.B(n_416),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_400),
.B(n_374),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_414),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_386),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_397),
.B(n_368),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_388),
.B(n_368),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_406),
.A2(n_383),
.B1(n_392),
.B2(n_388),
.Y(n_420)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_420),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_407),
.A2(n_390),
.B1(n_379),
.B2(n_391),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_424),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_405),
.A2(n_385),
.B1(n_379),
.B2(n_370),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_425),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_412),
.A2(n_386),
.B1(n_398),
.B2(n_380),
.Y(n_424)
);

INVx11_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_366),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_426),
.B(n_427),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_410),
.B(n_393),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_371),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_428),
.A2(n_221),
.B(n_205),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_421),
.A2(n_413),
.B(n_415),
.Y(n_429)
);

OAI221xp5_ASAP7_75t_L g440 ( 
.A1(n_429),
.A2(n_431),
.B1(n_436),
.B2(n_5),
.C(n_11),
.Y(n_440)
);

OAI21xp33_ASAP7_75t_L g431 ( 
.A1(n_417),
.A2(n_389),
.B(n_415),
.Y(n_431)
);

AOI322xp5_ASAP7_75t_L g438 ( 
.A1(n_431),
.A2(n_424),
.A3(n_428),
.B1(n_422),
.B2(n_420),
.C1(n_193),
.C2(n_14),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_418),
.C(n_428),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_434),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_425),
.B(n_221),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_3),
.Y(n_442)
);

A2O1A1Ixp33_ASAP7_75t_SL g445 ( 
.A1(n_438),
.A2(n_440),
.B(n_11),
.C(n_12),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_437),
.A2(n_430),
.B1(n_436),
.B2(n_432),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_439),
.B(n_442),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_429),
.B(n_11),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_443),
.B(n_15),
.Y(n_447)
);

MAJx2_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_446),
.C(n_0),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_438),
.C(n_14),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_447),
.A2(n_0),
.B(n_444),
.Y(n_448)
);

AOI21xp33_ASAP7_75t_L g450 ( 
.A1(n_448),
.A2(n_449),
.B(n_0),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_0),
.Y(n_451)
);


endmodule