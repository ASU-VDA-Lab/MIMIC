module real_jpeg_30012_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_0),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_0),
.A2(n_27),
.B1(n_48),
.B2(n_50),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_0),
.A2(n_27),
.B1(n_54),
.B2(n_55),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_1),
.B(n_48),
.Y(n_86)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_2),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_101),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_2),
.A2(n_48),
.B1(n_50),
.B2(n_101),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_101),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_3),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_3),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_145)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_6),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_6),
.A2(n_29),
.B(n_33),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_114),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_6),
.B(n_31),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_6),
.A2(n_54),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_6),
.B(n_54),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_6),
.B(n_68),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_6),
.A2(n_85),
.B1(n_240),
.B2(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_6),
.A2(n_32),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_7),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_99),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_99),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_7),
.A2(n_48),
.B1(n_50),
.B2(n_99),
.Y(n_234)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_9),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_9),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_10),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_104),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_104),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_10),
.A2(n_48),
.B1(n_50),
.B2(n_104),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_11),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_94),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_94),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_12),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_12),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_12),
.A2(n_50),
.A3(n_54),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_13),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_13),
.A2(n_36),
.B1(n_48),
.B2(n_50),
.Y(n_126)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_17),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_110),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_17),
.A2(n_54),
.B1(n_55),
.B2(n_110),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_17),
.A2(n_48),
.B1(n_50),
.B2(n_110),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_331),
.B(n_334),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_76),
.B(n_330),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_21),
.B(n_37),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_21),
.B(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_21),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_23),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_25),
.A2(n_34),
.B(n_114),
.C(n_115),
.Y(n_113)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_28),
.A2(n_31),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_28),
.A2(n_31),
.B1(n_100),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_28),
.A2(n_31),
.B1(n_109),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_28),
.A2(n_31),
.B(n_35),
.Y(n_333)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_31),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_60),
.Y(n_62)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_32),
.A2(n_55),
.A3(n_64),
.B1(n_257),
.B2(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_33),
.B(n_114),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_69),
.C(n_71),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_38),
.A2(n_39),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_57),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_40),
.B(n_314),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_42),
.A2(n_73),
.B1(n_75),
.B2(n_164),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_46),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_46),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_46),
.A2(n_57),
.B1(n_308),
.B2(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_52),
.B(n_56),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_47),
.A2(n_52),
.B1(n_92),
.B2(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_47),
.A2(n_52),
.B1(n_95),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_47),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_47),
.A2(n_52),
.B1(n_56),
.B2(n_137),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_47),
.A2(n_52),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_47),
.A2(n_52),
.B1(n_215),
.B2(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_47),
.B(n_114),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_47),
.A2(n_52),
.B1(n_182),
.B2(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_48),
.B(n_51),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_48),
.B(n_246),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_52),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_54),
.B(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_57),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_68),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_58),
.A2(n_68),
.B1(n_105),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_58),
.A2(n_68),
.B1(n_178),
.B2(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_58),
.A2(n_66),
.B1(n_68),
.B2(n_306),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_63),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_63),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_59),
.A2(n_63),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_59),
.A2(n_63),
.B1(n_122),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_59),
.A2(n_63),
.B1(n_190),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_64),
.Y(n_266)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_69),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_75),
.B1(n_108),
.B2(n_111),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_73),
.A2(n_75),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_323),
.B(n_329),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_299),
.A3(n_318),
.B1(n_321),
.B2(n_322),
.C(n_340),
.Y(n_77)
);

AOI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_148),
.A3(n_170),
.B1(n_293),
.B2(n_298),
.C(n_341),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_80),
.A2(n_294),
.B(n_297),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_129),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_81),
.B(n_129),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_106),
.C(n_124),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_82),
.B(n_124),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_96),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_97),
.C(n_102),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_84),
.B(n_91),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_90),
.B1(n_119),
.B2(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_85),
.A2(n_119),
.B(n_126),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_85),
.A2(n_89),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_85),
.A2(n_89),
.B1(n_234),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_85),
.A2(n_229),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_88),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_86),
.A2(n_117),
.B1(n_120),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_86),
.A2(n_120),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_89),
.B(n_114),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_93),
.A2(n_135),
.B1(n_138),
.B2(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_106),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.C(n_121),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_107),
.B(n_121),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_112),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_113),
.B(n_116),
.Y(n_185)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_SL g268 ( 
.A(n_120),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_127),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_128),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_147),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_141),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_141),
.C(n_147),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_139),
.B2(n_140),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_132),
.B(n_140),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_138),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_135),
.A2(n_138),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_140),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_139),
.A2(n_162),
.B(n_165),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_141),
.Y(n_338)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_144),
.CI(n_146),
.CON(n_141),
.SN(n_141)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_144),
.C(n_146),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_143),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_149),
.B(n_150),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_168),
.B2(n_169),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_153),
.B(n_159),
.C(n_169),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_157),
.B(n_158),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_157),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_156),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_158),
.B(n_301),
.C(n_310),
.Y(n_300)
);

FAx1_ASAP7_75t_L g320 ( 
.A(n_158),
.B(n_301),
.CI(n_310),
.CON(n_320),
.SN(n_320)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_168),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_200),
.C(n_205),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_194),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_172),
.B(n_194),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_185),
.C(n_186),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_173),
.B(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_183),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_180),
.C(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_185),
.Y(n_291)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_188),
.B(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_191),
.B(n_193),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_192),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_197),
.C(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_201),
.A2(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_202),
.B(n_203),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_287),
.B(n_292),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_273),
.B(n_286),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_250),
.B(n_272),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_230),
.B(n_249),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_210),
.B(n_220),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_236)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_225),
.C(n_227),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_226),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_228),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_237),
.B(n_248),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_236),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_242),
.B(n_247),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_251),
.B(n_252),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_263),
.B1(n_270),
.B2(n_271),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_258),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_262),
.C(n_271),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_260),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_263),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_267),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_274),
.B(n_275),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_282),
.C(n_284),
.Y(n_288)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_311),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_311),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_309),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_303),
.B1(n_313),
.B2(n_316),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_305),
.C(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_316),
.C(n_317),
.Y(n_324)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_313),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_320),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_333),
.B(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);


endmodule