module real_aes_6052_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1106;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_357;
wire n_635;
wire n_792;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_1113;
wire n_852;
wire n_766;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_1034;
wire n_923;
wire n_952;
wire n_429;
wire n_976;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_1021;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_626;
wire n_400;
wire n_539;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_1072;
wire n_370;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_1053;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_1025;
wire n_409;
wire n_781;
wire n_860;
wire n_748;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_769;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_756;
wire n_713;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_334;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_1105;
wire n_902;
wire n_853;
wire n_1079;
wire n_843;
wire n_810;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1028;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_1090;
wire n_359;
wire n_456;
wire n_717;
wire n_982;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_1045;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1102;
wire n_1076;
wire n_463;
wire n_661;
wire n_396;
wire n_804;
wire n_1101;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_0), .A2(n_210), .B1(n_454), .B2(n_463), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_1), .A2(n_5), .B1(n_801), .B2(n_802), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_2), .A2(n_159), .B1(n_455), .B2(n_461), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_3), .A2(n_164), .B1(n_604), .B2(n_605), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_4), .A2(n_120), .B1(n_457), .B2(n_458), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_6), .A2(n_132), .B1(n_382), .B2(n_387), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_7), .A2(n_265), .B1(n_455), .B2(n_461), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g753 ( .A1(n_8), .A2(n_207), .B1(n_573), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_9), .A2(n_272), .B1(n_423), .B2(n_1079), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_10), .A2(n_135), .B1(n_576), .B2(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g684 ( .A(n_11), .Y(n_684) );
INVx1_ASAP7_75t_SL g933 ( .A(n_12), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_13), .A2(n_74), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_14), .A2(n_280), .B1(n_382), .B2(n_471), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_15), .A2(n_253), .B1(n_398), .B2(n_414), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_16), .B(n_342), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_17), .A2(n_212), .B1(n_805), .B2(n_806), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_18), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_19), .A2(n_197), .B1(n_457), .B2(n_458), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_20), .A2(n_139), .B1(n_573), .B2(n_574), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_21), .A2(n_169), .B1(n_441), .B2(n_464), .Y(n_608) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_22), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_23), .A2(n_75), .B1(n_865), .B2(n_867), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g1082 ( .A1(n_24), .A2(n_281), .B1(n_370), .B2(n_574), .Y(n_1082) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_25), .A2(n_119), .B1(n_478), .B2(n_479), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_26), .A2(n_181), .B1(n_513), .B2(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g634 ( .A(n_27), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_28), .A2(n_588), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_29), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_30), .A2(n_189), .B1(n_850), .B2(n_854), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_31), .A2(n_76), .B1(n_463), .B2(n_464), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_32), .A2(n_168), .B1(n_583), .B2(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_33), .A2(n_309), .B1(n_441), .B2(n_464), .Y(n_663) );
XOR2x2_ASAP7_75t_L g593 ( .A(n_34), .B(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_35), .A2(n_298), .B1(n_442), .B2(n_654), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_36), .A2(n_42), .B1(n_583), .B2(n_584), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_37), .A2(n_118), .B1(n_382), .B2(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g894 ( .A(n_38), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_39), .A2(n_84), .B1(n_411), .B2(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g787 ( .A(n_40), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_41), .A2(n_106), .B1(n_411), .B2(n_414), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_43), .A2(n_133), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_44), .A2(n_146), .B1(n_476), .B2(n_756), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_45), .A2(n_81), .B1(n_457), .B2(n_458), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_46), .A2(n_157), .B1(n_573), .B2(n_624), .Y(n_623) );
OA22x2_ASAP7_75t_L g348 ( .A1(n_47), .A2(n_131), .B1(n_342), .B2(n_346), .Y(n_348) );
INVx1_ASAP7_75t_L g377 ( .A(n_47), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_48), .A2(n_258), .B1(n_478), .B2(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_49), .A2(n_252), .B1(n_335), .B2(n_360), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_50), .A2(n_53), .B1(n_457), .B2(n_458), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_51), .A2(n_248), .B1(n_604), .B2(n_605), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_52), .A2(n_295), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_54), .A2(n_203), .B1(n_444), .B2(n_445), .Y(n_610) );
INVx1_ASAP7_75t_L g507 ( .A(n_55), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_56), .A2(n_80), .B1(n_604), .B2(n_781), .Y(n_1110) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_57), .A2(n_152), .B1(n_596), .B2(n_598), .C(n_599), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_58), .B(n_147), .Y(n_322) );
INVx1_ASAP7_75t_L g345 ( .A(n_58), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g378 ( .A1(n_58), .A2(n_131), .B(n_379), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_59), .A2(n_1094), .B1(n_1095), .B2(n_1096), .Y(n_1093) );
CKINVDCx5p33_ASAP7_75t_R g1094 ( .A(n_59), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_60), .A2(n_292), .B1(n_457), .B2(n_458), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_61), .A2(n_249), .B1(n_442), .B2(n_444), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_62), .A2(n_93), .B1(n_517), .B2(n_518), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_63), .A2(n_114), .B1(n_365), .B2(n_479), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_64), .A2(n_150), .B1(n_365), .B2(n_1109), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_65), .A2(n_121), .B1(n_568), .B2(n_569), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_66), .A2(n_278), .B1(n_564), .B2(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_67), .B(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_68), .B(n_484), .Y(n_514) );
INVx1_ASAP7_75t_L g843 ( .A(n_69), .Y(n_843) );
AND2x4_ASAP7_75t_L g851 ( .A(n_69), .B(n_223), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_70), .A2(n_261), .B1(n_441), .B2(n_464), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_71), .A2(n_191), .B1(n_387), .B2(n_479), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_72), .A2(n_167), .B1(n_536), .B2(n_569), .Y(n_705) );
INVx1_ASAP7_75t_L g493 ( .A(n_73), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_77), .A2(n_161), .B1(n_445), .B2(n_534), .Y(n_659) );
INVx1_ASAP7_75t_L g823 ( .A(n_78), .Y(n_823) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_79), .A2(n_82), .B1(n_486), .B2(n_487), .C(n_490), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_83), .A2(n_460), .B(n_786), .Y(n_785) );
XNOR2x1_ASAP7_75t_L g501 ( .A(n_85), .B(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_86), .A2(n_487), .B(n_656), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_87), .A2(n_266), .B1(n_460), .B2(n_461), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_88), .B(n_1102), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_89), .A2(n_123), .B1(n_476), .B2(n_799), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_90), .A2(n_632), .B(n_633), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_91), .A2(n_124), .B1(n_391), .B2(n_393), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_92), .A2(n_116), .B1(n_710), .B2(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g491 ( .A(n_94), .Y(n_491) );
INVx1_ASAP7_75t_L g841 ( .A(n_95), .Y(n_841) );
AND2x4_ASAP7_75t_L g846 ( .A(n_95), .B(n_318), .Y(n_846) );
INVx1_ASAP7_75t_SL g866 ( .A(n_95), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_96), .A2(n_208), .B1(n_414), .B2(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_97), .A2(n_243), .B1(n_708), .B2(n_711), .Y(n_752) );
XNOR2x2_ASAP7_75t_SL g667 ( .A(n_98), .B(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_99), .A2(n_230), .B1(n_624), .B2(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g544 ( .A(n_100), .Y(n_544) );
CKINVDCx16_ASAP7_75t_R g847 ( .A(n_101), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_102), .A2(n_122), .B1(n_839), .B2(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g427 ( .A(n_103), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_104), .A2(n_214), .B1(n_391), .B2(n_520), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_105), .A2(n_284), .B1(n_576), .B2(n_756), .Y(n_755) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_107), .A2(n_301), .B1(n_598), .B2(n_688), .C(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g891 ( .A(n_108), .Y(n_891) );
XNOR2x1_ASAP7_75t_L g645 ( .A(n_109), .B(n_646), .Y(n_645) );
OAI22x1_ASAP7_75t_L g553 ( .A1(n_110), .A2(n_554), .B1(n_590), .B2(n_591), .Y(n_553) );
NAND3xp33_ASAP7_75t_SL g590 ( .A(n_110), .B(n_570), .C(n_585), .Y(n_590) );
INVx1_ASAP7_75t_L g652 ( .A(n_111), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_112), .A2(n_145), .B1(n_454), .B2(n_463), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_113), .A2(n_299), .B1(n_457), .B2(n_458), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_115), .A2(n_513), .B(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g678 ( .A(n_117), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_125), .B(n_632), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_126), .A2(n_251), .B1(n_335), .B2(n_360), .Y(n_334) );
INVx1_ASAP7_75t_L g643 ( .A(n_127), .Y(n_643) );
CKINVDCx6p67_ASAP7_75t_R g844 ( .A(n_128), .Y(n_844) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_129), .A2(n_288), .B1(n_441), .B2(n_464), .Y(n_539) );
INVx1_ASAP7_75t_L g359 ( .A(n_130), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_130), .B(n_178), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_130), .B(n_375), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_131), .B(n_233), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_134), .A2(n_226), .B1(n_398), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_136), .A2(n_142), .B1(n_398), .B2(n_400), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_137), .A2(n_193), .B1(n_360), .B2(n_476), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_138), .A2(n_148), .B1(n_418), .B2(n_486), .C(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_140), .A2(n_260), .B1(n_808), .B2(n_809), .Y(n_807) );
INVx1_ASAP7_75t_L g1106 ( .A(n_141), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_143), .A2(n_276), .B1(n_869), .B2(n_870), .Y(n_874) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_144), .A2(n_439), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_147), .B(n_352), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_149), .A2(n_173), .B1(n_517), .B2(n_520), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_151), .A2(n_310), .B1(n_360), .B2(n_476), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_153), .A2(n_311), .B1(n_360), .B2(n_523), .Y(n_522) );
AO22x2_ASAP7_75t_L g717 ( .A1(n_154), .A2(n_718), .B1(n_737), .B2(n_738), .Y(n_717) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_154), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_154), .A2(n_238), .B1(n_869), .B2(n_870), .Y(n_868) );
INVx1_ASAP7_75t_L g657 ( .A(n_155), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_156), .A2(n_199), .B1(n_562), .B2(n_565), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_158), .A2(n_250), .B1(n_391), .B2(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_160), .B(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_162), .A2(n_209), .B1(n_506), .B2(n_792), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_163), .A2(n_290), .B1(n_398), .B2(n_1100), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_165), .A2(n_331), .B1(n_332), .B2(n_434), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_165), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_166), .A2(n_256), .B1(n_839), .B2(n_860), .Y(n_879) );
XNOR2x1_ASAP7_75t_L g775 ( .A(n_170), .B(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_171), .A2(n_302), .B1(n_815), .B2(n_816), .Y(n_814) );
BUFx2_ASAP7_75t_L g726 ( .A(n_172), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_174), .A2(n_287), .B1(n_865), .B2(n_867), .Y(n_873) );
INVx1_ASAP7_75t_L g1071 ( .A(n_174), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_174), .A2(n_1091), .B1(n_1093), .B2(n_1113), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_175), .A2(n_231), .B1(n_854), .B2(n_878), .Y(n_902) );
INVx1_ASAP7_75t_L g527 ( .A(n_176), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_177), .A2(n_286), .B1(n_517), .B2(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g343 ( .A(n_178), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_179), .A2(n_202), .B1(n_628), .B2(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_180), .B(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_182), .A2(n_201), .B1(n_523), .B2(n_626), .Y(n_625) );
XNOR2x1_ASAP7_75t_L g435 ( .A(n_183), .B(n_436), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_183), .A2(n_188), .B1(n_858), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_184), .A2(n_228), .B1(n_536), .B2(n_765), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_185), .A2(n_192), .B1(n_506), .B2(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_186), .B(n_439), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_187), .A2(n_270), .B1(n_471), .B2(n_781), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_190), .A2(n_246), .B1(n_473), .B2(n_573), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_194), .A2(n_211), .B1(n_454), .B2(n_463), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_195), .A2(n_259), .B1(n_365), .B2(n_370), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_196), .A2(n_245), .B1(n_455), .B2(n_461), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_198), .A2(n_220), .B1(n_839), .B2(n_860), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_200), .A2(n_262), .B1(n_513), .B2(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_204), .A2(n_240), .B1(n_444), .B2(n_445), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_205), .A2(n_241), .B1(n_517), .B2(n_520), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_206), .A2(n_294), .B1(n_370), .B2(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_213), .B(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_215), .A2(n_304), .B1(n_697), .B2(n_698), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g1085 ( .A1(n_216), .A2(n_306), .B1(n_382), .B2(n_393), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_217), .A2(n_218), .B1(n_536), .B2(n_819), .C(n_822), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_219), .A2(n_254), .B1(n_454), .B2(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g686 ( .A(n_221), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_222), .A2(n_239), .B1(n_850), .B2(n_858), .Y(n_857) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_223), .Y(n_323) );
AND2x4_ASAP7_75t_L g842 ( .A(n_223), .B(n_843), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_224), .B(n_418), .Y(n_417) );
XNOR2x2_ASAP7_75t_L g795 ( .A(n_225), .B(n_796), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_227), .A2(n_305), .B1(n_565), .B2(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g509 ( .A(n_229), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_232), .A2(n_274), .B1(n_442), .B2(n_460), .Y(n_609) );
INVx1_ASAP7_75t_L g357 ( .A(n_233), .Y(n_357) );
INVxp67_ASAP7_75t_L g409 ( .A(n_233), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_234), .B(n_565), .Y(n_1077) );
AOI21xp33_ASAP7_75t_SL g720 ( .A1(n_235), .A2(n_534), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g600 ( .A(n_236), .Y(n_600) );
INVx1_ASAP7_75t_L g549 ( .A(n_237), .Y(n_549) );
AOI22xp5_ASAP7_75t_SL g585 ( .A1(n_242), .A2(n_282), .B1(n_586), .B2(n_588), .Y(n_585) );
INVxp67_ASAP7_75t_R g852 ( .A(n_244), .Y(n_852) );
INVx2_ASAP7_75t_L g318 ( .A(n_247), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_255), .A2(n_257), .B1(n_441), .B2(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g690 ( .A(n_263), .Y(n_690) );
INVx1_ASAP7_75t_L g722 ( .A(n_264), .Y(n_722) );
AOI21xp33_ASAP7_75t_L g446 ( .A1(n_267), .A2(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_268), .Y(n_449) );
INVx1_ASAP7_75t_L g511 ( .A(n_269), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_271), .B(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_273), .A2(n_300), .B1(n_576), .B2(n_578), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_275), .A2(n_285), .B1(n_414), .B2(n_654), .Y(n_788) );
OAI21xp5_ASAP7_75t_L g749 ( .A1(n_277), .A2(n_750), .B(n_769), .Y(n_749) );
INVx1_ASAP7_75t_L g771 ( .A(n_277), .Y(n_771) );
INVx1_ASAP7_75t_L g892 ( .A(n_279), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_283), .A2(n_303), .B1(n_812), .B2(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g550 ( .A(n_289), .Y(n_550) );
BUFx2_ASAP7_75t_L g729 ( .A(n_291), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_293), .A2(n_307), .B1(n_479), .B2(n_518), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_296), .A2(n_489), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g934 ( .A(n_297), .Y(n_934) );
AOI21xp33_ASAP7_75t_SL g422 ( .A1(n_308), .A2(n_423), .B(n_426), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_324), .B(n_829), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx4_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .C(n_323), .Y(n_315) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_316), .B(n_1088), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_316), .B(n_1089), .Y(n_1092) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OA21x2_ASAP7_75t_L g1114 ( .A1(n_317), .A2(n_866), .B(n_1115), .Y(n_1114) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g840 ( .A(n_318), .B(n_841), .Y(n_840) );
AND3x4_ASAP7_75t_L g865 ( .A(n_318), .B(n_842), .C(n_866), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g1088 ( .A(n_319), .B(n_1089), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_320), .A2(n_431), .B(n_432), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g1089 ( .A(n_323), .Y(n_1089) );
XNOR2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_614), .Y(n_324) );
XOR2x2_ASAP7_75t_SL g325 ( .A(n_326), .B(n_496), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_329), .B1(n_465), .B2(n_494), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
XOR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_435), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_331), .A2(n_849), .B1(n_852), .B2(n_853), .Y(n_848) );
INVx1_ASAP7_75t_L g434 ( .A(n_332), .Y(n_434) );
NAND4xp75_ASAP7_75t_L g332 ( .A(n_333), .B(n_380), .C(n_396), .D(n_416), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_364), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g577 ( .A(n_336), .Y(n_577) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx12f_ASAP7_75t_L g476 ( .A(n_337), .Y(n_476) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_337), .Y(n_523) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_349), .Y(n_337) );
AND2x2_ASAP7_75t_L g361 ( .A(n_338), .B(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g366 ( .A(n_338), .B(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g392 ( .A(n_338), .B(n_385), .Y(n_392) );
AND2x4_ASAP7_75t_L g441 ( .A(n_338), .B(n_389), .Y(n_441) );
AND2x4_ASAP7_75t_L g454 ( .A(n_338), .B(n_385), .Y(n_454) );
AND2x4_ASAP7_75t_L g457 ( .A(n_338), .B(n_349), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_338), .B(n_362), .Y(n_458) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_347), .Y(n_338) );
AND2x2_ASAP7_75t_L g413 ( .A(n_339), .B(n_348), .Y(n_413) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g384 ( .A(n_340), .B(n_348), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
NAND2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx2_ASAP7_75t_L g346 ( .A(n_342), .Y(n_346) );
INVx3_ASAP7_75t_L g352 ( .A(n_342), .Y(n_352) );
NAND2xp33_ASAP7_75t_L g358 ( .A(n_342), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g379 ( .A(n_342), .Y(n_379) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_342), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_343), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g408 ( .A1(n_345), .A2(n_379), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g407 ( .A(n_348), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g399 ( .A(n_349), .B(n_384), .Y(n_399) );
AND2x4_ASAP7_75t_L g425 ( .A(n_349), .B(n_413), .Y(n_425) );
AND2x4_ASAP7_75t_L g444 ( .A(n_349), .B(n_384), .Y(n_444) );
AND2x4_ASAP7_75t_L g460 ( .A(n_349), .B(n_413), .Y(n_460) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_354), .Y(n_349) );
INVx2_ASAP7_75t_L g363 ( .A(n_350), .Y(n_363) );
OR2x2_ASAP7_75t_L g368 ( .A(n_350), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g385 ( .A(n_350), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g403 ( .A(n_350), .B(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_352), .B(n_357), .Y(n_356) );
INVxp67_ASAP7_75t_L g375 ( .A(n_352), .Y(n_375) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_353), .B(n_374), .C(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g362 ( .A(n_354), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g369 ( .A(n_355), .Y(n_369) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g581 ( .A(n_361), .Y(n_581) );
BUFx5_ASAP7_75t_L g626 ( .A(n_361), .Y(n_626) );
BUFx3_ASAP7_75t_L g756 ( .A(n_361), .Y(n_756) );
AND2x4_ASAP7_75t_L g412 ( .A(n_362), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g415 ( .A(n_362), .B(n_373), .Y(n_415) );
AND2x2_ASAP7_75t_L g421 ( .A(n_362), .B(n_384), .Y(n_421) );
AND2x4_ASAP7_75t_L g442 ( .A(n_362), .B(n_373), .Y(n_442) );
AND2x2_ASAP7_75t_L g447 ( .A(n_362), .B(n_413), .Y(n_447) );
AND2x2_ASAP7_75t_L g489 ( .A(n_362), .B(n_384), .Y(n_489) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_366), .Y(n_478) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_366), .Y(n_518) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_366), .Y(n_672) );
AND2x4_ASAP7_75t_L g372 ( .A(n_367), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g455 ( .A(n_367), .B(n_384), .Y(n_455) );
AND2x4_ASAP7_75t_L g464 ( .A(n_367), .B(n_373), .Y(n_464) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g389 ( .A(n_368), .Y(n_389) );
INVx1_ASAP7_75t_L g386 ( .A(n_369), .Y(n_386) );
INVx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g708 ( .A(n_371), .Y(n_708) );
INVx5_ASAP7_75t_L g779 ( .A(n_371), .Y(n_779) );
INVx2_ASAP7_75t_L g1109 ( .A(n_371), .Y(n_1109) );
INVx6_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx12f_ASAP7_75t_L g479 ( .A(n_372), .Y(n_479) );
AND2x4_ASAP7_75t_L g395 ( .A(n_373), .B(n_385), .Y(n_395) );
AND2x4_ASAP7_75t_L g463 ( .A(n_373), .B(n_385), .Y(n_463) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_378), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_390), .Y(n_380) );
BUFx3_ASAP7_75t_L g805 ( .A(n_382), .Y(n_805) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx8_ASAP7_75t_L g573 ( .A(n_383), .Y(n_573) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AND2x4_ASAP7_75t_L g388 ( .A(n_384), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g461 ( .A(n_384), .B(n_385), .Y(n_461) );
AND2x2_ASAP7_75t_L g606 ( .A(n_384), .B(n_385), .Y(n_606) );
BUFx3_ASAP7_75t_L g754 ( .A(n_387), .Y(n_754) );
BUFx12f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_388), .Y(n_471) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_388), .Y(n_574) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_388), .Y(n_604) );
BUFx3_ASAP7_75t_L g624 ( .A(n_388), .Y(n_624) );
BUFx2_ASAP7_75t_SL g801 ( .A(n_391), .Y(n_801) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx12f_ASAP7_75t_L g517 ( .A(n_392), .Y(n_517) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_392), .Y(n_628) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx4_ASAP7_75t_L g473 ( .A(n_394), .Y(n_473) );
INVx2_ASAP7_75t_L g520 ( .A(n_394), .Y(n_520) );
INVx4_ASAP7_75t_L g584 ( .A(n_394), .Y(n_584) );
INVx1_ASAP7_75t_L g629 ( .A(n_394), .Y(n_629) );
INVx1_ASAP7_75t_L g650 ( .A(n_394), .Y(n_650) );
INVx8_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_410), .Y(n_396) );
INVx2_ASAP7_75t_L g587 ( .A(n_398), .Y(n_587) );
BUFx2_ASAP7_75t_L g813 ( .A(n_398), .Y(n_813) );
BUFx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_399), .Y(n_506) );
INVx2_ASAP7_75t_L g642 ( .A(n_399), .Y(n_642) );
INVx4_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx3_ASAP7_75t_L g536 ( .A(n_401), .Y(n_536) );
INVx2_ASAP7_75t_L g568 ( .A(n_401), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_401), .A2(n_634), .B(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g1100 ( .A(n_401), .Y(n_1100) );
INVx5_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx4f_ASAP7_75t_L g484 ( .A(n_402), .Y(n_484) );
BUFx2_ASAP7_75t_L g792 ( .A(n_402), .Y(n_792) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_407), .Y(n_402) );
AND2x2_ASAP7_75t_L g445 ( .A(n_403), .B(n_407), .Y(n_445) );
AND2x4_ASAP7_75t_L g681 ( .A(n_403), .B(n_407), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
BUFx3_ASAP7_75t_L g815 ( .A(n_411), .Y(n_815) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx3_ASAP7_75t_L g486 ( .A(n_412), .Y(n_486) );
BUFx8_ASAP7_75t_SL g546 ( .A(n_412), .Y(n_546) );
INVx2_ASAP7_75t_L g566 ( .A(n_412), .Y(n_566) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_412), .Y(n_654) );
INVx3_ASAP7_75t_L g508 ( .A(n_414), .Y(n_508) );
BUFx3_ASAP7_75t_L g768 ( .A(n_414), .Y(n_768) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_415), .Y(n_564) );
INVx3_ASAP7_75t_L g817 ( .A(n_415), .Y(n_817) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_422), .Y(n_416) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g560 ( .A(n_420), .Y(n_560) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g439 ( .A(n_421), .Y(n_439) );
INVx3_ASAP7_75t_L g597 ( .A(n_421), .Y(n_597) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx3_ASAP7_75t_L g483 ( .A(n_425), .Y(n_483) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_425), .Y(n_513) );
BUFx3_ASAP7_75t_L g534 ( .A(n_425), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_428), .B(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_428), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_428), .B(n_787), .Y(n_786) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_429), .Y(n_637) );
INVx2_ASAP7_75t_L g763 ( .A(n_429), .Y(n_763) );
INVx1_ASAP7_75t_L g1076 ( .A(n_429), .Y(n_1076) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g451 ( .A(n_430), .Y(n_451) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_452), .Y(n_436) );
NAND4xp25_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .C(n_443), .D(n_446), .Y(n_437) );
BUFx3_ASAP7_75t_L g632 ( .A(n_439), .Y(n_632) );
INVx1_ASAP7_75t_L g704 ( .A(n_439), .Y(n_704) );
INVx2_ASAP7_75t_L g685 ( .A(n_442), .Y(n_685) );
INVx1_ASAP7_75t_L g683 ( .A(n_444), .Y(n_683) );
INVx2_ASAP7_75t_L g730 ( .A(n_444), .Y(n_730) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_447), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx4_ASAP7_75t_L g529 ( .A(n_450), .Y(n_529) );
INVx1_ASAP7_75t_L g569 ( .A(n_450), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_450), .B(n_600), .Y(n_599) );
INVx4_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g492 ( .A(n_451), .Y(n_492) );
NAND4xp25_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .C(n_459), .D(n_462), .Y(n_452) );
INVx2_ASAP7_75t_L g679 ( .A(n_460), .Y(n_679) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g495 ( .A(n_467), .Y(n_495) );
XNOR2x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_493), .Y(n_467) );
NAND4xp75_ASAP7_75t_L g468 ( .A(n_469), .B(n_474), .C(n_480), .D(n_485), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_472), .Y(n_469) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
BUFx3_ASAP7_75t_L g711 ( .A(n_478), .Y(n_711) );
BUFx3_ASAP7_75t_L g809 ( .A(n_479), .Y(n_809) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
BUFx2_ASAP7_75t_L g812 ( .A(n_483), .Y(n_812) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_489), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_492), .B(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_492), .B(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_492), .B(n_823), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_498), .B1(n_551), .B2(n_613), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
XNOR2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_530), .Y(n_500) );
NAND4xp75_ASAP7_75t_L g502 ( .A(n_503), .B(n_515), .C(n_521), .D(n_525), .Y(n_502) );
NOR2xp67_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_514), .Y(n_510) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
BUFx12f_ASAP7_75t_L g583 ( .A(n_517), .Y(n_583) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_517), .Y(n_710) );
BUFx3_ASAP7_75t_L g808 ( .A(n_518), .Y(n_808) );
BUFx2_ASAP7_75t_SL g802 ( .A(n_520), .Y(n_802) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_524), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
XOR2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_550), .Y(n_530) );
NOR4xp75_ASAP7_75t_L g531 ( .A(n_532), .B(n_537), .C(n_540), .D(n_543), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
INVx2_ASAP7_75t_L g589 ( .A(n_534), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OAI21x1_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_545), .B(n_547), .Y(n_543) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
AO22x2_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B1(n_592), .B2(n_612), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_570), .C(n_585), .Y(n_555) );
INVx1_ASAP7_75t_L g591 ( .A(n_556), .Y(n_591) );
AND3x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .C(n_567), .Y(n_556) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx4_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g698 ( .A(n_564), .Y(n_698) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g639 ( .A(n_566), .Y(n_639) );
AND4x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .C(n_575), .D(n_582), .Y(n_570) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_574), .Y(n_806) );
BUFx4f_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_580), .Y(n_713) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_593), .Y(n_612) );
NAND3x1_ASAP7_75t_L g594 ( .A(n_595), .B(n_601), .C(n_607), .Y(n_594) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g790 ( .A(n_597), .Y(n_790) );
INVx2_ASAP7_75t_L g821 ( .A(n_597), .Y(n_821) );
INVx2_ASAP7_75t_L g1075 ( .A(n_597), .Y(n_1075) );
INVx2_ASAP7_75t_L g1102 ( .A(n_597), .Y(n_1102) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx4f_ASAP7_75t_L g781 ( .A(n_606), .Y(n_781) );
AND4x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .C(n_610), .D(n_611), .Y(n_607) );
XOR2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_742), .Y(n_614) );
XNOR2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_664), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
XNOR2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_644), .Y(n_618) );
XNOR2x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_643), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_630), .Y(n_620) );
NAND4xp25_ASAP7_75t_SL g621 ( .A(n_622), .B(n_623), .C(n_625), .D(n_627), .Y(n_621) );
BUFx3_ASAP7_75t_L g799 ( .A(n_626), .Y(n_799) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_638), .C(n_640), .Y(n_630) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g1105 ( .A(n_637), .B(n_1106), .Y(n_1105) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_642), .Y(n_701) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND4xp75_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .C(n_658), .D(n_661), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
OA21x2_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_655), .Y(n_651) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
BUFx3_ASAP7_75t_L g697 ( .A(n_654), .Y(n_697) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_691), .B1(n_692), .B2(n_741), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g741 ( .A(n_667), .Y(n_741) );
NAND4xp75_ASAP7_75t_L g668 ( .A(n_669), .B(n_673), .C(n_676), .D(n_687), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_682), .Y(n_676) );
OAI21xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B(n_680), .Y(n_677) );
INVx4_ASAP7_75t_L g727 ( .A(n_681), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_685), .B2(n_686), .Y(n_682) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OA22x2_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_716), .B1(n_739), .B2(n_740), .Y(n_692) );
INVx1_ASAP7_75t_L g739 ( .A(n_693), .Y(n_739) );
XOR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_715), .Y(n_693) );
NOR2x1_ASAP7_75t_L g694 ( .A(n_695), .B(n_706), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_696), .B(n_699), .C(n_702), .D(n_705), .Y(n_695) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g765 ( .A(n_701), .Y(n_765) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .C(n_712), .D(n_714), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_715), .A2(n_894), .B1(n_895), .B2(n_896), .Y(n_893) );
INVx1_ASAP7_75t_L g740 ( .A(n_716), .Y(n_740) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g738 ( .A(n_718), .Y(n_738) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_732), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_723), .C(n_731), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_727), .B1(n_728), .B2(n_730), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
CKINVDCx9p33_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
NAND4xp25_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .C(n_735), .D(n_736), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_794), .B(n_824), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g828 ( .A(n_747), .Y(n_828) );
OA22x2_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B1(n_773), .B2(n_793), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_758), .Y(n_750) );
INVxp67_ASAP7_75t_L g772 ( .A(n_751), .Y(n_772) );
NAND4xp25_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .C(n_755), .D(n_757), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_758), .B(n_771), .Y(n_770) );
NAND4xp25_ASAP7_75t_L g758 ( .A(n_759), .B(n_764), .C(n_766), .D(n_767), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx3_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g793 ( .A(n_775), .Y(n_793) );
NOR2x1_ASAP7_75t_L g776 ( .A(n_777), .B(n_784), .Y(n_776) );
NAND4xp25_ASAP7_75t_L g777 ( .A(n_778), .B(n_780), .C(n_782), .D(n_783), .Y(n_777) );
NAND4xp25_ASAP7_75t_SL g784 ( .A(n_785), .B(n_788), .C(n_789), .D(n_791), .Y(n_784) );
BUFx3_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_SL g826 ( .A(n_795), .Y(n_826) );
NAND4xp75_ASAP7_75t_L g796 ( .A(n_797), .B(n_803), .C(n_810), .D(n_818), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_800), .Y(n_797) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_807), .Y(n_803) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_814), .Y(n_810) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx3_ASAP7_75t_L g1079 ( .A(n_817), .Y(n_1079) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_827), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_1062), .B1(n_1064), .B2(n_1086), .C(n_1090), .Y(n_829) );
AOI211xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_975), .B(n_1023), .C(n_1048), .Y(n_830) );
NAND5xp2_ASAP7_75t_L g831 ( .A(n_832), .B(n_910), .C(n_939), .D(n_948), .E(n_968), .Y(n_831) );
NOR3xp33_ASAP7_75t_SL g832 ( .A(n_833), .B(n_880), .C(n_898), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_861), .Y(n_834) );
INVx1_ASAP7_75t_L g960 ( .A(n_835), .Y(n_960) );
AOI221xp5_ASAP7_75t_L g976 ( .A1(n_835), .A2(n_977), .B1(n_979), .B2(n_980), .C(n_981), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_835), .B(n_907), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_835), .B(n_887), .Y(n_1042) );
AND2x2_ASAP7_75t_L g835 ( .A(n_836), .B(n_855), .Y(n_835) );
AND2x2_ASAP7_75t_L g897 ( .A(n_836), .B(n_856), .Y(n_897) );
INVx2_ASAP7_75t_L g914 ( .A(n_836), .Y(n_914) );
INVx3_ASAP7_75t_L g921 ( .A(n_836), .Y(n_921) );
OR2x2_ASAP7_75t_L g950 ( .A(n_836), .B(n_856), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_836), .B(n_888), .Y(n_967) );
OR2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_848), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_844), .B1(n_845), .B2(n_847), .Y(n_837) );
OAI221xp5_ASAP7_75t_L g932 ( .A1(n_838), .A2(n_845), .B1(n_933), .B2(n_934), .C(n_935), .Y(n_932) );
INVx3_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
AND2x4_ASAP7_75t_L g839 ( .A(n_840), .B(n_842), .Y(n_839) );
AND2x4_ASAP7_75t_L g850 ( .A(n_840), .B(n_851), .Y(n_850) );
AND2x2_ASAP7_75t_L g869 ( .A(n_840), .B(n_851), .Y(n_869) );
AND2x2_ASAP7_75t_L g878 ( .A(n_840), .B(n_851), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_842), .B(n_846), .Y(n_845) );
AND2x4_ASAP7_75t_L g860 ( .A(n_842), .B(n_846), .Y(n_860) );
AND2x4_ASAP7_75t_L g867 ( .A(n_842), .B(n_846), .Y(n_867) );
CKINVDCx5p33_ASAP7_75t_R g1115 ( .A(n_842), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_845), .A2(n_890), .B1(n_891), .B2(n_892), .Y(n_889) );
BUFx2_ASAP7_75t_L g1063 ( .A(n_845), .Y(n_1063) );
AND2x4_ASAP7_75t_L g854 ( .A(n_846), .B(n_851), .Y(n_854) );
AND2x2_ASAP7_75t_L g858 ( .A(n_846), .B(n_851), .Y(n_858) );
AND2x2_ASAP7_75t_L g870 ( .A(n_846), .B(n_851), .Y(n_870) );
INVx3_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_855), .B(n_900), .Y(n_899) );
INVx3_ASAP7_75t_L g930 ( .A(n_855), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_855), .B(n_901), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1061 ( .A(n_855), .B(n_901), .Y(n_1061) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
AND2x2_ASAP7_75t_L g920 ( .A(n_856), .B(n_921), .Y(n_920) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_856), .B(n_901), .Y(n_1036) );
AND2x2_ASAP7_75t_L g856 ( .A(n_857), .B(n_859), .Y(n_856) );
O2A1O1Ixp33_ASAP7_75t_L g984 ( .A1(n_861), .A2(n_974), .B(n_985), .C(n_987), .Y(n_984) );
AOI222xp33_ASAP7_75t_L g1033 ( .A1(n_861), .A2(n_1034), .B1(n_1036), .B2(n_1037), .C1(n_1038), .C2(n_1041), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_861), .B(n_887), .Y(n_1035) );
AND2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_871), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_862), .B(n_882), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_862), .B(n_884), .Y(n_942) );
AND2x2_ASAP7_75t_SL g947 ( .A(n_862), .B(n_917), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g971 ( .A(n_862), .B(n_972), .Y(n_971) );
AND2x2_ASAP7_75t_L g978 ( .A(n_862), .B(n_887), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_862), .B(n_888), .Y(n_997) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_862), .B(n_875), .Y(n_1009) );
A2O1A1Ixp33_ASAP7_75t_L g1043 ( .A1(n_862), .A2(n_1044), .B(n_1045), .C(n_1046), .Y(n_1043) );
CKINVDCx6p67_ASAP7_75t_R g862 ( .A(n_863), .Y(n_862) );
AND2x2_ASAP7_75t_L g909 ( .A(n_863), .B(n_871), .Y(n_909) );
AND2x2_ASAP7_75t_L g916 ( .A(n_863), .B(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g925 ( .A(n_863), .Y(n_925) );
OR2x2_ASAP7_75t_L g994 ( .A(n_863), .B(n_872), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_863), .B(n_884), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_863), .B(n_979), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_863), .B(n_872), .Y(n_1053) );
AND2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_868), .Y(n_863) );
INVx1_ASAP7_75t_L g890 ( .A(n_865), .Y(n_890) );
INVx2_ASAP7_75t_SL g905 ( .A(n_867), .Y(n_905) );
INVx1_ASAP7_75t_L g896 ( .A(n_869), .Y(n_896) );
INVx1_ASAP7_75t_L g895 ( .A(n_870), .Y(n_895) );
INVx1_ASAP7_75t_L g1021 ( .A(n_871), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_871), .B(n_917), .Y(n_1044) );
AND2x2_ASAP7_75t_L g871 ( .A(n_872), .B(n_875), .Y(n_871) );
AND2x2_ASAP7_75t_L g882 ( .A(n_872), .B(n_876), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g885 ( .A(n_872), .Y(n_885) );
AND2x4_ASAP7_75t_SL g872 ( .A(n_873), .B(n_874), .Y(n_872) );
AND2x2_ASAP7_75t_L g884 ( .A(n_875), .B(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g923 ( .A(n_875), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_875), .B(n_924), .Y(n_951) );
AND2x2_ASAP7_75t_L g966 ( .A(n_875), .B(n_924), .Y(n_966) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AND2x2_ASAP7_75t_L g917 ( .A(n_876), .B(n_885), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_877), .B(n_879), .Y(n_876) );
AOI21xp33_ASAP7_75t_L g880 ( .A1(n_881), .A2(n_883), .B(n_886), .Y(n_880) );
INVx1_ASAP7_75t_L g1029 ( .A(n_881), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_881), .B(n_1056), .Y(n_1055) );
AND2x2_ASAP7_75t_L g962 ( .A(n_882), .B(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g972 ( .A(n_882), .Y(n_972) );
AND2x2_ASAP7_75t_L g979 ( .A(n_882), .B(n_888), .Y(n_979) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_882), .B(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
AND2x2_ASAP7_75t_L g958 ( .A(n_884), .B(n_888), .Y(n_958) );
OAI321xp33_ASAP7_75t_L g996 ( .A1(n_884), .A2(n_922), .A3(n_961), .B1(n_995), .B2(n_997), .C(n_998), .Y(n_996) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_884), .B(n_963), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_885), .B(n_924), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_897), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_887), .B(n_928), .Y(n_927) );
AND2x2_ASAP7_75t_L g963 ( .A(n_887), .B(n_924), .Y(n_963) );
NOR2x1p5_ASAP7_75t_L g993 ( .A(n_887), .B(n_994), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_887), .B(n_930), .Y(n_1007) );
INVx1_ASAP7_75t_L g1018 ( .A(n_887), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1059 ( .A(n_887), .B(n_921), .Y(n_1059) );
CKINVDCx6p67_ASAP7_75t_R g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g908 ( .A(n_888), .Y(n_908) );
AND2x2_ASAP7_75t_L g915 ( .A(n_888), .B(n_916), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_888), .B(n_951), .Y(n_986) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_888), .B(n_921), .Y(n_999) );
NOR2xp33_ASAP7_75t_L g1020 ( .A(n_888), .B(n_1021), .Y(n_1020) );
OR2x6_ASAP7_75t_SL g888 ( .A(n_889), .B(n_893), .Y(n_888) );
INVx1_ASAP7_75t_L g982 ( .A(n_897), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_897), .B(n_901), .Y(n_1047) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_906), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g940 ( .A(n_899), .B(n_907), .Y(n_940) );
INVx1_ASAP7_75t_L g1054 ( .A(n_899), .Y(n_1054) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_900), .B(n_938), .Y(n_937) );
INVx2_ASAP7_75t_L g955 ( .A(n_900), .Y(n_955) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_900), .Y(n_1000) );
INVx3_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g944 ( .A(n_901), .Y(n_944) );
AND2x2_ASAP7_75t_L g974 ( .A(n_901), .B(n_949), .Y(n_974) );
AND2x4_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
INVx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_909), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_907), .B(n_920), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_907), .B(n_947), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_907), .B(n_966), .Y(n_1028) );
INVx3_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g1056 ( .A(n_909), .Y(n_1056) );
OAI21xp33_ASAP7_75t_L g910 ( .A1(n_911), .A2(n_918), .B(n_936), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_915), .Y(n_912) );
INVx2_ASAP7_75t_L g980 ( .A(n_913), .Y(n_980) );
BUFx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_914), .B(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g1003 ( .A(n_914), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_914), .B(n_1031), .Y(n_1030) );
NOR2xp33_ASAP7_75t_L g1052 ( .A(n_914), .B(n_1053), .Y(n_1052) );
AND2x2_ASAP7_75t_L g977 ( .A(n_917), .B(n_978), .Y(n_977) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_919), .A2(n_922), .B1(n_926), .B2(n_929), .C(n_931), .Y(n_918) );
INVx1_ASAP7_75t_L g1010 ( .A(n_920), .Y(n_1010) );
O2A1O1Ixp33_ASAP7_75t_L g1024 ( .A1(n_920), .A2(n_1025), .B(n_1029), .C(n_1030), .Y(n_1024) );
INVx1_ASAP7_75t_L g992 ( .A(n_921), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_921), .B(n_955), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_921), .B(n_962), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_922), .B(n_942), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g987 ( .A(n_922), .B(n_988), .Y(n_987) );
O2A1O1Ixp33_ASAP7_75t_L g1016 ( .A1(n_922), .A2(n_1017), .B(n_1019), .C(n_1022), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_924), .B(n_958), .Y(n_1004) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_927), .B(n_1027), .Y(n_1026) );
OAI22xp33_ASAP7_75t_L g1006 ( .A1(n_928), .A2(n_1007), .B1(n_1008), .B2(n_1010), .Y(n_1006) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_929), .B(n_965), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g981 ( .A1(n_929), .A2(n_938), .B1(n_970), .B2(n_982), .C(n_983), .Y(n_981) );
INVx3_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_930), .A2(n_957), .B1(n_959), .B2(n_961), .Y(n_956) );
INVx1_ASAP7_75t_L g995 ( .A(n_930), .Y(n_995) );
OAI221xp5_ASAP7_75t_L g1048 ( .A1(n_930), .A2(n_953), .B1(n_1049), .B2(n_1050), .C(n_1051), .Y(n_1048) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
BUFx3_ASAP7_75t_L g938 ( .A(n_932), .Y(n_938) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_941), .B1(n_943), .B2(n_945), .Y(n_939) );
INVx1_ASAP7_75t_L g1022 ( .A(n_943), .Y(n_1022) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
AOI311xp33_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_951), .A3(n_952), .B(n_956), .C(n_964), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_951), .B(n_967), .Y(n_983) );
OAI211xp5_ASAP7_75t_L g1023 ( .A1(n_952), .A2(n_1024), .B(n_1033), .C(n_1043), .Y(n_1023) );
INVx3_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_953), .B(n_960), .Y(n_959) );
INVx3_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_954), .B(n_1059), .Y(n_1058) );
INVx3_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_962), .B(n_1003), .Y(n_1050) );
AOI21xp33_ASAP7_75t_L g1060 ( .A1(n_965), .A2(n_1013), .B(n_1061), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_966), .B(n_967), .Y(n_965) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_970), .B(n_973), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
NAND5xp2_ASAP7_75t_L g975 ( .A(n_976), .B(n_984), .C(n_989), .D(n_1001), .E(n_1005), .Y(n_975) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_988), .B(n_1058), .Y(n_1057) );
A2O1A1Ixp33_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_995), .B(n_996), .C(n_1000), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_993), .Y(n_991) );
INVx1_ASAP7_75t_L g1032 ( .A(n_997), .Y(n_1032) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1000), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1004), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1003), .B(n_1039), .Y(n_1038) );
AOI221xp5_ASAP7_75t_L g1005 ( .A1(n_1006), .A2(n_1011), .B1(n_1012), .B2(n_1014), .C(n_1016), .Y(n_1005) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
CKINVDCx14_ASAP7_75t_R g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVxp67_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1054), .B1(n_1055), .B2(n_1057), .C(n_1060), .Y(n_1051) );
BUFx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVxp67_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
XNOR2xp5_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1072), .Y(n_1069) );
CKINVDCx5p33_ASAP7_75t_R g1070 ( .A(n_1071), .Y(n_1070) );
NOR2x1_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1081), .Y(n_1072) );
NAND4xp25_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1077), .C(n_1078), .D(n_1080), .Y(n_1073) );
NAND4xp25_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1083), .C(n_1084), .D(n_1085), .Y(n_1081) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
BUFx2_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
NOR2xp67_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1107), .Y(n_1097) );
NAND4xp25_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1101), .C(n_1103), .D(n_1104), .Y(n_1098) );
NAND4xp25_ASAP7_75t_SL g1107 ( .A(n_1108), .B(n_1110), .C(n_1111), .D(n_1112), .Y(n_1107) );
BUFx2_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
endmodule