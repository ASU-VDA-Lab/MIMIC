module fake_netlist_6_4896_n_1989 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1989);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1989;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1851;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1890;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_60),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_120),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_124),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_35),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_36),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_38),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_9),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_17),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_121),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_23),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_194),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_72),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_97),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_43),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_187),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_59),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_22),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_38),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_138),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_40),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_64),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_81),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_100),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_145),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_76),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_195),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_98),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_96),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_63),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_61),
.Y(n_236)
);

BUFx8_ASAP7_75t_SL g237 ( 
.A(n_12),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_42),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_86),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_87),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_165),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_131),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_45),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_170),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_126),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_29),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_42),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_119),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_30),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_130),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_78),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_57),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_49),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_46),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_180),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_19),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_122),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_70),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_21),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_28),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_40),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_54),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_22),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_134),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_5),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_32),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_12),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_70),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_142),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_162),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_103),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_58),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_58),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_99),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_143),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_75),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_20),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_62),
.Y(n_282)
);

BUFx8_ASAP7_75t_SL g283 ( 
.A(n_16),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_175),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_71),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_36),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_65),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_104),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_71),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_34),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_108),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_33),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_8),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_146),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_105),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_24),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_101),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_54),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_110),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_59),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_74),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_160),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_139),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_88),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_183),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_148),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_147),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_82),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_178),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_129),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_21),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_51),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_118),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_114),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_192),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_155),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_179),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_63),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_31),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_37),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_64),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_17),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_123),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_115),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_125),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_157),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_0),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_68),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_158),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_23),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_186),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_6),
.Y(n_332)
);

BUFx2_ASAP7_75t_SL g333 ( 
.A(n_109),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_79),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_133),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_73),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_41),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_90),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_31),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_116),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_6),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_136),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_185),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_56),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_69),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_111),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_161),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_73),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_15),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_50),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_20),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_95),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_176),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_189),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_94),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_173),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_113),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_191),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_76),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_75),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_10),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_15),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_61),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_48),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_117),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_18),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_77),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_137),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_84),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_7),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_7),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_57),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_83),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_28),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_10),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_151),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_80),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_1),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_3),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_39),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_37),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_60),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_135),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_152),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_3),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_8),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_66),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_2),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_14),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_52),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_35),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_92),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_181),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_0),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_236),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_236),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_251),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_291),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_237),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_279),
.B(n_1),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_236),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_236),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_226),
.B(n_2),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_236),
.Y(n_404)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_203),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_283),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_236),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_229),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_386),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_199),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_226),
.B(n_4),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_309),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_321),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_201),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_225),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_229),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_205),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_321),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_209),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_203),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_211),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_215),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_217),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_321),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_224),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_321),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_279),
.B(n_213),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_225),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_227),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_212),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_213),
.B(n_4),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_273),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_321),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_321),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_262),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_230),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_231),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_R g440 ( 
.A(n_273),
.B(n_305),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_305),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_297),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_206),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_239),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_262),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_240),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_241),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_297),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_242),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_244),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_249),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_200),
.B(n_5),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_262),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_262),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_257),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_212),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_259),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_200),
.B(n_9),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_262),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_340),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_363),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_363),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_200),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_221),
.B(n_11),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_363),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_221),
.B(n_11),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_266),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_228),
.B(n_13),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_372),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_372),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_275),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_284),
.Y(n_474)
);

INVxp33_ASAP7_75t_SL g475 ( 
.A(n_202),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_372),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_212),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_294),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g479 ( 
.A(n_206),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_295),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_200),
.B(n_13),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_372),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_372),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_268),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_268),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_292),
.B(n_14),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_292),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_299),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_349),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_303),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_349),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_212),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_456),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_395),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_456),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_395),
.B(n_235),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_456),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_396),
.B(n_235),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_456),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_456),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_401),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_432),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_432),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_432),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_465),
.B(n_228),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_465),
.B(n_232),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_232),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_452),
.B(n_278),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_477),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_477),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_429),
.B(n_266),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_404),
.B(n_278),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_477),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_400),
.B(n_285),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_406),
.B(n_233),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_404),
.Y(n_521)
);

AND3x2_ASAP7_75t_L g522 ( 
.A(n_403),
.B(n_323),
.C(n_313),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_313),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_408),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_492),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_408),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_492),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_415),
.B(n_323),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_420),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_420),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_426),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_428),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_437),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_428),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_435),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_435),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_436),
.B(n_233),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_436),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_437),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_411),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_445),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_445),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_406),
.B(n_245),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_453),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_453),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_417),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_454),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_454),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_459),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_430),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_459),
.B(n_245),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_460),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_452),
.B(n_247),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_406),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_460),
.B(n_247),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_434),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_461),
.B(n_252),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_463),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_463),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_464),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_464),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_467),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_467),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_476),
.Y(n_569)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_481),
.A2(n_267),
.B(n_252),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_476),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_483),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_549),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_550),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_539),
.B(n_409),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_519),
.A2(n_413),
.B1(n_410),
.B2(n_451),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_539),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_516),
.B(n_475),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_516),
.B(n_412),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_523),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_523),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_536),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_501),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_536),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_549),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_519),
.B(n_416),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_549),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_552),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_544),
.A2(n_285),
.B1(n_254),
.B2(n_281),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_513),
.A2(n_557),
.B1(n_481),
.B2(n_458),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_513),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_558),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_552),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_558),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_522),
.Y(n_595)
);

OAI22xp33_ASAP7_75t_L g596 ( 
.A1(n_544),
.A2(n_469),
.B1(n_409),
.B2(n_400),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_542),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_520),
.B(n_442),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_510),
.B(n_471),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_513),
.A2(n_458),
.B1(n_466),
.B2(n_433),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_513),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_501),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_536),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_510),
.B(n_472),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_531),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_542),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_513),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_542),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_531),
.B(n_419),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_536),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_536),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_531),
.B(n_421),
.Y(n_613)
);

INVxp33_ASAP7_75t_L g614 ( 
.A(n_550),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_542),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_510),
.B(n_470),
.C(n_468),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_542),
.Y(n_617)
);

NAND3xp33_ASAP7_75t_L g618 ( 
.A(n_510),
.B(n_483),
.C(n_486),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_557),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_494),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_513),
.A2(n_462),
.B1(n_486),
.B2(n_482),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_513),
.A2(n_256),
.B1(n_405),
.B2(n_214),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_511),
.B(n_423),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_531),
.B(n_424),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_544),
.B(n_469),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_543),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_557),
.A2(n_256),
.B1(n_214),
.B2(n_248),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_543),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_543),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_543),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_494),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_501),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_511),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_494),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_543),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_545),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_497),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_545),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_550),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_511),
.B(n_425),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_545),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_511),
.B(n_427),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_520),
.B(n_431),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_497),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_501),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_557),
.A2(n_238),
.B1(n_261),
.B2(n_255),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_512),
.B(n_438),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_512),
.B(n_439),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_520),
.B(n_547),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_552),
.Y(n_650)
);

AND3x2_ASAP7_75t_L g651 ( 
.A(n_550),
.B(n_443),
.C(n_269),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_501),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_564),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_522),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_SL g655 ( 
.A(n_520),
.B(n_441),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_512),
.B(n_444),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_497),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_512),
.B(n_446),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_547),
.B(n_447),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_547),
.B(n_422),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_547),
.Y(n_661)
);

BUFx8_ASAP7_75t_SL g662 ( 
.A(n_554),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_545),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_501),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_501),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_503),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_555),
.A2(n_362),
.B1(n_479),
.B2(n_207),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_564),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_503),
.Y(n_669)
);

CKINVDCx16_ASAP7_75t_R g670 ( 
.A(n_554),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_557),
.B(n_449),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_523),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_564),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_503),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_565),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_545),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_551),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_504),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_570),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_504),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_570),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_523),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_570),
.B(n_333),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_504),
.B(n_450),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_505),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_501),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_501),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_555),
.B(n_455),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_555),
.B(n_457),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_505),
.B(n_473),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_554),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_505),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_559),
.A2(n_208),
.B1(n_216),
.B2(n_210),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_508),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_R g695 ( 
.A(n_554),
.B(n_399),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_559),
.A2(n_218),
.B1(n_220),
.B2(n_219),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_570),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_551),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_541),
.A2(n_339),
.B1(n_348),
.B2(n_198),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_508),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_559),
.B(n_333),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_565),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_565),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_523),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_541),
.A2(n_345),
.B1(n_289),
.B2(n_261),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_508),
.B(n_474),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_521),
.B(n_480),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_562),
.B(n_490),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_566),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_521),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_521),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_524),
.B(n_422),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_523),
.B(n_212),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_524),
.Y(n_714)
);

AND3x2_ASAP7_75t_L g715 ( 
.A(n_560),
.B(n_443),
.C(n_269),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_514),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_524),
.Y(n_717)
);

INVx5_ASAP7_75t_L g718 ( 
.A(n_523),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_562),
.B(n_267),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_514),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_526),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_500),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_689),
.B(n_526),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_695),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_625),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_661),
.B(n_529),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_598),
.B(n_422),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_633),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_625),
.B(n_560),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_633),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_573),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_590),
.B(n_529),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_649),
.B(n_529),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_633),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_649),
.B(n_598),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_578),
.A2(n_488),
.B1(n_478),
.B2(n_397),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_576),
.B(n_560),
.C(n_407),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_585),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_582),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_591),
.B(n_347),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_600),
.A2(n_414),
.B1(n_398),
.B2(n_288),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_575),
.B(n_592),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_591),
.B(n_347),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_585),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_643),
.B(n_530),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_599),
.B(n_605),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_582),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_623),
.B(n_530),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_640),
.A2(n_288),
.B1(n_306),
.B2(n_274),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_587),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_587),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_660),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_693),
.A2(n_541),
.B(n_562),
.C(n_499),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_642),
.B(n_530),
.Y(n_754)
);

OAI221xp5_ASAP7_75t_L g755 ( 
.A1(n_705),
.A2(n_322),
.B1(n_366),
.B2(n_319),
.C(n_312),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_647),
.B(n_533),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_586),
.B(n_688),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_648),
.B(n_533),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_656),
.B(n_533),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_658),
.B(n_537),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_591),
.B(n_347),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_708),
.B(n_560),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_588),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_671),
.B(n_537),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_682),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_619),
.A2(n_306),
.B1(n_326),
.B2(n_274),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_591),
.B(n_537),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_588),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_592),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_601),
.B(n_540),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_584),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_601),
.B(n_347),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_584),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_593),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_593),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_594),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_616),
.B(n_448),
.C(n_223),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_579),
.B(n_302),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_594),
.B(n_448),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_682),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_719),
.B(n_540),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_601),
.B(n_540),
.Y(n_782)
);

INVxp33_ASAP7_75t_L g783 ( 
.A(n_577),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_650),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_601),
.B(n_566),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_608),
.B(n_566),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_608),
.B(n_571),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_575),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_608),
.B(n_347),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_574),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_608),
.B(n_571),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_595),
.A2(n_307),
.B1(n_308),
.B2(n_304),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_619),
.B(n_681),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_604),
.B(n_611),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_655),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_611),
.B(n_572),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_639),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_612),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_L g799 ( 
.A(n_618),
.B(n_496),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_612),
.B(n_572),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_660),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_650),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_606),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_722),
.B(n_534),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_684),
.B(n_222),
.Y(n_805)
);

INVxp33_ASAP7_75t_L g806 ( 
.A(n_699),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_719),
.B(n_534),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_719),
.B(n_534),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_653),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_620),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_719),
.B(n_534),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_690),
.B(n_234),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_616),
.A2(n_343),
.B1(n_353),
.B2(n_326),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_670),
.B(n_271),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_622),
.B(n_484),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_706),
.B(n_534),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_619),
.A2(n_701),
.B1(n_654),
.B2(n_595),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_707),
.B(n_534),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_679),
.B(n_373),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_631),
.B(n_534),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_682),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_631),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_634),
.B(n_535),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_619),
.B(n_373),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_L g825 ( 
.A(n_670),
.B(n_246),
.C(n_243),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_653),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_634),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_668),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_637),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_681),
.A2(n_391),
.B(n_289),
.C(n_287),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_637),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_668),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_644),
.B(n_657),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_644),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_L g835 ( 
.A(n_679),
.B(n_373),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_657),
.B(n_535),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_683),
.A2(n_358),
.B1(n_354),
.B2(n_383),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_666),
.B(n_535),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_666),
.B(n_535),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_691),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_683),
.A2(n_358),
.B1(n_354),
.B2(n_383),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_681),
.B(n_373),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_669),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_701),
.B(n_484),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_610),
.B(n_250),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_654),
.A2(n_352),
.B1(n_310),
.B2(n_314),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_L g847 ( 
.A(n_596),
.B(n_258),
.C(n_253),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_669),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_613),
.B(n_260),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_662),
.Y(n_850)
);

OAI221xp5_ASAP7_75t_L g851 ( 
.A1(n_646),
.A2(n_627),
.B1(n_621),
.B2(n_699),
.C(n_589),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_697),
.B(n_373),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_683),
.A2(n_697),
.B1(n_701),
.B2(n_618),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_674),
.B(n_535),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_674),
.B(n_535),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_678),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_678),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_701),
.A2(n_365),
.B1(n_353),
.B2(n_343),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_680),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_659),
.A2(n_324),
.B1(n_315),
.B2(n_316),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_624),
.B(n_263),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_614),
.B(n_264),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_680),
.B(n_535),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_685),
.B(n_561),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_692),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_692),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_697),
.B(n_317),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_694),
.B(n_561),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_683),
.A2(n_365),
.B1(n_523),
.B2(n_276),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_701),
.A2(n_683),
.B1(n_696),
.B2(n_667),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_651),
.B(n_265),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_694),
.B(n_561),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_700),
.B(n_710),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_589),
.Y(n_874)
);

OR2x6_ASAP7_75t_SL g875 ( 
.A(n_712),
.B(n_270),
.Y(n_875)
);

BUFx5_ASAP7_75t_L g876 ( 
.A(n_682),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_700),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_710),
.B(n_561),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_711),
.A2(n_325),
.B1(n_329),
.B2(n_331),
.Y(n_879)
);

NOR2x1p5_ASAP7_75t_L g880 ( 
.A(n_715),
.B(n_272),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_711),
.B(n_335),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_714),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_714),
.B(n_338),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_SL g884 ( 
.A(n_580),
.B(n_378),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_717),
.B(n_561),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_717),
.B(n_721),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_673),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_723),
.B(n_721),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_765),
.A2(n_821),
.B(n_780),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_745),
.B(n_673),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_851),
.A2(n_271),
.B(n_277),
.C(n_276),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_735),
.B(n_675),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_765),
.A2(n_665),
.B(n_664),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_765),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_765),
.A2(n_665),
.B(n_664),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_727),
.B(n_204),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_765),
.A2(n_665),
.B(n_664),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_780),
.A2(n_665),
.B(n_664),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_746),
.B(n_675),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_748),
.B(n_702),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_780),
.A2(n_664),
.B(n_632),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_740),
.A2(n_703),
.B(n_702),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_876),
.B(n_632),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_780),
.A2(n_664),
.B(n_632),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_769),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_842),
.A2(n_852),
.B(n_808),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_754),
.B(n_703),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_780),
.A2(n_632),
.B(n_716),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_757),
.A2(n_359),
.B(n_301),
.C(n_298),
.Y(n_909)
);

NOR3xp33_ASAP7_75t_L g910 ( 
.A(n_778),
.B(n_286),
.C(n_280),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_731),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_756),
.B(n_709),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_731),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_758),
.B(n_709),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_856),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_876),
.B(n_821),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_759),
.B(n_583),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_856),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_813),
.A2(n_388),
.B1(n_330),
.B2(n_298),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_790),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_870),
.A2(n_287),
.B(n_282),
.C(n_277),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_742),
.B(n_290),
.Y(n_922)
);

BUFx12f_ASAP7_75t_L g923 ( 
.A(n_850),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_760),
.B(n_583),
.Y(n_924)
);

NOR3xp33_ASAP7_75t_L g925 ( 
.A(n_741),
.B(n_762),
.C(n_797),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_821),
.A2(n_632),
.B(n_716),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_821),
.A2(n_632),
.B(n_716),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_738),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_842),
.A2(n_602),
.B(n_583),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_805),
.B(n_602),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_812),
.B(n_602),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_845),
.B(n_296),
.C(n_293),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_779),
.B(n_603),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_852),
.A2(n_645),
.B(n_603),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_807),
.A2(n_645),
.B(n_603),
.Y(n_935)
);

O2A1O1Ixp5_ASAP7_75t_L g936 ( 
.A1(n_824),
.A2(n_720),
.B(n_496),
.C(n_517),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_819),
.A2(n_645),
.B(n_603),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_776),
.Y(n_938)
);

INVx11_ASAP7_75t_L g939 ( 
.A(n_783),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_882),
.B(n_645),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_728),
.B(n_652),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_730),
.B(n_652),
.Y(n_942)
);

AOI33xp33_ASAP7_75t_L g943 ( 
.A1(n_815),
.A2(n_385),
.A3(n_282),
.B1(n_330),
.B2(n_332),
.B3(n_334),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_817),
.A2(n_342),
.B1(n_346),
.B2(n_355),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_876),
.B(n_652),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_725),
.B(n_394),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_738),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_734),
.B(n_652),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_752),
.B(n_686),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_724),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_884),
.A2(n_356),
.B1(n_357),
.B2(n_368),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_867),
.A2(n_369),
.B1(n_376),
.B2(n_377),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_801),
.B(n_332),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_819),
.A2(n_687),
.B(n_686),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_830),
.A2(n_496),
.B(n_499),
.C(n_528),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_876),
.B(n_686),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_811),
.A2(n_687),
.B(n_607),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_801),
.B(n_687),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_744),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_806),
.B(n_687),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_835),
.A2(n_720),
.B(n_713),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_742),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_835),
.A2(n_732),
.B(n_793),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_776),
.B(n_204),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_764),
.B(n_720),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_793),
.A2(n_720),
.B(n_581),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_799),
.A2(n_818),
.B(n_816),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_806),
.B(n_300),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_853),
.A2(n_499),
.B1(n_528),
.B2(n_517),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_840),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_744),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_876),
.B(n_580),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_830),
.A2(n_517),
.B(n_528),
.C(n_351),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_810),
.B(n_597),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_788),
.B(n_311),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_781),
.A2(n_824),
.B(n_804),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_753),
.A2(n_351),
.B(n_334),
.C(n_345),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_749),
.A2(n_359),
.B(n_366),
.C(n_388),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_767),
.A2(n_581),
.B(n_580),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_876),
.B(n_580),
.Y(n_980)
);

NOR3xp33_ASAP7_75t_L g981 ( 
.A(n_849),
.B(n_320),
.C(n_318),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_858),
.A2(n_385),
.B(n_379),
.C(n_391),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_770),
.A2(n_581),
.B(n_580),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_820),
.A2(n_836),
.B(n_823),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_750),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_782),
.A2(n_581),
.B(n_580),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_837),
.A2(n_841),
.B1(n_733),
.B2(n_833),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_861),
.A2(n_607),
.B(n_609),
.C(n_615),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_785),
.A2(n_672),
.B(n_581),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_822),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_827),
.B(n_597),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_876),
.B(n_581),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_829),
.B(n_607),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_750),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_867),
.A2(n_766),
.B(n_886),
.C(n_873),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_831),
.B(n_609),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_834),
.B(n_609),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_755),
.A2(n_379),
.B(n_327),
.C(n_344),
.Y(n_998)
);

AND2x2_ASAP7_75t_SL g999 ( 
.A(n_847),
.B(n_485),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_781),
.B(n_672),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_729),
.B(n_328),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_794),
.A2(n_617),
.B(n_615),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_803),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_843),
.B(n_617),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_795),
.B(n_672),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_729),
.B(n_336),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_777),
.A2(n_630),
.B(n_698),
.C(n_677),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_751),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_814),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_814),
.B(n_337),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_862),
.A2(n_341),
.B(n_350),
.Y(n_1011)
);

AND3x1_ASAP7_75t_L g1012 ( 
.A(n_737),
.B(n_485),
.C(n_487),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_881),
.A2(n_636),
.B(n_677),
.C(n_676),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_848),
.B(n_626),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_857),
.B(n_626),
.Y(n_1015)
);

BUFx8_ASAP7_75t_L g1016 ( 
.A(n_840),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_786),
.A2(n_718),
.B(n_704),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_859),
.B(n_626),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_783),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_815),
.A2(n_375),
.B(n_380),
.C(n_374),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_787),
.A2(n_718),
.B(n_704),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_844),
.B(n_487),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_844),
.A2(n_393),
.B1(n_384),
.B2(n_392),
.Y(n_1023)
);

CKINVDCx11_ASAP7_75t_R g1024 ( 
.A(n_803),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_871),
.A2(n_382),
.B(n_361),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_795),
.B(n_360),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_724),
.B(n_364),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_791),
.A2(n_718),
.B(n_704),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_751),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_865),
.B(n_628),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_866),
.B(n_628),
.Y(n_1031)
);

AO21x1_ASAP7_75t_L g1032 ( 
.A1(n_740),
.A2(n_698),
.B(n_676),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_736),
.B(n_204),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_763),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_881),
.A2(n_698),
.B(n_676),
.C(n_663),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_877),
.B(n_628),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_743),
.A2(n_718),
.B(n_704),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_726),
.A2(n_771),
.B1(n_739),
.B2(n_798),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_L g1039 ( 
.A(n_747),
.B(n_523),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_763),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_773),
.B(n_768),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_874),
.B(n_370),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_850),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_792),
.A2(n_371),
.B(n_390),
.Y(n_1044)
);

AOI21x1_ASAP7_75t_L g1045 ( 
.A1(n_761),
.A2(n_638),
.B(n_629),
.Y(n_1045)
);

AOI21xp33_ASAP7_75t_L g1046 ( 
.A1(n_874),
.A2(n_381),
.B(n_387),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_875),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_825),
.B(n_489),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_883),
.B(n_389),
.Y(n_1049)
);

OR2x6_ASAP7_75t_L g1050 ( 
.A(n_880),
.B(n_489),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_869),
.A2(n_636),
.B1(n_630),
.B2(n_635),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_768),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_774),
.B(n_672),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_883),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_838),
.A2(n_630),
.B(n_635),
.C(n_636),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_761),
.A2(n_718),
.B(n_704),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_772),
.A2(n_638),
.B(n_635),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_774),
.B(n_638),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_775),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_839),
.A2(n_663),
.B(n_641),
.Y(n_1060)
);

AO21x1_ASAP7_75t_L g1061 ( 
.A1(n_772),
.A2(n_789),
.B(n_796),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_789),
.A2(n_718),
.B(n_704),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_846),
.B(n_16),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_775),
.B(n_641),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_784),
.B(n_672),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_784),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_875),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_800),
.A2(n_500),
.B(n_493),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_920),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_963),
.A2(n_854),
.B(n_863),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_915),
.B(n_918),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_SL g1072 ( 
.A(n_923),
.B(n_802),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_925),
.A2(n_879),
.B1(n_860),
.B2(n_887),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_915),
.B(n_809),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_888),
.B(n_826),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_939),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_1019),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_918),
.B(n_894),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_SL g1079 ( 
.A(n_1003),
.B(n_826),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_1049),
.A2(n_885),
.B(n_878),
.C(n_872),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1009),
.B(n_828),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_947),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_894),
.B(n_828),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_970),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_1042),
.B(n_832),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_L g1086 ( 
.A(n_1046),
.B(n_491),
.C(n_855),
.Y(n_1086)
);

O2A1O1Ixp5_ASAP7_75t_L g1087 ( 
.A1(n_1061),
.A2(n_832),
.B(n_868),
.C(n_864),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_947),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_889),
.A2(n_500),
.B(n_493),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_899),
.B(n_532),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_SL g1091 ( 
.A(n_1043),
.B(n_491),
.Y(n_1091)
);

BUFx2_ASAP7_75t_SL g1092 ( 
.A(n_970),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_906),
.B(n_532),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_916),
.A2(n_500),
.B(n_495),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_916),
.A2(n_500),
.B(n_495),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_R g1096 ( 
.A(n_950),
.B(n_85),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_1024),
.B(n_89),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1022),
.B(n_93),
.Y(n_1098)
);

AO32x2_ASAP7_75t_L g1099 ( 
.A1(n_969),
.A2(n_987),
.A3(n_1038),
.B1(n_1051),
.B2(n_921),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_1016),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_938),
.B(n_532),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_995),
.B(n_532),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1045),
.A2(n_567),
.B(n_563),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_990),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_903),
.A2(n_967),
.B(n_895),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1001),
.B(n_561),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1042),
.B(n_18),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_890),
.B(n_561),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_905),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_900),
.A2(n_567),
.B1(n_563),
.B2(n_551),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_903),
.A2(n_493),
.B(n_495),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_1006),
.B(n_563),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1049),
.A2(n_523),
.B1(n_567),
.B2(n_563),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_962),
.B(n_946),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_922),
.B(n_563),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_893),
.A2(n_493),
.B(n_495),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1016),
.Y(n_1117)
);

NAND2x1p5_ASAP7_75t_L g1118 ( 
.A(n_1000),
.B(n_563),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1022),
.B(n_563),
.Y(n_1119)
);

NAND2xp33_ASAP7_75t_L g1120 ( 
.A(n_1054),
.B(n_523),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_976),
.B(n_532),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_960),
.A2(n_567),
.B(n_551),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_897),
.A2(n_493),
.B(n_495),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1063),
.A2(n_567),
.B(n_569),
.C(n_553),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_994),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_907),
.B(n_567),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1033),
.A2(n_569),
.B1(n_553),
.B2(n_551),
.C(n_26),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_898),
.A2(n_498),
.B(n_502),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1057),
.A2(n_498),
.B(n_502),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_960),
.A2(n_569),
.B(n_553),
.C(n_498),
.Y(n_1130)
);

AOI221x1_ASAP7_75t_L g1131 ( 
.A1(n_977),
.A2(n_569),
.B1(n_553),
.B2(n_525),
.C(n_514),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_908),
.A2(n_498),
.B(n_502),
.Y(n_1132)
);

AOI21x1_ASAP7_75t_L g1133 ( 
.A1(n_902),
.A2(n_569),
.B(n_553),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_912),
.B(n_506),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_919),
.A2(n_523),
.B1(n_556),
.B2(n_548),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_921),
.A2(n_527),
.B(n_518),
.C(n_515),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1041),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_914),
.A2(n_498),
.B1(n_502),
.B2(n_548),
.Y(n_1138)
);

AOI21x1_ASAP7_75t_L g1139 ( 
.A1(n_930),
.A2(n_502),
.B(n_515),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1001),
.B(n_19),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_946),
.B(n_968),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_926),
.A2(n_506),
.B(n_507),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1050),
.B(n_102),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_927),
.A2(n_506),
.B(n_507),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1027),
.B(n_24),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1052),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_892),
.A2(n_568),
.B1(n_556),
.B2(n_548),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_SL g1148 ( 
.A1(n_1005),
.A2(n_515),
.B(n_518),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_896),
.B(n_506),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1043),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_999),
.B(n_532),
.Y(n_1151)
);

O2A1O1Ixp5_ASAP7_75t_SL g1152 ( 
.A1(n_1067),
.A2(n_506),
.B(n_507),
.C(n_509),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1005),
.A2(n_568),
.B1(n_556),
.B2(n_548),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1020),
.A2(n_515),
.B(n_518),
.C(n_527),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_994),
.Y(n_1155)
);

NOR3xp33_ASAP7_75t_SL g1156 ( 
.A(n_1027),
.B(n_25),
.C(n_26),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1059),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_901),
.A2(n_506),
.B(n_507),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1010),
.B(n_506),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_904),
.A2(n_507),
.B(n_509),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1010),
.B(n_25),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_931),
.A2(n_568),
.B1(n_556),
.B2(n_548),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1066),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_945),
.A2(n_507),
.B(n_509),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_SL g1165 ( 
.A1(n_910),
.A2(n_507),
.B(n_509),
.C(n_527),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1026),
.B(n_891),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_945),
.A2(n_956),
.B(n_972),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_956),
.A2(n_509),
.B(n_527),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_972),
.A2(n_509),
.B(n_527),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_999),
.B(n_532),
.Y(n_1170)
);

AO21x1_ASAP7_75t_L g1171 ( 
.A1(n_973),
.A2(n_933),
.B(n_955),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_980),
.A2(n_509),
.B(n_515),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_964),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1034),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_919),
.A2(n_523),
.B1(n_556),
.B2(n_548),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1041),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1026),
.A2(n_518),
.B(n_538),
.C(n_532),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_981),
.A2(n_523),
.B1(n_556),
.B2(n_548),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_980),
.A2(n_518),
.B(n_514),
.Y(n_1179)
);

AND2x6_ASAP7_75t_L g1180 ( 
.A(n_1048),
.B(n_514),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_891),
.B(n_538),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_975),
.B(n_27),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_917),
.B(n_538),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1034),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1047),
.B(n_568),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_924),
.B(n_538),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_992),
.A2(n_514),
.B(n_525),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_975),
.B(n_953),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1011),
.B(n_27),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_SL g1190 ( 
.A(n_1025),
.B(n_568),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_977),
.A2(n_514),
.B(n_525),
.Y(n_1191)
);

BUFx2_ASAP7_75t_SL g1192 ( 
.A(n_953),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_992),
.A2(n_514),
.B(n_525),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1000),
.B(n_538),
.Y(n_1194)
);

NAND3xp33_ASAP7_75t_SL g1195 ( 
.A(n_932),
.B(n_29),
.C(n_30),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1020),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1050),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1044),
.B(n_39),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_909),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_909),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1023),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1050),
.B(n_47),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_965),
.A2(n_514),
.B(n_525),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_943),
.B(n_538),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_935),
.A2(n_525),
.B(n_538),
.Y(n_1205)
);

O2A1O1Ixp5_ASAP7_75t_L g1206 ( 
.A1(n_1032),
.A2(n_132),
.B(n_197),
.C(n_188),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_940),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_998),
.A2(n_538),
.B(n_532),
.C(n_548),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_957),
.A2(n_525),
.B(n_538),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_998),
.A2(n_532),
.B(n_556),
.C(n_548),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1012),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_911),
.B(n_568),
.Y(n_1212)
);

OAI22x1_ASAP7_75t_L g1213 ( 
.A1(n_944),
.A2(n_951),
.B1(n_952),
.B2(n_1065),
.Y(n_1213)
);

BUFx8_ASAP7_75t_SL g1214 ( 
.A(n_913),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1013),
.A2(n_568),
.B(n_556),
.C(n_548),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1007),
.A2(n_112),
.B(n_184),
.C(n_177),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_928),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_R g1218 ( 
.A(n_1039),
.B(n_107),
.Y(n_1218)
);

CKINVDCx11_ASAP7_75t_R g1219 ( 
.A(n_928),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_959),
.B(n_568),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1105),
.A2(n_961),
.B(n_937),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1188),
.B(n_978),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1131),
.A2(n_988),
.A3(n_1055),
.B(n_954),
.Y(n_1223)
);

AOI21xp33_ASAP7_75t_L g1224 ( 
.A1(n_1141),
.A2(n_982),
.B(n_1035),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1077),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1102),
.A2(n_929),
.B(n_934),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1214),
.Y(n_1227)
);

NOR4xp25_ASAP7_75t_L g1228 ( 
.A(n_1196),
.B(n_1199),
.C(n_1200),
.D(n_1107),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1219),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1104),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1141),
.A2(n_949),
.B(n_958),
.C(n_1065),
.Y(n_1231)
);

OA22x2_ASAP7_75t_L g1232 ( 
.A1(n_1069),
.A2(n_1053),
.B1(n_971),
.B2(n_985),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1102),
.A2(n_1002),
.B(n_966),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1152),
.A2(n_936),
.B(n_984),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1070),
.A2(n_1159),
.B(n_1075),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1080),
.A2(n_1015),
.B(n_974),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1215),
.A2(n_1060),
.B(n_1068),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1079),
.B(n_971),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1171),
.A2(n_1014),
.B(n_1018),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1107),
.A2(n_1008),
.B1(n_1029),
.B2(n_985),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1085),
.B(n_1008),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1087),
.A2(n_1004),
.B(n_997),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1085),
.B(n_1029),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_SL g1244 ( 
.A(n_1150),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1133),
.A2(n_1058),
.B(n_1064),
.Y(n_1245)
);

NAND2x2_ASAP7_75t_L g1246 ( 
.A(n_1076),
.B(n_993),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1166),
.B(n_1040),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1129),
.A2(n_1103),
.B(n_1139),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1146),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1208),
.A2(n_1053),
.B(n_942),
.C(n_948),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_SL g1251 ( 
.A(n_1145),
.B(n_991),
.C(n_996),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1210),
.A2(n_1030),
.B(n_1036),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1167),
.A2(n_1031),
.B(n_941),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1121),
.A2(n_1028),
.B(n_979),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1121),
.A2(n_989),
.B(n_983),
.Y(n_1255)
);

OA21x2_ASAP7_75t_L g1256 ( 
.A1(n_1177),
.A2(n_1017),
.B(n_986),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1116),
.A2(n_1021),
.B(n_1056),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1145),
.A2(n_1062),
.B(n_1037),
.C(n_50),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1092),
.B(n_556),
.Y(n_1259)
);

AOI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1093),
.A2(n_568),
.B(n_546),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1109),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1093),
.A2(n_546),
.B(n_174),
.Y(n_1262)
);

AO32x2_ASAP7_75t_L g1263 ( 
.A1(n_1207),
.A2(n_47),
.A3(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_1263)
);

INVx3_ASAP7_75t_SL g1264 ( 
.A(n_1100),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1197),
.B(n_127),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1123),
.A2(n_546),
.B(n_172),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1181),
.A2(n_53),
.A3(n_55),
.B(n_56),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1182),
.A2(n_546),
.B(n_55),
.C(n_62),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1128),
.A2(n_546),
.B(n_128),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1084),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1132),
.A2(n_1209),
.B(n_1095),
.Y(n_1271)
);

AOI221xp5_ASAP7_75t_L g1272 ( 
.A1(n_1182),
.A2(n_1198),
.B1(n_1189),
.B2(n_1140),
.C(n_1161),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_1084),
.Y(n_1273)
);

INVx6_ASAP7_75t_SL g1274 ( 
.A(n_1143),
.Y(n_1274)
);

AO21x1_ASAP7_75t_L g1275 ( 
.A1(n_1189),
.A2(n_1198),
.B(n_1170),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1091),
.B(n_546),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1114),
.B(n_53),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1201),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1278)
);

AOI221xp5_ASAP7_75t_L g1279 ( 
.A1(n_1127),
.A2(n_546),
.B1(n_68),
.B2(n_69),
.C(n_72),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1192),
.A2(n_67),
.B1(n_74),
.B2(n_77),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1211),
.A2(n_546),
.B1(n_79),
.B2(n_78),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1173),
.B(n_140),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1205),
.A2(n_141),
.A3(n_149),
.B(n_153),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1149),
.A2(n_546),
.B(n_163),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_SL g1285 ( 
.A1(n_1170),
.A2(n_156),
.B(n_164),
.C(n_166),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1117),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1094),
.A2(n_169),
.B(n_171),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1111),
.A2(n_1203),
.B(n_1089),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1213),
.A2(n_1124),
.A3(n_1162),
.B(n_1138),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1206),
.A2(n_1090),
.B(n_1122),
.Y(n_1290)
);

INVx8_ASAP7_75t_L g1291 ( 
.A(n_1098),
.Y(n_1291)
);

AO21x1_ASAP7_75t_L g1292 ( 
.A1(n_1151),
.A2(n_1190),
.B(n_1073),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_SL g1293 ( 
.A1(n_1165),
.A2(n_1071),
.B(n_1078),
.C(n_1194),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1114),
.B(n_1106),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1072),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1098),
.A2(n_1157),
.B1(n_1163),
.B2(n_1143),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1090),
.A2(n_1134),
.B(n_1183),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1154),
.A2(n_1108),
.B(n_1186),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1126),
.A2(n_1078),
.B(n_1071),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1185),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1195),
.A2(n_1086),
.B1(n_1202),
.B2(n_1156),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1083),
.A2(n_1074),
.B(n_1120),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1112),
.A2(n_1115),
.B(n_1156),
.C(n_1204),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_SL g1304 ( 
.A(n_1197),
.B(n_1176),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1187),
.A2(n_1193),
.B(n_1142),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1144),
.A2(n_1179),
.B(n_1168),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1164),
.A2(n_1220),
.B(n_1160),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1137),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1119),
.A2(n_1165),
.B(n_1184),
.C(n_1081),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1158),
.A2(n_1172),
.B(n_1169),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1082),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1217),
.A2(n_1184),
.B1(n_1074),
.B2(n_1155),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1088),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1125),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1147),
.A2(n_1153),
.A3(n_1110),
.B(n_1130),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1194),
.A2(n_1212),
.B(n_1216),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1096),
.B(n_1097),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1130),
.A2(n_1101),
.B(n_1174),
.C(n_1113),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1148),
.A2(n_1136),
.B(n_1191),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1191),
.A2(n_1178),
.B(n_1118),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1118),
.A2(n_1191),
.B(n_1178),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1217),
.Y(n_1322)
);

AND2x2_ASAP7_75t_SL g1323 ( 
.A(n_1217),
.B(n_1099),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1217),
.A2(n_1099),
.B(n_1135),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1099),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1097),
.B(n_1096),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1099),
.A2(n_1135),
.B(n_1175),
.C(n_1218),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1180),
.B(n_1218),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1180),
.Y(n_1329)
);

OAI22x1_ASAP7_75t_L g1330 ( 
.A1(n_1180),
.A2(n_1107),
.B1(n_1141),
.B2(n_1182),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1175),
.A2(n_889),
.B(n_780),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1180),
.A2(n_889),
.B(n_780),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1180),
.A2(n_1133),
.B(n_1129),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1141),
.A2(n_1182),
.B(n_757),
.C(n_778),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1188),
.B(n_1141),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1141),
.A2(n_1182),
.B(n_757),
.C(n_778),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1131),
.A2(n_1171),
.A3(n_1210),
.B(n_1208),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1141),
.B(n_1085),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1105),
.A2(n_889),
.B(n_780),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1104),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1141),
.A2(n_1107),
.B(n_1145),
.C(n_1182),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1105),
.A2(n_889),
.B(n_780),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1131),
.A2(n_1171),
.A3(n_1210),
.B(n_1208),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1197),
.B(n_1084),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1131),
.A2(n_1102),
.B(n_1215),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1131),
.A2(n_1171),
.A3(n_1210),
.B(n_1208),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1077),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1131),
.A2(n_1171),
.A3(n_1210),
.B(n_1208),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1133),
.A2(n_1129),
.B(n_1103),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1069),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1105),
.A2(n_889),
.B(n_780),
.Y(n_1351)
);

AND2x6_ASAP7_75t_L g1352 ( 
.A(n_1143),
.B(n_1098),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1105),
.A2(n_889),
.B(n_780),
.Y(n_1353)
);

OAI22x1_ASAP7_75t_L g1354 ( 
.A1(n_1107),
.A2(n_1141),
.B1(n_1182),
.B2(n_1145),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1133),
.A2(n_1129),
.B(n_1103),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1105),
.A2(n_889),
.B(n_780),
.Y(n_1356)
);

OAI22x1_ASAP7_75t_L g1357 ( 
.A1(n_1107),
.A2(n_1141),
.B1(n_1182),
.B2(n_1145),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1141),
.B(n_578),
.C(n_1107),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1141),
.A2(n_1107),
.B(n_1145),
.C(n_1182),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1141),
.B(n_1085),
.Y(n_1360)
);

AOI221x1_ASAP7_75t_L g1361 ( 
.A1(n_1141),
.A2(n_1107),
.B1(n_1145),
.B2(n_1182),
.C(n_977),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1133),
.A2(n_1129),
.B(n_1103),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1131),
.A2(n_1171),
.A3(n_1210),
.B(n_1208),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1141),
.A2(n_1182),
.B(n_757),
.C(n_778),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1105),
.A2(n_889),
.B(n_780),
.Y(n_1365)
);

AOI221x1_ASAP7_75t_L g1366 ( 
.A1(n_1141),
.A2(n_1107),
.B1(n_1145),
.B2(n_1182),
.C(n_977),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1104),
.Y(n_1367)
);

NOR4xp25_ASAP7_75t_L g1368 ( 
.A(n_1196),
.B(n_1200),
.C(n_1199),
.D(n_1107),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1131),
.A2(n_1171),
.A3(n_1210),
.B(n_1208),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1141),
.B(n_1085),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1104),
.Y(n_1371)
);

AOI221xp5_ASAP7_75t_L g1372 ( 
.A1(n_1107),
.A2(n_1141),
.B1(n_576),
.B2(n_1182),
.C(n_1046),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1150),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1105),
.A2(n_889),
.B(n_780),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1152),
.A2(n_963),
.B(n_1087),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1225),
.Y(n_1376)
);

BUFx4f_ASAP7_75t_L g1377 ( 
.A(n_1229),
.Y(n_1377)
);

BUFx10_ASAP7_75t_L g1378 ( 
.A(n_1229),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1244),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1358),
.A2(n_1372),
.B1(n_1360),
.B2(n_1370),
.Y(n_1380)
);

CKINVDCx6p67_ASAP7_75t_R g1381 ( 
.A(n_1264),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1358),
.A2(n_1272),
.B1(n_1354),
.B2(n_1357),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1350),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1291),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1352),
.A2(n_1295),
.B1(n_1280),
.B2(n_1330),
.Y(n_1385)
);

BUFx12f_ASAP7_75t_L g1386 ( 
.A(n_1229),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1344),
.B(n_1270),
.Y(n_1387)
);

BUFx2_ASAP7_75t_SL g1388 ( 
.A(n_1227),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1322),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1340),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1347),
.Y(n_1391)
);

AOI22x1_ASAP7_75t_SL g1392 ( 
.A1(n_1350),
.A2(n_1341),
.B1(n_1359),
.B2(n_1249),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1367),
.Y(n_1393)
);

INVx3_ASAP7_75t_SL g1394 ( 
.A(n_1326),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1371),
.Y(n_1395)
);

AOI21xp33_ASAP7_75t_L g1396 ( 
.A1(n_1334),
.A2(n_1364),
.B(n_1336),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1335),
.B(n_1294),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1279),
.A2(n_1275),
.B1(n_1278),
.B2(n_1281),
.Y(n_1398)
);

CKINVDCx11_ASAP7_75t_R g1399 ( 
.A(n_1286),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1280),
.A2(n_1352),
.B1(n_1323),
.B2(n_1296),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1301),
.A2(n_1366),
.B(n_1361),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1352),
.A2(n_1277),
.B1(n_1296),
.B2(n_1222),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1301),
.A2(n_1304),
.B1(n_1227),
.B2(n_1326),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1352),
.A2(n_1262),
.B1(n_1291),
.B2(n_1227),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1261),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1292),
.A2(n_1224),
.B1(n_1251),
.B2(n_1262),
.Y(n_1406)
);

INVx4_ASAP7_75t_L g1407 ( 
.A(n_1270),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1373),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1291),
.Y(n_1409)
);

INVx6_ASAP7_75t_L g1410 ( 
.A(n_1270),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1317),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1224),
.A2(n_1246),
.B1(n_1274),
.B2(n_1238),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1311),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1326),
.Y(n_1414)
);

OAI21xp33_ASAP7_75t_L g1415 ( 
.A1(n_1228),
.A2(n_1368),
.B(n_1268),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1308),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1241),
.B(n_1243),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1274),
.A2(n_1300),
.B1(n_1232),
.B2(n_1265),
.Y(n_1418)
);

BUFx2_ASAP7_75t_SL g1419 ( 
.A(n_1273),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1265),
.A2(n_1247),
.B1(n_1313),
.B2(n_1314),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_1282),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1303),
.B(n_1228),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1259),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1328),
.A2(n_1327),
.B1(n_1240),
.B2(n_1309),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1304),
.A2(n_1240),
.B1(n_1324),
.B2(n_1226),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1368),
.B(n_1276),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1267),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1302),
.A2(n_1299),
.B1(n_1329),
.B2(n_1235),
.Y(n_1428)
);

INVx4_ASAP7_75t_L g1429 ( 
.A(n_1256),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1312),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1331),
.A2(n_1239),
.B1(n_1312),
.B2(n_1258),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1285),
.A2(n_1284),
.B1(n_1332),
.B2(n_1290),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1298),
.A2(n_1290),
.B1(n_1325),
.B2(n_1320),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1316),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1293),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1267),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1267),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1298),
.A2(n_1320),
.B1(n_1252),
.B2(n_1236),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1252),
.A2(n_1242),
.B1(n_1375),
.B2(n_1256),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1263),
.A2(n_1345),
.B1(n_1375),
.B2(n_1237),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1231),
.A2(n_1242),
.B1(n_1374),
.B2(n_1365),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1263),
.A2(n_1345),
.B1(n_1297),
.B2(n_1233),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1254),
.A2(n_1255),
.B1(n_1253),
.B2(n_1221),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1339),
.A2(n_1353),
.B1(n_1356),
.B2(n_1351),
.Y(n_1444)
);

BUFx2_ASAP7_75t_SL g1445 ( 
.A(n_1342),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1237),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1263),
.B(n_1283),
.Y(n_1447)
);

INVx8_ASAP7_75t_L g1448 ( 
.A(n_1318),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1287),
.Y(n_1449)
);

INVx8_ASAP7_75t_L g1450 ( 
.A(n_1283),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1234),
.A2(n_1319),
.B1(n_1321),
.B2(n_1307),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1234),
.A2(n_1319),
.B1(n_1260),
.B2(n_1348),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1337),
.B(n_1369),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1337),
.B(n_1369),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1250),
.A2(n_1266),
.B1(n_1269),
.B2(n_1310),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1283),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1289),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1289),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1343),
.A2(n_1369),
.B1(n_1363),
.B2(n_1348),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1346),
.A2(n_1363),
.B1(n_1348),
.B2(n_1289),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1346),
.B(n_1363),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1346),
.A2(n_1223),
.B1(n_1315),
.B2(n_1245),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1271),
.A2(n_1288),
.B1(n_1306),
.B2(n_1305),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1257),
.A2(n_1333),
.B1(n_1349),
.B2(n_1355),
.Y(n_1464)
);

OAI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1223),
.A2(n_1315),
.B1(n_1362),
.B2(n_1248),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1358),
.A2(n_1107),
.B1(n_1141),
.B2(n_1182),
.Y(n_1466)
);

BUFx10_ASAP7_75t_L g1467 ( 
.A(n_1229),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1358),
.A2(n_1107),
.B1(n_1141),
.B2(n_1182),
.Y(n_1468)
);

BUFx12f_ASAP7_75t_L g1469 ( 
.A(n_1229),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1350),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1230),
.Y(n_1471)
);

CKINVDCx12_ASAP7_75t_R g1472 ( 
.A(n_1326),
.Y(n_1472)
);

BUFx10_ASAP7_75t_L g1473 ( 
.A(n_1229),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1372),
.A2(n_1358),
.B1(n_1272),
.B2(n_1141),
.Y(n_1474)
);

CKINVDCx6p67_ASAP7_75t_R g1475 ( 
.A(n_1264),
.Y(n_1475)
);

INVx11_ASAP7_75t_L g1476 ( 
.A(n_1286),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1358),
.A2(n_1107),
.B1(n_1141),
.B2(n_1182),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1358),
.A2(n_1107),
.B1(n_1141),
.B2(n_1182),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1372),
.A2(n_1358),
.B1(n_1272),
.B2(n_1141),
.Y(n_1479)
);

INVx6_ASAP7_75t_L g1480 ( 
.A(n_1270),
.Y(n_1480)
);

INVx5_ASAP7_75t_L g1481 ( 
.A(n_1352),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1358),
.A2(n_1107),
.B1(n_1141),
.B2(n_1182),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1230),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1358),
.A2(n_1372),
.B1(n_1334),
.B2(n_1364),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1372),
.A2(n_1358),
.B1(n_1272),
.B2(n_1141),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1358),
.A2(n_1372),
.B1(n_1334),
.B2(n_1364),
.Y(n_1486)
);

BUFx4f_ASAP7_75t_SL g1487 ( 
.A(n_1274),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1358),
.A2(n_1372),
.B1(n_1334),
.B2(n_1364),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1372),
.A2(n_1358),
.B1(n_1272),
.B2(n_1141),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1322),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1372),
.A2(n_1141),
.B1(n_1358),
.B2(n_1107),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1230),
.Y(n_1492)
);

INVx6_ASAP7_75t_L g1493 ( 
.A(n_1270),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1225),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1358),
.A2(n_1372),
.B1(n_1360),
.B2(n_1338),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1372),
.A2(n_1358),
.B1(n_1272),
.B2(n_1141),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1225),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1225),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1372),
.A2(n_1358),
.B1(n_1272),
.B2(n_1141),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1344),
.B(n_1084),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1358),
.A2(n_1107),
.B1(n_1141),
.B2(n_1182),
.Y(n_1501)
);

CKINVDCx11_ASAP7_75t_R g1502 ( 
.A(n_1264),
.Y(n_1502)
);

OR2x6_ASAP7_75t_L g1503 ( 
.A(n_1291),
.B(n_1296),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1344),
.B(n_1137),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1358),
.A2(n_1372),
.B1(n_1334),
.B2(n_1364),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1230),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1358),
.A2(n_1107),
.B1(n_1141),
.B2(n_1182),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1230),
.Y(n_1508)
);

INVx8_ASAP7_75t_L g1509 ( 
.A(n_1291),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1372),
.A2(n_1358),
.B1(n_1272),
.B2(n_1141),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1427),
.Y(n_1511)
);

CKINVDCx14_ASAP7_75t_R g1512 ( 
.A(n_1502),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1390),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1393),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1391),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1437),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1422),
.B(n_1457),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1453),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1401),
.B(n_1447),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1395),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1503),
.B(n_1450),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1464),
.A2(n_1444),
.B(n_1441),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1454),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1471),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1458),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1461),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1494),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1483),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1460),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1459),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1380),
.B(n_1495),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1446),
.Y(n_1532)
);

AOI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1431),
.A2(n_1486),
.B(n_1484),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1492),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1383),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1503),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1506),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1503),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1508),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1382),
.B(n_1433),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1429),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1497),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1429),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1426),
.B(n_1488),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1481),
.B(n_1402),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1376),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1382),
.B(n_1505),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1481),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1481),
.B(n_1423),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1397),
.B(n_1424),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1479),
.A2(n_1510),
.B1(n_1485),
.B2(n_1499),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1479),
.A2(n_1510),
.B1(n_1485),
.B2(n_1499),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1434),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1396),
.B(n_1400),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1491),
.A2(n_1474),
.B1(n_1489),
.B2(n_1496),
.C(n_1501),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1481),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1435),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1440),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1440),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1435),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1435),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1413),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1403),
.A2(n_1380),
.B1(n_1495),
.B2(n_1394),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1400),
.B(n_1385),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1381),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1462),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1464),
.A2(n_1463),
.B(n_1443),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1462),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1439),
.A2(n_1406),
.B(n_1438),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1376),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1498),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1442),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1442),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1425),
.Y(n_1574)
);

OR2x6_ASAP7_75t_L g1575 ( 
.A(n_1445),
.B(n_1448),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1425),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1465),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1449),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1465),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1466),
.A2(n_1468),
.B1(n_1507),
.B2(n_1482),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1452),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1463),
.A2(n_1455),
.B(n_1428),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1452),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1498),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1410),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1410),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1436),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1430),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1448),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1496),
.B(n_1466),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1456),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1406),
.B(n_1415),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1451),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1470),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1417),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1432),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_SL g1597 ( 
.A1(n_1392),
.A2(n_1478),
.B1(n_1507),
.B2(n_1468),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1403),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1477),
.B(n_1482),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1504),
.Y(n_1600)
);

CKINVDCx6p67_ASAP7_75t_R g1601 ( 
.A(n_1399),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1420),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1477),
.A2(n_1501),
.B1(n_1478),
.B2(n_1398),
.Y(n_1603)
);

AOI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1500),
.A2(n_1404),
.B(n_1412),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1420),
.A2(n_1412),
.B(n_1418),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1504),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1394),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1404),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1419),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1387),
.A2(n_1490),
.B(n_1389),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1398),
.A2(n_1421),
.B(n_1405),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1472),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1384),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1389),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1411),
.A2(n_1408),
.B(n_1500),
.Y(n_1615)
);

CKINVDCx12_ASAP7_75t_R g1616 ( 
.A(n_1377),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1475),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1379),
.B(n_1414),
.Y(n_1618)
);

OAI21xp33_ASAP7_75t_L g1619 ( 
.A1(n_1416),
.A2(n_1490),
.B(n_1409),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1601),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1519),
.B(n_1388),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1595),
.B(n_1407),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1525),
.B(n_1517),
.Y(n_1623)
);

BUFx4f_ASAP7_75t_SL g1624 ( 
.A(n_1601),
.Y(n_1624)
);

O2A1O1Ixp33_ASAP7_75t_SL g1625 ( 
.A1(n_1531),
.A2(n_1377),
.B(n_1509),
.C(n_1487),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1555),
.B(n_1409),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1603),
.A2(n_1580),
.B1(n_1591),
.B2(n_1547),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1562),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1562),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_R g1630 ( 
.A(n_1545),
.B(n_1509),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1519),
.B(n_1378),
.Y(n_1631)
);

NAND2x1_ASAP7_75t_L g1632 ( 
.A(n_1575),
.B(n_1493),
.Y(n_1632)
);

NOR2x1_ASAP7_75t_SL g1633 ( 
.A(n_1575),
.B(n_1386),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1558),
.B(n_1378),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1570),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1558),
.B(n_1467),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1597),
.A2(n_1487),
.B1(n_1480),
.B2(n_1410),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1562),
.Y(n_1638)
);

OAI31xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1563),
.A2(n_1467),
.A3(n_1473),
.B(n_1469),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1551),
.A2(n_1480),
.B1(n_1476),
.B2(n_1473),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1549),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1552),
.A2(n_1590),
.B1(n_1599),
.B2(n_1554),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1559),
.B(n_1581),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1533),
.A2(n_1592),
.B(n_1605),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1608),
.B(n_1587),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1535),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_SL g1647 ( 
.A(n_1575),
.B(n_1521),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1592),
.A2(n_1554),
.B1(n_1612),
.B2(n_1564),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1544),
.A2(n_1550),
.B1(n_1591),
.B2(n_1564),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1550),
.A2(n_1587),
.B1(n_1611),
.B2(n_1612),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1533),
.A2(n_1605),
.B(n_1522),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1616),
.A2(n_1512),
.B1(n_1615),
.B2(n_1617),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1521),
.B(n_1545),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1540),
.A2(n_1576),
.B(n_1574),
.C(n_1598),
.Y(n_1654)
);

BUFx4f_ASAP7_75t_SL g1655 ( 
.A(n_1594),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1583),
.B(n_1593),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1522),
.A2(n_1540),
.B(n_1582),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1572),
.B(n_1573),
.Y(n_1658)
);

AO22x2_ASAP7_75t_L g1659 ( 
.A1(n_1566),
.A2(n_1568),
.B1(n_1577),
.B2(n_1579),
.Y(n_1659)
);

OAI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1574),
.A2(n_1576),
.B(n_1569),
.C(n_1598),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1582),
.A2(n_1596),
.B(n_1567),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1570),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1588),
.B(n_1619),
.Y(n_1663)
);

AO21x1_ASAP7_75t_L g1664 ( 
.A1(n_1609),
.A2(n_1614),
.B(n_1516),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1596),
.A2(n_1567),
.B(n_1569),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1515),
.B(n_1527),
.Y(n_1666)
);

OA21x2_ASAP7_75t_L g1667 ( 
.A1(n_1577),
.A2(n_1579),
.B(n_1568),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1532),
.B(n_1513),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1588),
.B(n_1542),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1569),
.A2(n_1604),
.B(n_1553),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1619),
.B(n_1604),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1537),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1553),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1569),
.A2(n_1602),
.B1(n_1546),
.B2(n_1584),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1553),
.A2(n_1602),
.B(n_1609),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1514),
.B(n_1520),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1536),
.B(n_1538),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_SL g1678 ( 
.A1(n_1514),
.A2(n_1539),
.B(n_1534),
.Y(n_1678)
);

OA21x2_ASAP7_75t_L g1679 ( 
.A1(n_1566),
.A2(n_1511),
.B(n_1529),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1545),
.A2(n_1560),
.B1(n_1561),
.B2(n_1557),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1520),
.B(n_1524),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1669),
.B(n_1571),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1628),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1629),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1666),
.B(n_1635),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1662),
.B(n_1516),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1643),
.B(n_1529),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1667),
.B(n_1530),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1643),
.B(n_1530),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1673),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1638),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1627),
.A2(n_1610),
.B(n_1545),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1667),
.B(n_1523),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1647),
.B(n_1536),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1642),
.A2(n_1538),
.B1(n_1561),
.B2(n_1575),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1667),
.B(n_1526),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1626),
.A2(n_1607),
.B1(n_1549),
.B2(n_1600),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_1541),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1653),
.B(n_1543),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1655),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1642),
.A2(n_1575),
.B1(n_1607),
.B2(n_1589),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1671),
.A2(n_1556),
.B1(n_1548),
.B2(n_1589),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_SL g1703 ( 
.A1(n_1650),
.A2(n_1626),
.B1(n_1671),
.B2(n_1637),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1649),
.A2(n_1549),
.B1(n_1600),
.B2(n_1606),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1653),
.B(n_1511),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1645),
.B(n_1623),
.Y(n_1706)
);

AND2x2_ASAP7_75t_SL g1707 ( 
.A(n_1674),
.B(n_1556),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1653),
.B(n_1578),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1672),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1677),
.B(n_1518),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1676),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1681),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1679),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1679),
.B(n_1518),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1677),
.B(n_1523),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1648),
.B(n_1528),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1641),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1641),
.B(n_1578),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1668),
.Y(n_1719)
);

OAI321xp33_ASAP7_75t_L g1720 ( 
.A1(n_1695),
.A2(n_1644),
.A3(n_1657),
.B1(n_1651),
.B2(n_1670),
.C(n_1674),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1711),
.B(n_1712),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_SL g1722 ( 
.A1(n_1707),
.A2(n_1652),
.B1(n_1675),
.B2(n_1663),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1688),
.B(n_1665),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1694),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1705),
.B(n_1717),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1683),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1711),
.B(n_1661),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1690),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1705),
.B(n_1717),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1683),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1713),
.Y(n_1731)
);

OAI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1703),
.A2(n_1639),
.B1(n_1654),
.B2(n_1640),
.C(n_1663),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1684),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_L g1734 ( 
.A1(n_1707),
.A2(n_1660),
.B(n_1622),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1712),
.B(n_1659),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1694),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1717),
.B(n_1659),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1716),
.B(n_1631),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1710),
.B(n_1715),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1701),
.A2(n_1654),
.B1(n_1634),
.B2(n_1636),
.Y(n_1740)
);

AO21x2_ASAP7_75t_L g1741 ( 
.A1(n_1688),
.A2(n_1664),
.B(n_1678),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1709),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1684),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1710),
.B(n_1659),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1693),
.B(n_1658),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1692),
.A2(n_1646),
.B1(n_1656),
.B2(n_1625),
.C(n_1658),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1698),
.Y(n_1747)
);

OAI31xp33_ASAP7_75t_L g1748 ( 
.A1(n_1700),
.A2(n_1625),
.A3(n_1680),
.B(n_1621),
.Y(n_1748)
);

OAI222xp33_ASAP7_75t_L g1749 ( 
.A1(n_1697),
.A2(n_1685),
.B1(n_1621),
.B2(n_1682),
.C1(n_1704),
.C2(n_1702),
.Y(n_1749)
);

INVx5_ASAP7_75t_L g1750 ( 
.A(n_1694),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1718),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1691),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1714),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1726),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1735),
.B(n_1719),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1726),
.Y(n_1756)
);

NOR2x1_ASAP7_75t_L g1757 ( 
.A(n_1741),
.B(n_1693),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1723),
.B(n_1696),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1724),
.B(n_1707),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1724),
.B(n_1702),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1724),
.B(n_1694),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1736),
.B(n_1706),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1730),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1723),
.B(n_1696),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1730),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1736),
.B(n_1706),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1735),
.B(n_1727),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1736),
.B(n_1708),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1733),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1735),
.B(n_1687),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1738),
.B(n_1620),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1723),
.B(n_1686),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1725),
.B(n_1708),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1725),
.B(n_1708),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1751),
.B(n_1718),
.Y(n_1775)
);

INVxp67_ASAP7_75t_SL g1776 ( 
.A(n_1731),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1745),
.B(n_1727),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1727),
.B(n_1687),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1733),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1745),
.B(n_1689),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1743),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1743),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1725),
.B(n_1708),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1745),
.B(n_1744),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1744),
.B(n_1689),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1725),
.B(n_1698),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1725),
.B(n_1729),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1750),
.B(n_1698),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1752),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1752),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1721),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1729),
.B(n_1698),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1729),
.B(n_1744),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1742),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1750),
.B(n_1699),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1729),
.B(n_1699),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1721),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1767),
.B(n_1728),
.Y(n_1798)
);

NAND2xp33_ASAP7_75t_L g1799 ( 
.A(n_1760),
.B(n_1620),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1754),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1772),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1754),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1767),
.B(n_1728),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1759),
.B(n_1760),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1756),
.Y(n_1805)
);

OAI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1771),
.A2(n_1722),
.B(n_1720),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1756),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1759),
.B(n_1750),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1794),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1759),
.B(n_1750),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1793),
.B(n_1750),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1762),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1763),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1772),
.B(n_1741),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1793),
.B(n_1750),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1778),
.B(n_1738),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1778),
.B(n_1739),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1763),
.Y(n_1818)
);

INVxp33_ASAP7_75t_L g1819 ( 
.A(n_1768),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1757),
.A2(n_1722),
.B(n_1720),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1773),
.B(n_1624),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1788),
.B(n_1748),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1786),
.B(n_1750),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1765),
.Y(n_1824)
);

NAND2x1_ASAP7_75t_L g1825 ( 
.A(n_1788),
.B(n_1729),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1784),
.B(n_1741),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1788),
.B(n_1748),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1786),
.B(n_1750),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1792),
.B(n_1747),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1792),
.B(n_1747),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1788),
.B(n_1795),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1765),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1762),
.B(n_1739),
.Y(n_1833)
);

INVxp33_ASAP7_75t_SL g1834 ( 
.A(n_1762),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1769),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1795),
.A2(n_1732),
.B1(n_1746),
.B2(n_1740),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1766),
.B(n_1739),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1784),
.B(n_1741),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1794),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1777),
.B(n_1741),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1769),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1779),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1779),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1822),
.Y(n_1844)
);

AND2x4_ASAP7_75t_SL g1845 ( 
.A(n_1831),
.B(n_1795),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1798),
.B(n_1777),
.Y(n_1846)
);

OAI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1820),
.A2(n_1806),
.B(n_1836),
.C(n_1827),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1804),
.B(n_1796),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1816),
.B(n_1766),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1804),
.B(n_1796),
.Y(n_1850)
);

NOR2x1_ASAP7_75t_L g1851 ( 
.A(n_1799),
.B(n_1757),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1799),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1809),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1798),
.B(n_1758),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1801),
.B(n_1803),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1812),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1803),
.B(n_1834),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1805),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1805),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1825),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1834),
.B(n_1781),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1809),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1842),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1831),
.B(n_1795),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1831),
.B(n_1773),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1829),
.B(n_1774),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1821),
.B(n_1565),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1815),
.B(n_1787),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1839),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1817),
.B(n_1833),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1800),
.B(n_1781),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1842),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1802),
.B(n_1782),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1837),
.B(n_1766),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1826),
.B(n_1758),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1829),
.B(n_1830),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1819),
.B(n_1785),
.Y(n_1877)
);

BUFx2_ASAP7_75t_L g1878 ( 
.A(n_1815),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1830),
.B(n_1808),
.Y(n_1879)
);

NAND3xp33_ASAP7_75t_L g1880 ( 
.A(n_1826),
.B(n_1732),
.C(n_1746),
.Y(n_1880)
);

INVxp67_ASAP7_75t_SL g1881 ( 
.A(n_1851),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1856),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1858),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1852),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1847),
.A2(n_1815),
.B1(n_1808),
.B2(n_1810),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1862),
.Y(n_1886)
);

NAND2xp33_ASAP7_75t_SL g1887 ( 
.A(n_1857),
.B(n_1825),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1858),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1859),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1859),
.Y(n_1890)
);

O2A1O1Ixp33_ASAP7_75t_L g1891 ( 
.A1(n_1844),
.A2(n_1749),
.B(n_1838),
.C(n_1840),
.Y(n_1891)
);

AOI321xp33_ASAP7_75t_L g1892 ( 
.A1(n_1851),
.A2(n_1740),
.A3(n_1838),
.B1(n_1810),
.B2(n_1840),
.C(n_1734),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_R g1893 ( 
.A(n_1852),
.B(n_1616),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1853),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1876),
.B(n_1785),
.Y(n_1895)
);

O2A1O1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1880),
.A2(n_1749),
.B(n_1814),
.C(n_1839),
.Y(n_1896)
);

OAI21xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1880),
.A2(n_1734),
.B(n_1811),
.Y(n_1897)
);

AOI211xp5_ASAP7_75t_L g1898 ( 
.A1(n_1855),
.A2(n_1811),
.B(n_1814),
.C(n_1823),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1876),
.B(n_1823),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1879),
.B(n_1755),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1860),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1863),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1855),
.A2(n_1618),
.B(n_1807),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1864),
.B(n_1828),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1879),
.B(n_1828),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1878),
.Y(n_1906)
);

AOI22x1_ASAP7_75t_L g1907 ( 
.A1(n_1878),
.A2(n_1761),
.B1(n_1776),
.B2(n_1764),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_SL g1908 ( 
.A1(n_1845),
.A2(n_1867),
.B(n_1864),
.Y(n_1908)
);

AOI31xp33_ASAP7_75t_L g1909 ( 
.A1(n_1884),
.A2(n_1881),
.A3(n_1906),
.B(n_1882),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1893),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_SL g1911 ( 
.A1(n_1886),
.A2(n_1860),
.B1(n_1864),
.B2(n_1861),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1886),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1903),
.B(n_1848),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1894),
.Y(n_1914)
);

AOI33xp33_ASAP7_75t_L g1915 ( 
.A1(n_1896),
.A2(n_1853),
.A3(n_1869),
.B1(n_1872),
.B2(n_1863),
.B3(n_1845),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1894),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1897),
.B(n_1848),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1891),
.A2(n_1861),
.B(n_1877),
.Y(n_1918)
);

INVxp67_ASAP7_75t_L g1919 ( 
.A(n_1887),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1883),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1888),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1905),
.B(n_1865),
.Y(n_1922)
);

OAI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1892),
.A2(n_1870),
.B1(n_1846),
.B2(n_1849),
.C(n_1860),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1899),
.B(n_1850),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1899),
.B(n_1850),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1889),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1890),
.Y(n_1927)
);

OAI322xp33_ASAP7_75t_L g1928 ( 
.A1(n_1907),
.A2(n_1846),
.A3(n_1854),
.B1(n_1869),
.B2(n_1853),
.C1(n_1872),
.C2(n_1875),
.Y(n_1928)
);

AOI21xp33_ASAP7_75t_SL g1929 ( 
.A1(n_1908),
.A2(n_1854),
.B(n_1860),
.Y(n_1929)
);

OAI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1885),
.A2(n_1874),
.B1(n_1864),
.B2(n_1869),
.Y(n_1930)
);

OAI211xp5_ASAP7_75t_L g1931 ( 
.A1(n_1929),
.A2(n_1887),
.B(n_1907),
.C(n_1898),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1912),
.Y(n_1932)
);

AOI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1909),
.A2(n_1904),
.B(n_1901),
.Y(n_1933)
);

AOI31xp33_ASAP7_75t_SL g1934 ( 
.A1(n_1911),
.A2(n_1901),
.A3(n_1895),
.B(n_1900),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1912),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1910),
.B(n_1904),
.Y(n_1936)
);

INVx1_ASAP7_75t_SL g1937 ( 
.A(n_1922),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1919),
.B(n_1905),
.Y(n_1938)
);

O2A1O1Ixp33_ASAP7_75t_L g1939 ( 
.A1(n_1928),
.A2(n_1902),
.B(n_1873),
.C(n_1871),
.Y(n_1939)
);

INVx1_ASAP7_75t_SL g1940 ( 
.A(n_1922),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1913),
.B(n_1845),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1915),
.B(n_1866),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1914),
.Y(n_1943)
);

NAND2x1_ASAP7_75t_SL g1944 ( 
.A(n_1920),
.B(n_1868),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1931),
.B(n_1915),
.Y(n_1945)
);

NOR3xp33_ASAP7_75t_L g1946 ( 
.A(n_1936),
.B(n_1917),
.C(n_1918),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1937),
.B(n_1920),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1940),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1941),
.B(n_1923),
.Y(n_1949)
);

OAI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1933),
.A2(n_1930),
.B1(n_1924),
.B2(n_1925),
.Y(n_1950)
);

NOR4xp25_ASAP7_75t_L g1951 ( 
.A(n_1934),
.B(n_1927),
.C(n_1926),
.D(n_1921),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1938),
.B(n_1916),
.Y(n_1952)
);

NAND4xp25_ASAP7_75t_L g1953 ( 
.A(n_1938),
.B(n_1868),
.C(n_1865),
.D(n_1875),
.Y(n_1953)
);

AOI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1939),
.A2(n_1873),
.B(n_1871),
.Y(n_1954)
);

AOI211xp5_ASAP7_75t_L g1955 ( 
.A1(n_1945),
.A2(n_1942),
.B(n_1935),
.C(n_1932),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1947),
.B(n_1943),
.Y(n_1956)
);

AOI222xp33_ASAP7_75t_L g1957 ( 
.A1(n_1949),
.A2(n_1944),
.B1(n_1868),
.B2(n_1866),
.C1(n_1776),
.C2(n_1843),
.Y(n_1957)
);

NOR3xp33_ASAP7_75t_L g1958 ( 
.A(n_1946),
.B(n_1868),
.C(n_1843),
.Y(n_1958)
);

AOI211xp5_ASAP7_75t_SL g1959 ( 
.A1(n_1950),
.A2(n_1841),
.B(n_1835),
.C(n_1832),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1947),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1958),
.A2(n_1948),
.B1(n_1953),
.B2(n_1951),
.Y(n_1961)
);

O2A1O1Ixp33_ASAP7_75t_L g1962 ( 
.A1(n_1955),
.A2(n_1952),
.B(n_1954),
.C(n_1824),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1956),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1960),
.B(n_1813),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1957),
.A2(n_1818),
.B1(n_1634),
.B2(n_1636),
.Y(n_1965)
);

NOR2x1_ASAP7_75t_SL g1966 ( 
.A(n_1959),
.B(n_1761),
.Y(n_1966)
);

OAI21xp5_ASAP7_75t_SL g1967 ( 
.A1(n_1959),
.A2(n_1768),
.B(n_1787),
.Y(n_1967)
);

NOR2x1_ASAP7_75t_L g1968 ( 
.A(n_1963),
.B(n_1962),
.Y(n_1968)
);

NAND4xp75_ASAP7_75t_L g1969 ( 
.A(n_1961),
.B(n_1737),
.C(n_1585),
.D(n_1586),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1966),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1964),
.B(n_1774),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1967),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1965),
.B(n_1764),
.Y(n_1973)
);

NOR3xp33_ASAP7_75t_L g1974 ( 
.A(n_1968),
.B(n_1632),
.C(n_1755),
.Y(n_1974)
);

OAI31xp33_ASAP7_75t_L g1975 ( 
.A1(n_1970),
.A2(n_1753),
.A3(n_1783),
.B(n_1747),
.Y(n_1975)
);

NAND4xp75_ASAP7_75t_L g1976 ( 
.A(n_1972),
.B(n_1737),
.C(n_1585),
.D(n_1586),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1975),
.B(n_1973),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1977),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1978),
.A2(n_1969),
.B1(n_1976),
.B2(n_1974),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1978),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1980),
.A2(n_1979),
.B1(n_1971),
.B2(n_1775),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1979),
.A2(n_1783),
.B(n_1770),
.Y(n_1982)
);

OAI21x1_ASAP7_75t_L g1983 ( 
.A1(n_1981),
.A2(n_1770),
.B(n_1789),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1982),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1780),
.B(n_1633),
.Y(n_1985)
);

OAI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1985),
.A2(n_1984),
.B(n_1983),
.Y(n_1986)
);

OAI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1986),
.A2(n_1797),
.B1(n_1791),
.B2(n_1790),
.Y(n_1987)
);

OAI221xp5_ASAP7_75t_R g1988 ( 
.A1(n_1987),
.A2(n_1630),
.B1(n_1753),
.B2(n_1790),
.C(n_1789),
.Y(n_1988)
);

AOI211xp5_ASAP7_75t_L g1989 ( 
.A1(n_1988),
.A2(n_1613),
.B(n_1548),
.C(n_1556),
.Y(n_1989)
);


endmodule