module fake_netlist_6_3273_n_591 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_591);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_591;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_581;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_311;
wire n_403;
wire n_253;
wire n_583;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

BUFx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_16),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_28),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_30),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_96),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_8),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_9),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_20),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_26),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_9),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_75),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_3),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_87),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_4),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_13),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_56),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_63),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_19),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_2),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_36),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_27),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_111),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_66),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_21),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_50),
.B(n_76),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_67),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_14),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_5),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_54),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_83),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_43),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_106),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_64),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_8),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_53),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_48),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_25),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_15),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_113),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_7),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_13),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_91),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_80),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_90),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_12),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_L g194 ( 
.A(n_71),
.B(n_100),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_29),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_118),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_157),
.Y(n_200)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_134),
.B(n_0),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_142),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_135),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_17),
.Y(n_214)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_136),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_144),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_139),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_151),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_1),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_143),
.B(n_18),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_147),
.B(n_22),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_147),
.B(n_4),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_153),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_155),
.B(n_161),
.Y(n_234)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_185),
.A2(n_186),
.B1(n_166),
.B2(n_172),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_154),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_159),
.B(n_5),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_214),
.B(n_194),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_137),
.B1(n_149),
.B2(n_187),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_160),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_214),
.B(n_141),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_162),
.Y(n_249)
);

AOI21x1_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_198),
.B(n_164),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

BUFx4f_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_214),
.B(n_150),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_218),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_209),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_170),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_205),
.A2(n_196),
.B1(n_171),
.B2(n_174),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_218),
.B(n_176),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

NOR3xp33_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_224),
.C(n_231),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_211),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_169),
.C(n_192),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_232),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_237),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_201),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_217),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_200),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_226),
.B(n_227),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_216),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_239),
.A2(n_181),
.B1(n_183),
.B2(n_169),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_227),
.B1(n_226),
.B2(n_225),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_285),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_226),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_242),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_247),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_247),
.B(n_222),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_249),
.B(n_235),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_240),
.Y(n_302)
);

O2A1O1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_240),
.A2(n_203),
.B(n_204),
.C(n_208),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_201),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_246),
.B(n_201),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_265),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_227),
.B1(n_228),
.B2(n_233),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_278),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_270),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_276),
.Y(n_312)
);

OR2x6_ASAP7_75t_L g313 ( 
.A(n_254),
.B(n_220),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g315 ( 
.A1(n_275),
.A2(n_230),
.B1(n_204),
.B2(n_208),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_257),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_247),
.B(n_235),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_244),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_283),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_258),
.B(n_229),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_258),
.B1(n_268),
.B2(n_238),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_287),
.B(n_230),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_241),
.B(n_238),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_287),
.A2(n_156),
.B1(n_165),
.B2(n_197),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_217),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_L g330 ( 
.A(n_250),
.B(n_206),
.C(n_168),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_199),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_264),
.B(n_217),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_244),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_264),
.B(n_217),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_248),
.Y(n_340)
);

OAI22x1_ASAP7_75t_R g341 ( 
.A1(n_255),
.A2(n_207),
.B1(n_191),
.B2(n_190),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_248),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_267),
.B(n_274),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_255),
.A2(n_206),
.B1(n_199),
.B2(n_202),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_277),
.B(n_175),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_295),
.B(n_282),
.Y(n_347)
);

AOI22x1_ASAP7_75t_L g348 ( 
.A1(n_295),
.A2(n_282),
.B1(n_262),
.B2(n_261),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_311),
.B(n_255),
.Y(n_349)
);

O2A1O1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_296),
.A2(n_202),
.B(n_251),
.C(n_261),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_288),
.A2(n_262),
.B(n_260),
.C(n_251),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_288),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_260),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_296),
.A2(n_184),
.B1(n_180),
.B2(n_178),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_252),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_325),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_346),
.A2(n_281),
.B(n_252),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_301),
.A2(n_177),
.B1(n_207),
.B2(n_252),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_301),
.B(n_6),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_299),
.B(n_252),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_23),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_318),
.A2(n_309),
.B1(n_298),
.B2(n_326),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_340),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_24),
.Y(n_369)
);

AOI21x1_ASAP7_75t_L g370 ( 
.A1(n_343),
.A2(n_70),
.B(n_130),
.Y(n_370)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_313),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_304),
.A2(n_69),
.B(n_129),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_330),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_315),
.B(n_10),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_305),
.A2(n_72),
.B1(n_31),
.B2(n_32),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_303),
.A2(n_11),
.B(n_33),
.C(n_34),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_320),
.A2(n_78),
.B(n_35),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_334),
.A2(n_79),
.B1(n_37),
.B2(n_38),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_335),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_297),
.B(n_11),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_330),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_320),
.A2(n_42),
.B(n_44),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_303),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_383)
);

O2A1O1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_315),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_316),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_338),
.A2(n_55),
.B(n_57),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_338),
.A2(n_58),
.B(n_59),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_317),
.B(n_60),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_328),
.A2(n_61),
.B(n_62),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_65),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_327),
.B(n_68),
.Y(n_392)
);

O2A1O1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_342),
.A2(n_339),
.B(n_337),
.C(n_324),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_292),
.B(n_74),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_289),
.Y(n_395)
);

NAND3xp33_ASAP7_75t_L g396 ( 
.A(n_319),
.B(n_77),
.C(n_81),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_291),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_293),
.A2(n_88),
.B(n_89),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_300),
.A2(n_92),
.B(n_93),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_306),
.B(n_95),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_294),
.A2(n_97),
.B(n_98),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_289),
.B(n_99),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_352),
.A2(n_333),
.B(n_344),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_358),
.B(n_329),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_362),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_314),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_380),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_356),
.A2(n_332),
.B(n_312),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_308),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_371),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_307),
.Y(n_412)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_348),
.A2(n_103),
.B(n_105),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_379),
.A2(n_341),
.B1(n_333),
.B2(n_336),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_361),
.B(n_107),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_347),
.A2(n_108),
.B(n_109),
.Y(n_416)
);

AOI221xp5_ASAP7_75t_L g417 ( 
.A1(n_374),
.A2(n_110),
.B1(n_114),
.B2(n_115),
.C(n_119),
.Y(n_417)
);

OAI21xp33_ASAP7_75t_L g418 ( 
.A1(n_354),
.A2(n_121),
.B(n_125),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_365),
.A2(n_336),
.B(n_126),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_357),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_369),
.A2(n_336),
.B(n_133),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_353),
.A2(n_336),
.B(n_393),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g423 ( 
.A1(n_366),
.A2(n_336),
.B(n_391),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_373),
.B(n_359),
.C(n_355),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_386),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_349),
.B(n_401),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_385),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_351),
.A2(n_350),
.B(n_403),
.Y(n_429)
);

AO31x2_ASAP7_75t_L g430 ( 
.A1(n_376),
.A2(n_383),
.A3(n_394),
.B(n_375),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_392),
.A2(n_395),
.B(n_384),
.Y(n_431)
);

AO21x2_ASAP7_75t_L g432 ( 
.A1(n_370),
.A2(n_387),
.B(n_388),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_360),
.A2(n_377),
.B(n_382),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_385),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_395),
.A2(n_400),
.B(n_381),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_389),
.B(n_396),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_390),
.A2(n_399),
.B(n_398),
.Y(n_437)
);

AO31x2_ASAP7_75t_L g438 ( 
.A1(n_402),
.A2(n_372),
.A3(n_378),
.B(n_397),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_371),
.A2(n_352),
.B(n_356),
.Y(n_439)
);

OAI21x1_ASAP7_75t_L g440 ( 
.A1(n_433),
.A2(n_423),
.B(n_437),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_408),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_413),
.A2(n_429),
.B(n_422),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_407),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_404),
.A2(n_435),
.B(n_406),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_412),
.Y(n_446)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_407),
.Y(n_448)
);

AO31x2_ASAP7_75t_L g449 ( 
.A1(n_419),
.A2(n_421),
.A3(n_427),
.B(n_428),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_420),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_409),
.A2(n_416),
.B(n_439),
.Y(n_451)
);

AO21x2_ASAP7_75t_L g452 ( 
.A1(n_431),
.A2(n_432),
.B(n_418),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_434),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_417),
.A2(n_436),
.B1(n_410),
.B2(n_426),
.Y(n_454)
);

INVx4_ASAP7_75t_SL g455 ( 
.A(n_425),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_415),
.B(n_430),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_411),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_436),
.A2(n_405),
.B(n_430),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_430),
.A2(n_438),
.B(n_405),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_438),
.A2(n_433),
.B(n_423),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_438),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_406),
.B(n_296),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_426),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_425),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_433),
.A2(n_423),
.B(n_437),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_446),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_450),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_463),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_453),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_455),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_463),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_459),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_458),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_458),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_447),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_447),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_443),
.B(n_448),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_443),
.Y(n_484)
);

INVx5_ASAP7_75t_SL g485 ( 
.A(n_443),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_454),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_441),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_481),
.Y(n_489)
);

BUFx12f_ASAP7_75t_L g490 ( 
.A(n_467),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_468),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_471),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_467),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_448),
.Y(n_494)
);

OAI22xp33_ASAP7_75t_L g495 ( 
.A1(n_469),
.A2(n_444),
.B1(n_461),
.B2(n_457),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_448),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_466),
.B(n_464),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_473),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_466),
.B(n_461),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_464),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

AOI31xp33_ASAP7_75t_L g504 ( 
.A1(n_469),
.A2(n_488),
.A3(n_454),
.B(n_479),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_485),
.B(n_449),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_481),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_449),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_449),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_449),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_482),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_484),
.B(n_452),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_480),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_487),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_475),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_442),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_452),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_451),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_491),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_486),
.Y(n_519)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_478),
.C(n_470),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_493),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_499),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_476),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_512),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_476),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_500),
.B(n_472),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_497),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_497),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_502),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_498),
.B(n_480),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_460),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_494),
.B(n_477),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_509),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_490),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_490),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_440),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_514),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_518),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_533),
.B(n_509),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_522),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_521),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_495),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_527),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_524),
.B(n_495),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_528),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_519),
.B(n_523),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_524),
.B(n_513),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_526),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_519),
.B(n_517),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_525),
.B(n_514),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_534),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_509),
.Y(n_552)
);

OAI32xp33_ASAP7_75t_L g553 ( 
.A1(n_544),
.A2(n_520),
.A3(n_547),
.B1(n_542),
.B2(n_541),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_543),
.B(n_523),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_538),
.Y(n_555)
);

OAI22xp33_ASAP7_75t_L g556 ( 
.A1(n_541),
.A2(n_532),
.B1(n_535),
.B2(n_534),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_R g557 ( 
.A(n_549),
.B(n_536),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_546),
.B(n_536),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_540),
.B(n_526),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_552),
.B(n_525),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_539),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_558),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_554),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_555),
.B(n_545),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_554),
.B(n_539),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_559),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_553),
.A2(n_440),
.B(n_465),
.Y(n_567)
);

OAI321xp33_ASAP7_75t_L g568 ( 
.A1(n_564),
.A2(n_556),
.A3(n_551),
.B1(n_550),
.B2(n_548),
.C(n_535),
.Y(n_568)
);

AOI221xp5_ASAP7_75t_L g569 ( 
.A1(n_566),
.A2(n_550),
.B1(n_510),
.B2(n_501),
.C(n_537),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_567),
.A2(n_511),
.B(n_515),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_564),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_563),
.Y(n_572)
);

NAND4xp25_ASAP7_75t_L g573 ( 
.A(n_570),
.B(n_567),
.C(n_557),
.D(n_565),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_SL g574 ( 
.A(n_569),
.B(n_561),
.C(n_516),
.Y(n_574)
);

AO21x1_ASAP7_75t_L g575 ( 
.A1(n_571),
.A2(n_529),
.B(n_531),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_568),
.A2(n_572),
.B(n_562),
.Y(n_576)
);

NAND4xp25_ASAP7_75t_L g577 ( 
.A(n_570),
.B(n_501),
.C(n_496),
.D(n_494),
.Y(n_577)
);

AOI211xp5_ASAP7_75t_L g578 ( 
.A1(n_573),
.A2(n_501),
.B(n_496),
.C(n_494),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_574),
.B(n_576),
.Y(n_579)
);

AOI211x1_ASAP7_75t_SL g580 ( 
.A1(n_577),
.A2(n_506),
.B(n_489),
.C(n_492),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_579),
.B(n_575),
.Y(n_581)
);

NOR3xp33_ASAP7_75t_L g582 ( 
.A(n_578),
.B(n_503),
.C(n_496),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_581),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_583),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_584),
.A2(n_582),
.B(n_580),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_585),
.A2(n_506),
.B1(n_489),
.B2(n_503),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_586),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_587),
.A2(n_477),
.B(n_503),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_588),
.B(n_506),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_589),
.B(n_531),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_590),
.A2(n_506),
.B1(n_489),
.B2(n_481),
.Y(n_591)
);


endmodule