module fake_jpeg_531_n_216 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_45),
.Y(n_59)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_1),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_79),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_49),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_64),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_94),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_60),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_97),
.Y(n_134)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_80),
.B1(n_76),
.B2(n_58),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_109),
.B1(n_110),
.B2(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_95),
.A2(n_73),
.B1(n_69),
.B2(n_65),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_108),
.Y(n_127)
);

INVx2_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_107),
.B(n_54),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_69),
.B(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_61),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_80),
.B1(n_76),
.B2(n_73),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_74),
.B1(n_71),
.B2(n_53),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_66),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_114),
.B(n_52),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_126),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_109),
.B1(n_98),
.B2(n_105),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_120),
.B1(n_129),
.B2(n_115),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_67),
.B(n_72),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_0),
.B(n_2),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_96),
.B1(n_71),
.B2(n_66),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_125),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_0),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_54),
.B1(n_62),
.B2(n_56),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_63),
.B1(n_47),
.B2(n_41),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_28),
.B(n_22),
.C(n_40),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_24),
.B(n_21),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_139),
.B1(n_143),
.B2(n_5),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_127),
.B1(n_134),
.B2(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_146),
.Y(n_170)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_141),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_51),
.B(n_59),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_144),
.A2(n_5),
.B(n_6),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_150),
.Y(n_161)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_39),
.C(n_33),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_160),
.C(n_151),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_160),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_167)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_4),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_158),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_10),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_164),
.B(n_176),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_12),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_27),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_178),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_181),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_8),
.B(n_9),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_162),
.B(n_172),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_143),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_10),
.C(n_12),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_13),
.C(n_14),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_149),
.B(n_19),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_153),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_152),
.B(n_141),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_183),
.A2(n_187),
.B(n_173),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_148),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_193),
.C(n_180),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_167),
.B1(n_164),
.B2(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_189),
.B(n_185),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_176),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_198),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_192),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_200),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_166),
.B1(n_169),
.B2(n_177),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_190),
.B(n_174),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_201),
.C(n_192),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_205),
.Y(n_209)
);

OAI21x1_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_196),
.B(n_194),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_194),
.Y(n_205)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_203),
.B(n_209),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_186),
.B1(n_188),
.B2(n_199),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_19),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_210),
.A2(n_211),
.B1(n_13),
.B2(n_14),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_15),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_213),
.A2(n_15),
.B(n_16),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_17),
.C(n_18),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_215),
.B(n_17),
.Y(n_216)
);


endmodule