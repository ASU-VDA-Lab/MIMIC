module fake_jpeg_25928_n_63 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_3),
.B(n_4),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_37),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_39),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_1),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_19),
.A2(n_23),
.B1(n_31),
.B2(n_26),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_22),
.C(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_32),
.B1(n_36),
.B2(n_33),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.C(n_30),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_42),
.C(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_48),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_27),
.B1(n_30),
.B2(n_22),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_44),
.B(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_56),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_53),
.C(n_35),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_25),
.C(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_24),
.B2(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_34),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_2),
.C(n_4),
.Y(n_63)
);


endmodule