module fake_netlist_6_1541_n_418 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_108, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_103, n_111, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_418);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_108;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_418;

wire n_326;
wire n_256;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_141;
wire n_383;
wire n_200;
wire n_176;
wire n_114;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_344;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_397;
wire n_155;
wire n_122;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_417;
wire n_374;
wire n_366;
wire n_407;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_406;
wire n_204;
wire n_261;
wire n_312;
wire n_394;
wire n_130;
wire n_164;
wire n_292;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_317;
wire n_149;
wire n_347;
wire n_328;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_391;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_43),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_16),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_56),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_30),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_39),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_38),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_24),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_51),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_19),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_27),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_37),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_50),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_44),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx8_ASAP7_75t_SL g142 ( 
.A(n_32),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g144 ( 
.A(n_33),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_47),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_46),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_108),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_59),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_45),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_55),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_48),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_25),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_4),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_9),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_81),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_20),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_67),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_90),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_28),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_14),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_26),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_12),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_15),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_36),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_4),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_0),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_2),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_3),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_49),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_54),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_31),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

BUFx8_ASAP7_75t_SL g186 ( 
.A(n_142),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

BUFx8_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_124),
.B(n_2),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

AND2x4_ASAP7_75t_L g198 ( 
.A(n_125),
.B(n_5),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

OAI22x1_ASAP7_75t_R g200 ( 
.A1(n_133),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_163),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_119),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_141),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

INVxp33_ASAP7_75t_SL g211 ( 
.A(n_148),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_114),
.Y(n_215)
);

OAI22x1_ASAP7_75t_R g216 ( 
.A1(n_159),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_216)
);

AND2x4_ASAP7_75t_SL g217 ( 
.A(n_152),
.B(n_29),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

BUFx8_ASAP7_75t_SL g219 ( 
.A(n_153),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_113),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_147),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_156),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_116),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_117),
.Y(n_226)
);

BUFx8_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_118),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_123),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_130),
.Y(n_230)
);

CKINVDCx11_ASAP7_75t_R g231 ( 
.A(n_162),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_134),
.B(n_21),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_137),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_139),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_174),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_121),
.B(n_22),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_186),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_207),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_219),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_231),
.Y(n_248)
);

NAND2xp33_ASAP7_75t_R g249 ( 
.A(n_211),
.B(n_180),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_215),
.Y(n_250)
);

BUFx2_ASAP7_75t_SL g251 ( 
.A(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_226),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_188),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_187),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_202),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_227),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_201),
.A2(n_128),
.B1(n_167),
.B2(n_166),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_189),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_237),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_157),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_239),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_158),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_240),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_238),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_191),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_238),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_212),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_217),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_190),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

OR2x6_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_204),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_242),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_222),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_277),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_222),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_250),
.B(n_254),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_260),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_194),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_221),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_194),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_198),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_194),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_206),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_251),
.B(n_206),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_262),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_171),
.C(n_112),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_233),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_284),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_264),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_200),
.B1(n_216),
.B2(n_248),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_290),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_193),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_R g318 ( 
.A(n_298),
.B(n_245),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_160),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_291),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_297),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_278),
.B(n_165),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_297),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_288),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_181),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_182),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_307),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_285),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_306),
.B(n_122),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_300),
.A2(n_225),
.B1(n_235),
.B2(n_224),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_246),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_318),
.Y(n_335)
);

OR2x6_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_205),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_129),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g338 ( 
.A1(n_331),
.A2(n_295),
.B(n_287),
.C(n_195),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_312),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_322),
.A2(n_214),
.B(n_209),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_261),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_321),
.A2(n_218),
.B(n_214),
.Y(n_343)
);

AOI21x1_ASAP7_75t_L g344 ( 
.A1(n_328),
.A2(n_301),
.B(n_299),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_323),
.A2(n_218),
.B(n_196),
.Y(n_345)
);

A2O1A1Ixp33_ASAP7_75t_L g346 ( 
.A1(n_319),
.A2(n_136),
.B(n_138),
.C(n_135),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_140),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_145),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_324),
.B(n_146),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_150),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_324),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_320),
.B(n_151),
.Y(n_352)
);

A2O1A1Ixp33_ASAP7_75t_SL g353 ( 
.A1(n_311),
.A2(n_327),
.B(n_329),
.C(n_326),
.Y(n_353)
);

AO21x2_ASAP7_75t_L g354 ( 
.A1(n_338),
.A2(n_332),
.B(n_333),
.Y(n_354)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_340),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g357 ( 
.A1(n_344),
.A2(n_197),
.B(n_203),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_325),
.Y(n_358)
);

OR2x6_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_313),
.Y(n_359)
);

OR2x4_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_234),
.Y(n_360)
);

NOR2x1_ASAP7_75t_R g361 ( 
.A(n_335),
.B(n_352),
.Y(n_361)
);

AO21x2_ASAP7_75t_L g362 ( 
.A1(n_353),
.A2(n_236),
.B(n_234),
.Y(n_362)
);

AO21x2_ASAP7_75t_L g363 ( 
.A1(n_346),
.A2(n_236),
.B(n_234),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_348),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_350),
.Y(n_365)
);

NAND2x1p5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_208),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_347),
.A2(n_345),
.B(n_343),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_356),
.Y(n_369)
);

NAND2x1p5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_342),
.Y(n_370)
);

AOI21x1_ASAP7_75t_L g371 ( 
.A1(n_357),
.A2(n_341),
.B(n_241),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_364),
.A2(n_175),
.B1(n_184),
.B2(n_183),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g373 ( 
.A1(n_364),
.A2(n_360),
.B1(n_358),
.B2(n_367),
.Y(n_373)
);

NAND2x1p5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_208),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_L g375 ( 
.A1(n_360),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_365),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_369),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_359),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_354),
.Y(n_379)
);

AO21x2_ASAP7_75t_L g380 ( 
.A1(n_371),
.A2(n_362),
.B(n_363),
.Y(n_380)
);

NOR3xp33_ASAP7_75t_SL g381 ( 
.A(n_375),
.B(n_361),
.C(n_366),
.Y(n_381)
);

OR2x6_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_368),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_374),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_377),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_382),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_376),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_382),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_382),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_380),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_381),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_385),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_387),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_383),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_390),
.B(n_388),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_385),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_391),
.B(n_389),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_394),
.B(n_393),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_395),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_398),
.Y(n_399)
);

AND2x4_ASAP7_75t_SL g400 ( 
.A(n_399),
.B(n_397),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_400),
.B(n_396),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_401),
.Y(n_402)
);

OAI221xp5_ASAP7_75t_L g403 ( 
.A1(n_402),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.C(n_65),
.Y(n_403)
);

NOR2x1_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_71),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_404),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_405),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_407),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_409),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_408),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_410),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_411),
.A2(n_85),
.B(n_86),
.Y(n_413)
);

AOI31xp33_ASAP7_75t_L g414 ( 
.A1(n_412),
.A2(n_87),
.A3(n_88),
.B(n_89),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_413),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_415),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_416)
);

OR2x6_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_414),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_417),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_418)
);


endmodule