module real_aes_7655_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_623;
wire n_249;
wire n_446;
wire n_221;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_0), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_1), .Y(n_604) );
XOR2x2_ASAP7_75t_L g541 ( .A(n_2), .B(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_3), .A2(n_13), .B1(n_379), .B2(n_614), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_4), .A2(n_48), .B1(n_325), .B2(n_437), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_5), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_6), .A2(n_183), .B1(n_303), .B2(n_412), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_7), .Y(n_419) );
AOI222xp33_ASAP7_75t_L g554 ( .A1(n_8), .A2(n_24), .B1(n_172), .B2(n_537), .C1(n_555), .C2(n_556), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_9), .A2(n_595), .B1(n_622), .B2(n_623), .Y(n_594) );
INVx1_ASAP7_75t_L g622 ( .A(n_9), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_10), .A2(n_136), .B1(n_343), .B2(n_344), .Y(n_342) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_11), .A2(n_84), .B1(n_276), .B2(n_412), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_12), .A2(n_60), .B1(n_337), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_14), .A2(n_51), .B1(n_477), .B2(n_478), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_15), .A2(n_174), .B1(n_663), .B2(n_664), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_16), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_17), .A2(n_204), .B1(n_322), .B2(n_440), .Y(n_470) );
INVx1_ASAP7_75t_L g443 ( .A(n_18), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_19), .A2(n_62), .B1(n_223), .B2(n_507), .Y(n_506) );
AO22x2_ASAP7_75t_L g236 ( .A1(n_20), .A2(n_68), .B1(n_228), .B2(n_233), .Y(n_236) );
INVx1_ASAP7_75t_L g638 ( .A(n_20), .Y(n_638) );
XOR2xp5_ASAP7_75t_L g641 ( .A(n_21), .B(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_22), .A2(n_123), .B1(n_335), .B2(n_407), .Y(n_406) );
AOI222xp33_ASAP7_75t_L g535 ( .A1(n_23), .A2(n_83), .B1(n_104), .B2(n_460), .C1(n_536), .C2(n_537), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_25), .A2(n_27), .B1(n_347), .B2(n_614), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_26), .A2(n_179), .B1(n_360), .B2(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g291 ( .A(n_28), .Y(n_291) );
AOI222xp33_ASAP7_75t_L g416 ( .A1(n_29), .A2(n_74), .B1(n_189), .B2(n_275), .C1(n_417), .C2(n_418), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_30), .A2(n_145), .B1(n_418), .B2(n_445), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_31), .A2(n_52), .B1(n_322), .B2(n_653), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_32), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_33), .A2(n_41), .B1(n_429), .B2(n_430), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_34), .A2(n_35), .B1(n_325), .B2(n_327), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_36), .A2(n_162), .B1(n_300), .B2(n_344), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_37), .Y(n_377) );
AO22x2_ASAP7_75t_L g238 ( .A1(n_38), .A2(n_70), .B1(n_228), .B2(n_229), .Y(n_238) );
INVx1_ASAP7_75t_L g639 ( .A(n_38), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_39), .A2(n_127), .B1(n_286), .B2(n_507), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g329 ( .A1(n_40), .A2(n_168), .B1(n_272), .B2(n_330), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_42), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_43), .A2(n_119), .B1(n_477), .B2(n_478), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_44), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g515 ( .A(n_45), .Y(n_515) );
AOI22xp5_ASAP7_75t_SL g424 ( .A1(n_46), .A2(n_195), .B1(n_367), .B2(n_425), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_47), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_49), .A2(n_99), .B1(n_619), .B2(n_620), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_50), .A2(n_164), .B1(n_509), .B2(n_568), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_53), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_54), .A2(n_190), .B1(n_440), .B2(n_441), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_55), .A2(n_161), .B1(n_343), .B2(n_509), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_56), .A2(n_75), .B1(n_512), .B2(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_57), .B(n_437), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_58), .A2(n_128), .B1(n_373), .B2(n_475), .Y(n_534) );
INVx1_ASAP7_75t_L g591 ( .A(n_59), .Y(n_591) );
AOI22xp33_ASAP7_75t_SL g320 ( .A1(n_61), .A2(n_122), .B1(n_321), .B2(n_322), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_63), .A2(n_126), .B1(n_298), .B2(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_64), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_65), .A2(n_97), .B1(n_241), .B2(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_66), .A2(n_194), .B1(n_264), .B2(n_384), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_67), .A2(n_201), .B1(n_328), .B2(n_383), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_69), .A2(n_118), .B1(n_253), .B2(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g333 ( .A1(n_71), .A2(n_166), .B1(n_334), .B2(n_335), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_72), .A2(n_197), .B1(n_241), .B2(n_339), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_73), .A2(n_160), .B1(n_433), .B2(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g214 ( .A(n_76), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_77), .A2(n_105), .B1(n_293), .B2(n_533), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_78), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_79), .A2(n_147), .B1(n_347), .B2(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_80), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g211 ( .A(n_81), .Y(n_211) );
INVx1_ASAP7_75t_L g446 ( .A(n_82), .Y(n_446) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_85), .A2(n_208), .B(n_216), .C(n_640), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_86), .Y(n_365) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_87), .A2(n_200), .B1(n_293), .B2(n_348), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_88), .A2(n_181), .B1(n_253), .B2(n_344), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_89), .A2(n_137), .B1(n_295), .B2(n_343), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_90), .A2(n_100), .B1(n_344), .B2(n_348), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_91), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_92), .Y(n_490) );
INVx1_ASAP7_75t_L g296 ( .A(n_93), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_94), .B(n_307), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_95), .A2(n_132), .B1(n_303), .B2(n_418), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g394 ( .A1(n_96), .A2(n_109), .B1(n_169), .B2(n_395), .C1(n_398), .C2(n_399), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_98), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_101), .A2(n_106), .B1(n_303), .B2(n_412), .Y(n_545) );
INVx1_ASAP7_75t_L g281 ( .A(n_102), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_103), .Y(n_579) );
AO22x2_ASAP7_75t_L g351 ( .A1(n_107), .A2(n_352), .B1(n_400), .B2(n_401), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_107), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_108), .A2(n_202), .B1(n_334), .B2(n_347), .Y(n_552) );
INVx1_ASAP7_75t_L g289 ( .A(n_110), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_111), .A2(n_113), .B1(n_223), .B2(n_239), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_112), .A2(n_188), .B1(n_367), .B2(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_114), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g301 ( .A1(n_115), .A2(n_143), .B1(n_149), .B2(n_302), .C1(n_303), .C2(n_307), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_116), .B(n_398), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_117), .A2(n_206), .B1(n_382), .B2(n_384), .C(n_385), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_120), .A2(n_148), .B1(n_434), .B2(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g215 ( .A(n_121), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_124), .A2(n_191), .B1(n_525), .B2(n_526), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_125), .Y(n_600) );
AND2x6_ASAP7_75t_L g210 ( .A(n_129), .B(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_129), .Y(n_632) );
AO22x2_ASAP7_75t_L g227 ( .A1(n_130), .A2(n_178), .B1(n_228), .B2(n_229), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_131), .A2(n_198), .B1(n_245), .B2(n_252), .Y(n_244) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_133), .A2(n_155), .B1(n_307), .B2(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g349 ( .A(n_134), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_135), .A2(n_177), .B1(n_360), .B2(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_138), .B(n_383), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_139), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_140), .A2(n_192), .B1(n_429), .B2(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_141), .Y(n_590) );
INVx1_ASAP7_75t_L g258 ( .A(n_142), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_144), .Y(n_539) );
INVx1_ASAP7_75t_L g310 ( .A(n_146), .Y(n_310) );
AOI22xp33_ASAP7_75t_SL g336 ( .A1(n_150), .A2(n_171), .B1(n_337), .B2(n_339), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_151), .B(n_327), .Y(n_326) );
AO22x2_ASAP7_75t_L g232 ( .A1(n_152), .A2(n_184), .B1(n_228), .B2(n_233), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_153), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_154), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_156), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_157), .A2(n_187), .B1(n_270), .B2(n_275), .Y(n_269) );
INVx1_ASAP7_75t_L g503 ( .A(n_158), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_159), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_163), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_165), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_167), .B(n_263), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_170), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_173), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_175), .Y(n_589) );
XOR2x2_ASAP7_75t_L g455 ( .A(n_176), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_178), .B(n_637), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_180), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_182), .Y(n_386) );
INVx1_ASAP7_75t_L g635 ( .A(n_184), .Y(n_635) );
INVx1_ASAP7_75t_L g461 ( .A(n_185), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_186), .Y(n_674) );
OA22x2_ASAP7_75t_L g675 ( .A1(n_186), .A2(n_642), .B1(n_643), .B2(n_674), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_193), .Y(n_648) );
INVx1_ASAP7_75t_L g228 ( .A(n_196), .Y(n_228) );
INVx1_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g598 ( .A(n_199), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_203), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_205), .Y(n_494) );
INVx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_210), .B(n_212), .Y(n_209) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_211), .Y(n_631) );
OA21x2_ASAP7_75t_L g672 ( .A1(n_212), .A2(n_630), .B(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_215), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_451), .B1(n_625), .B2(n_626), .C(n_627), .Y(n_216) );
INVx1_ASAP7_75t_L g625 ( .A(n_217), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_311), .B1(n_449), .B2(n_450), .Y(n_217) );
INVx1_ASAP7_75t_SL g449 ( .A(n_218), .Y(n_449) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
XOR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_310), .Y(n_219) );
NAND4xp75_ASAP7_75t_L g220 ( .A(n_221), .B(n_257), .C(n_279), .D(n_301), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_244), .Y(n_221) );
BUFx2_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_224), .Y(n_343) );
INVx2_ASAP7_75t_L g356 ( .A(n_224), .Y(n_356) );
BUFx2_ASAP7_75t_SL g533 ( .A(n_224), .Y(n_533) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_234), .Y(n_224) );
AND2x6_ASAP7_75t_L g295 ( .A(n_225), .B(n_267), .Y(n_295) );
AND2x4_ASAP7_75t_L g300 ( .A(n_225), .B(n_251), .Y(n_300) );
AND2x6_ASAP7_75t_L g302 ( .A(n_225), .B(n_278), .Y(n_302) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_231), .Y(n_225) );
AND2x2_ASAP7_75t_L g243 ( .A(n_226), .B(n_232), .Y(n_243) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g249 ( .A(n_227), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_227), .B(n_232), .Y(n_256) );
AND2x2_ASAP7_75t_L g274 ( .A(n_227), .B(n_236), .Y(n_274) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g233 ( .A(n_230), .Y(n_233) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g250 ( .A(n_232), .Y(n_250) );
INVx1_ASAP7_75t_L g306 ( .A(n_232), .Y(n_306) );
AND2x4_ASAP7_75t_L g242 ( .A(n_234), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_234), .B(n_249), .Y(n_284) );
AND2x4_ASAP7_75t_L g287 ( .A(n_234), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g345 ( .A(n_234), .B(n_249), .Y(n_345) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
AND2x2_ASAP7_75t_L g251 ( .A(n_235), .B(n_238), .Y(n_251) );
OR2x2_ASAP7_75t_L g268 ( .A(n_235), .B(n_238), .Y(n_268) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g278 ( .A(n_236), .B(n_238), .Y(n_278) );
AND2x2_ASAP7_75t_L g305 ( .A(n_237), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g340 ( .A(n_237), .Y(n_340) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g255 ( .A(n_238), .Y(n_255) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx4_ASAP7_75t_L g433 ( .A(n_240), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_240), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_572) );
INVx4_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g338 ( .A(n_242), .Y(n_338) );
BUFx3_ASAP7_75t_L g360 ( .A(n_242), .Y(n_360) );
BUFx3_ASAP7_75t_L g620 ( .A(n_242), .Y(n_620) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_243), .B(n_251), .Y(n_261) );
AND2x4_ASAP7_75t_L g266 ( .A(n_243), .B(n_267), .Y(n_266) );
AND2x6_ASAP7_75t_L g328 ( .A(n_243), .B(n_251), .Y(n_328) );
INVx1_ASAP7_75t_L g493 ( .A(n_243), .Y(n_493) );
INVx3_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx5_ASAP7_75t_L g335 ( .A(n_247), .Y(n_335) );
INVx4_ASAP7_75t_L g426 ( .A(n_247), .Y(n_426) );
INVx2_ASAP7_75t_L g509 ( .A(n_247), .Y(n_509) );
INVx3_ASAP7_75t_L g525 ( .A(n_247), .Y(n_525) );
INVx1_ASAP7_75t_L g659 ( .A(n_247), .Y(n_659) );
INVx8_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_249), .B(n_251), .Y(n_364) );
INVx1_ASAP7_75t_L g277 ( .A(n_250), .Y(n_277) );
BUFx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
BUFx2_ASAP7_75t_L g367 ( .A(n_253), .Y(n_367) );
BUFx2_ASAP7_75t_L g478 ( .A(n_253), .Y(n_478) );
BUFx2_ASAP7_75t_L g526 ( .A(n_253), .Y(n_526) );
INVx6_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g568 ( .A(n_254), .Y(n_568) );
OR2x6_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g273 ( .A(n_255), .Y(n_273) );
INVx1_ASAP7_75t_L g288 ( .A(n_256), .Y(n_288) );
OA211x2_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B(n_262), .C(n_269), .Y(n_257) );
OA211x2_ASAP7_75t_L g527 ( .A1(n_259), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
BUFx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g496 ( .A(n_261), .Y(n_496) );
BUFx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g325 ( .A(n_265), .Y(n_325) );
INVx5_ASAP7_75t_L g383 ( .A(n_265), .Y(n_383) );
INVx2_ASAP7_75t_L g469 ( .A(n_265), .Y(n_469) );
INVx4_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g492 ( .A(n_268), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
BUFx3_ASAP7_75t_L g412 ( .A(n_272), .Y(n_412) );
BUFx2_ASAP7_75t_L g440 ( .A(n_272), .Y(n_440) );
BUFx2_ASAP7_75t_L g653 ( .A(n_272), .Y(n_653) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AND2x4_ASAP7_75t_L g304 ( .A(n_274), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g308 ( .A(n_274), .B(n_309), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_274), .B(n_340), .Y(n_388) );
BUFx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx2_ASAP7_75t_SL g322 ( .A(n_276), .Y(n_322) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_276), .Y(n_441) );
BUFx2_ASAP7_75t_SL g556 ( .A(n_276), .Y(n_556) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g393 ( .A(n_277), .Y(n_393) );
INVx1_ASAP7_75t_L g392 ( .A(n_278), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_290), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_285), .B2(n_289), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_282), .A2(n_297), .B1(n_570), .B2(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g376 ( .A(n_283), .Y(n_376) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx3_ASAP7_75t_L g348 ( .A(n_287), .Y(n_348) );
BUFx3_ASAP7_75t_L g380 ( .A(n_287), .Y(n_380) );
BUFx2_ASAP7_75t_SL g434 ( .A(n_287), .Y(n_434) );
BUFx2_ASAP7_75t_L g514 ( .A(n_287), .Y(n_514) );
INVx1_ASAP7_75t_L g550 ( .A(n_287), .Y(n_550) );
BUFx2_ASAP7_75t_SL g576 ( .A(n_287), .Y(n_576) );
AND2x2_ASAP7_75t_L g339 ( .A(n_288), .B(n_340), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B1(n_296), .B2(n_297), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx4_ASAP7_75t_L g334 ( .A(n_294), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_294), .A2(n_370), .B1(n_371), .B2(n_372), .Y(n_369) );
INVx11_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx11_ASAP7_75t_L g431 ( .A(n_295), .Y(n_431) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g484 ( .A(n_299), .Y(n_484) );
INVx2_ASAP7_75t_L g616 ( .A(n_299), .Y(n_616) );
INVx6_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx3_ASAP7_75t_L g347 ( .A(n_300), .Y(n_347) );
BUFx3_ASAP7_75t_L g373 ( .A(n_300), .Y(n_373) );
BUFx3_ASAP7_75t_L g407 ( .A(n_300), .Y(n_407) );
INVx2_ASAP7_75t_L g318 ( .A(n_302), .Y(n_318) );
INVx4_ASAP7_75t_L g397 ( .A(n_302), .Y(n_397) );
BUFx3_ASAP7_75t_L g417 ( .A(n_302), .Y(n_417) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_302), .Y(n_555) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_303), .Y(n_536) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx4f_ASAP7_75t_SL g330 ( .A(n_304), .Y(n_330) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_304), .Y(n_398) );
BUFx2_ASAP7_75t_L g445 ( .A(n_304), .Y(n_445) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_304), .Y(n_465) );
INVx1_ASAP7_75t_L g309 ( .A(n_306), .Y(n_309) );
INVx1_ASAP7_75t_L g649 ( .A(n_307), .Y(n_649) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_308), .Y(n_321) );
BUFx12f_ASAP7_75t_L g418 ( .A(n_308), .Y(n_418) );
INVx1_ASAP7_75t_L g450 ( .A(n_311), .Y(n_450) );
XOR2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_350), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
XOR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_349), .Y(n_314) );
NAND2x1_ASAP7_75t_L g315 ( .A(n_316), .B(n_331), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_323), .Y(n_316) );
OAI21xp5_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_319), .B(n_320), .Y(n_317) );
BUFx3_ASAP7_75t_L g399 ( .A(n_321), .Y(n_399) );
INVx2_ASAP7_75t_L g585 ( .A(n_321), .Y(n_585) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .C(n_329), .Y(n_323) );
BUFx4f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g384 ( .A(n_328), .Y(n_384) );
INVx1_ASAP7_75t_SL g438 ( .A(n_328), .Y(n_438) );
INVx1_ASAP7_75t_L g647 ( .A(n_330), .Y(n_647) );
NOR2x1_ASAP7_75t_L g331 ( .A(n_332), .B(n_341), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_336), .Y(n_332) );
BUFx2_ASAP7_75t_L g477 ( .A(n_335), .Y(n_477) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_346), .Y(n_341) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_343), .Y(n_429) );
BUFx3_ASAP7_75t_L g619 ( .A(n_343), .Y(n_619) );
BUFx3_ASAP7_75t_L g663 ( .A(n_343), .Y(n_663) );
INVx1_ASAP7_75t_L g482 ( .A(n_344), .Y(n_482) );
BUFx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g507 ( .A(n_345), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_402), .B1(n_447), .B2(n_448), .Y(n_350) );
INVx1_ASAP7_75t_L g447 ( .A(n_351), .Y(n_447) );
INVx1_ASAP7_75t_L g401 ( .A(n_352), .Y(n_401) );
AND4x1_ASAP7_75t_L g352 ( .A(n_353), .B(n_368), .C(n_381), .D(n_394), .Y(n_352) );
NOR2xp33_ASAP7_75t_SL g353 ( .A(n_354), .B(n_361), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_357), .B2(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B1(n_365), .B2(n_366), .Y(n_361) );
BUFx2_ASAP7_75t_R g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_SL g368 ( .A(n_369), .B(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_377), .B2(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_389), .B2(n_390), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_387), .A2(n_391), .B1(n_502), .B2(n_503), .Y(n_501) );
BUFx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx4_ASAP7_75t_L g581 ( .A(n_388), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_388), .A2(n_390), .B1(n_609), .B2(n_610), .Y(n_608) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_391), .A2(n_579), .B1(n_580), .B2(n_582), .Y(n_578) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI21xp5_ASAP7_75t_SL g442 ( .A1(n_396), .A2(n_443), .B(n_444), .Y(n_442) );
BUFx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx4_ASAP7_75t_L g460 ( .A(n_397), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g583 ( .A1(n_397), .A2(n_584), .B1(n_585), .B2(n_586), .C(n_587), .Y(n_583) );
INVx1_ASAP7_75t_L g448 ( .A(n_402), .Y(n_448) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_420), .Y(n_402) );
XOR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_419), .Y(n_403) );
NAND4xp75_ASAP7_75t_L g404 ( .A(n_405), .B(n_409), .C(n_413), .D(n_416), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
AND2x2_ASAP7_75t_SL g409 ( .A(n_410), .B(n_411), .Y(n_409) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx3_ASAP7_75t_L g499 ( .A(n_417), .Y(n_499) );
INVx2_ASAP7_75t_L g538 ( .A(n_418), .Y(n_538) );
XOR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_446), .Y(n_420) );
NOR4xp75_ASAP7_75t_L g421 ( .A(n_422), .B(n_427), .C(n_435), .D(n_442), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_423), .B(n_424), .Y(n_422) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2x1_ASAP7_75t_L g427 ( .A(n_428), .B(n_432), .Y(n_427) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g475 ( .A(n_431), .Y(n_475) );
INVx4_ASAP7_75t_L g512 ( .A(n_431), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_436), .B(n_439), .Y(n_435) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g626 ( .A(n_451), .Y(n_626) );
AOI22xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_558), .B1(n_559), .B2(n_624), .Y(n_451) );
INVx1_ASAP7_75t_L g624 ( .A(n_452), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_517), .B2(n_518), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_485), .B1(n_486), .B2(n_516), .Y(n_454) );
INVx2_ASAP7_75t_L g516 ( .A(n_455), .Y(n_516) );
NAND3x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_471), .C(n_479), .Y(n_456) );
NOR2x1_ASAP7_75t_SL g457 ( .A(n_458), .B(n_466), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_461), .B(n_462), .Y(n_458) );
OAI222xp33_ASAP7_75t_L g645 ( .A1(n_459), .A2(n_646), .B1(n_647), .B2(n_648), .C1(n_649), .C2(n_650), .Y(n_645) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx4_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .C(n_470), .Y(n_466) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
XOR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_515), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_504), .Y(n_487) );
NOR3xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_497), .C(n_501), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_494), .B2(n_495), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_491), .A2(n_495), .B1(n_589), .B2(n_590), .Y(n_588) );
BUFx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_492), .Y(n_599) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_SL g601 ( .A(n_496), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_500), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_510), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
BUFx3_ASAP7_75t_L g614 ( .A(n_507), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_520), .B1(n_540), .B2(n_557), .Y(n_518) );
INVx3_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
XOR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_539), .Y(n_520) );
NAND4xp75_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .C(n_531), .D(n_535), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
INVx2_ASAP7_75t_SL g605 ( .A(n_536), .Y(n_605) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g557 ( .A(n_541), .Y(n_557) );
NAND4xp75_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .C(n_551), .D(n_554), .Y(n_542) );
AND2x2_ASAP7_75t_SL g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_SL g603 ( .A(n_555), .Y(n_603) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B1(n_592), .B2(n_593), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
XOR2xp5_ASAP7_75t_SL g562 ( .A(n_563), .B(n_591), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_577), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_569), .C(n_572), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .C(n_588), .Y(n_577) );
INVx3_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g623 ( .A(n_595), .Y(n_623) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_611), .Y(n_595) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_602), .C(n_608), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_600), .B2(n_601), .Y(n_597) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_605), .B2(n_606), .C(n_607), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_617), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .Y(n_617) );
INVx1_ASAP7_75t_L g665 ( .A(n_620), .Y(n_665) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_629), .B(n_633), .Y(n_628) );
OR2x2_ASAP7_75t_SL g678 ( .A(n_629), .B(n_634), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_630), .Y(n_667) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_631), .B(n_671), .Y(n_673) );
CKINVDCx16_ASAP7_75t_R g671 ( .A(n_632), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OAI322xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_666), .A3(n_668), .B1(n_672), .B2(n_674), .C1(n_675), .C2(n_676), .Y(n_640) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND3x1_ASAP7_75t_L g643 ( .A(n_644), .B(n_655), .C(n_660), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_651), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_677), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
endmodule