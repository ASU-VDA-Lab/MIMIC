module fake_ariane_2673_n_1957 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1957);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1957;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g201 ( 
.A(n_20),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_112),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_106),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_190),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_43),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_50),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_25),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_22),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_1),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_94),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_86),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_172),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_39),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_137),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_156),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_82),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_120),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_27),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_87),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_29),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_45),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_58),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_76),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_169),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_194),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_108),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_27),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_49),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_114),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_4),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_21),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_93),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_70),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_0),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_38),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_79),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_53),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_25),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_61),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_121),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_142),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_153),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_149),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_80),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_92),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_146),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_148),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_188),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_36),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_90),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_130),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_199),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_64),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_173),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_98),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_99),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_126),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_124),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_67),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_21),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_127),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_26),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_7),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_166),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_50),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_41),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_44),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_140),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_70),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_64),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_128),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_182),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_83),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_35),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_3),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_7),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_45),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_56),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_41),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_167),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_200),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_192),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_110),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_102),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_129),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_154),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_113),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_133),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_81),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_180),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_139),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_59),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_179),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_183),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_109),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_138),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_20),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_66),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_103),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_165),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_13),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_69),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_54),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_28),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_52),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_174),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_175),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_187),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_52),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_135),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_68),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_59),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_123),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_168),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_160),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_10),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_161),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_176),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_51),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_18),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_47),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_97),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_60),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_91),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_189),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_85),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_23),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_144),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_15),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_32),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_186),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_24),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_67),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_162),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_197),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_36),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_5),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_63),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_115),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_185),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_35),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_51),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_159),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_16),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_117),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_151),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_23),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_0),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_96),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_2),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_34),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_47),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_141),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_32),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_56),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_6),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_40),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_107),
.Y(n_369)
);

BUFx10_ASAP7_75t_L g370 ( 
.A(n_19),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_136),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_15),
.Y(n_372)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_10),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_122),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_42),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_195),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_30),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_198),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_31),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_60),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_28),
.Y(n_381)
);

BUFx10_ASAP7_75t_L g382 ( 
.A(n_4),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_145),
.Y(n_383)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_2),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_101),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_66),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_132),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_54),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_191),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_31),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_14),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_177),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_163),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_74),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_143),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_77),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_58),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_43),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_116),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_218),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_368),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_223),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_268),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_291),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_311),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_396),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_240),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_248),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_238),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_277),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_260),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_373),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_250),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_278),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_251),
.B(n_1),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_241),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_373),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_271),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_219),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_273),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_207),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_276),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_384),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_289),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_207),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_384),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_235),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_241),
.B(n_3),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_384),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_370),
.B(n_5),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_384),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_280),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_314),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_286),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_206),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_287),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_365),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_375),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_R g450 ( 
.A(n_318),
.B(n_105),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_339),
.B(n_6),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_384),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_285),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_288),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_377),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_285),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_201),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_208),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_290),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_390),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_309),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_312),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_315),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_210),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_235),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_316),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_233),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_211),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_208),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_242),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_395),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_226),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_320),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_215),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_356),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_229),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_345),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_215),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_272),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_272),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_319),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_319),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_331),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_247),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_264),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_322),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_327),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_356),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_274),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_334),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_356),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_281),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_249),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_340),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_341),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_308),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_426),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_236),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_371),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_406),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_426),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_426),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_426),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_465),
.B(n_299),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_458),
.A2(n_204),
.B(n_203),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_407),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_371),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_305),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_416),
.B(n_424),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_412),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_417),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_417),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_421),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_423),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_416),
.B(n_371),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_445),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_400),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_436),
.B(n_494),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_402),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_439),
.B(n_378),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_434),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_427),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_436),
.B(n_305),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_431),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_424),
.B(n_378),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_431),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_439),
.B(n_249),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_435),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_435),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_438),
.Y(n_541)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_438),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_440),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_440),
.B(n_209),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_442),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_485),
.B(n_378),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_442),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_448),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_448),
.B(n_452),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

NOR2x1_ASAP7_75t_L g553 ( 
.A(n_458),
.B(n_335),
.Y(n_553)
);

NAND2x1p5_ASAP7_75t_L g554 ( 
.A(n_437),
.B(n_369),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_470),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_470),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_475),
.A2(n_216),
.B(n_213),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_475),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_479),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_479),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_L g561 ( 
.A(n_410),
.B(n_369),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_480),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_480),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_420),
.B(n_202),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_481),
.B(n_313),
.Y(n_565)
);

NAND2x1_ASAP7_75t_L g566 ( 
.A(n_481),
.B(n_219),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_482),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_482),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_483),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_483),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_453),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_456),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_456),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_485),
.Y(n_575)
);

CKINVDCx11_ASAP7_75t_R g576 ( 
.A(n_411),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_457),
.B(n_221),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_523),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_532),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_500),
.B(n_415),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_548),
.B(n_425),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_527),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_523),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_532),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_548),
.B(n_484),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_523),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_523),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_561),
.A2(n_531),
.B1(n_548),
.B2(n_512),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_524),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_524),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_500),
.B(n_428),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_500),
.B(n_468),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_522),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_524),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_564),
.B(n_430),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_524),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_542),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_533),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_533),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_533),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_561),
.A2(n_451),
.B1(n_450),
.B2(n_441),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_512),
.B(n_477),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_533),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_539),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_532),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_531),
.A2(n_444),
.B1(n_454),
.B2(n_446),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_513),
.B(n_459),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_511),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_514),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_511),
.B(n_461),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_539),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_539),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_525),
.B(n_486),
.Y(n_613)
);

INVx6_ASAP7_75t_L g614 ( 
.A(n_542),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_513),
.B(n_462),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_538),
.B(n_486),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_511),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_539),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_525),
.B(n_463),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_541),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_541),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_541),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_541),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_525),
.B(n_490),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_514),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_529),
.B(n_490),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_544),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_536),
.B(n_466),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_534),
.B(n_474),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_536),
.B(n_487),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_534),
.B(n_488),
.Y(n_631)
);

AND2x6_ASAP7_75t_L g632 ( 
.A(n_536),
.B(n_219),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_544),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_544),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_544),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_554),
.B(n_491),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_522),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_554),
.B(n_495),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_575),
.B(n_493),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_511),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_564),
.B(n_496),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_514),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_542),
.B(n_469),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_511),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_538),
.A2(n_409),
.B1(n_414),
.B2(n_401),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_551),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_551),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_508),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_529),
.B(n_429),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_511),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_542),
.B(n_478),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_545),
.A2(n_352),
.B1(n_332),
.B2(n_422),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_508),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_508),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_501),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_501),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_501),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_522),
.Y(n_658)
);

AND2x2_ASAP7_75t_SL g659 ( 
.A(n_509),
.B(n_219),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_577),
.B(n_464),
.C(n_212),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_526),
.B(n_527),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_529),
.B(n_403),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_517),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_522),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_517),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_522),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_538),
.A2(n_386),
.B1(n_338),
.B2(n_353),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_517),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_511),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_529),
.B(n_493),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_518),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_511),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_542),
.B(n_467),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_515),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_515),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_L g676 ( 
.A(n_515),
.B(n_219),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_515),
.Y(n_677)
);

INVx6_ASAP7_75t_L g678 ( 
.A(n_542),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_515),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_515),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_545),
.A2(n_270),
.B1(n_372),
.B2(n_367),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_575),
.B(n_497),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_518),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_515),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_542),
.B(n_471),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_515),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_518),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_519),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_519),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_520),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_545),
.B(n_473),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_526),
.B(n_497),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_538),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_577),
.A2(n_472),
.B1(n_245),
.B2(n_344),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_575),
.B(n_380),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_530),
.A2(n_210),
.B1(n_361),
.B2(n_303),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_553),
.B(n_202),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_553),
.B(n_205),
.Y(n_698)
);

INVxp33_ASAP7_75t_L g699 ( 
.A(n_576),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_519),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_530),
.B(n_205),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_520),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_519),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_499),
.B(n_217),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_519),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_565),
.B(n_380),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_519),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_565),
.B(n_382),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_519),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_519),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_535),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_SL g712 ( 
.A(n_507),
.B(n_489),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_520),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_507),
.B(n_492),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_565),
.B(n_382),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_503),
.B(n_404),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_503),
.B(n_217),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_521),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_509),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_535),
.Y(n_720)
);

INVx8_ASAP7_75t_L g721 ( 
.A(n_565),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_565),
.B(n_222),
.Y(n_722)
);

OA22x2_ASAP7_75t_L g723 ( 
.A1(n_565),
.A2(n_362),
.B1(n_363),
.B2(n_355),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_602),
.B(n_510),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_585),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_693),
.B(n_521),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_585),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_693),
.B(n_521),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_588),
.A2(n_546),
.B1(n_510),
.B2(n_543),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_723),
.A2(n_509),
.B1(n_563),
.B2(n_546),
.Y(n_730)
);

OAI221xp5_ASAP7_75t_L g731 ( 
.A1(n_601),
.A2(n_379),
.B1(n_381),
.B2(n_388),
.C(n_323),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_579),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_579),
.B(n_405),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_646),
.B(n_528),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_655),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_655),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_584),
.B(n_408),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_602),
.B(n_592),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_721),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_646),
.B(n_528),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_647),
.B(n_528),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_647),
.B(n_537),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_656),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_657),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_602),
.B(n_516),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_657),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_663),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_593),
.B(n_537),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_663),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_665),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_592),
.B(n_516),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_665),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_593),
.B(n_537),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_L g754 ( 
.A(n_721),
.B(n_535),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_648),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_629),
.B(n_543),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_723),
.A2(n_509),
.B1(n_563),
.B2(n_556),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_631),
.B(n_547),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_691),
.B(n_573),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_714),
.A2(n_443),
.B1(n_460),
.B2(n_418),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_721),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_721),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_607),
.B(n_547),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_615),
.B(n_549),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_605),
.B(n_609),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_648),
.Y(n_766)
);

AO221x1_ASAP7_75t_L g767 ( 
.A1(n_652),
.A2(n_391),
.B1(n_397),
.B2(n_300),
.C(n_560),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_668),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_595),
.B(n_549),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_641),
.B(n_550),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_653),
.Y(n_771)
);

AND2x6_ASAP7_75t_SL g772 ( 
.A(n_716),
.B(n_576),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_668),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_653),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_695),
.B(n_550),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_661),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_593),
.B(n_535),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_637),
.B(n_535),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_695),
.B(n_560),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_654),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_580),
.B(n_419),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_613),
.A2(n_567),
.B(n_560),
.C(n_562),
.Y(n_782)
);

AND2x6_ASAP7_75t_L g783 ( 
.A(n_706),
.B(n_558),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_637),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_614),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_613),
.B(n_560),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_624),
.B(n_560),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_624),
.B(n_562),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_654),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_586),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_582),
.B(n_562),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_609),
.B(n_562),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_582),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_637),
.B(n_535),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_586),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_591),
.B(n_562),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_632),
.B(n_639),
.Y(n_797)
);

AO221x1_ASAP7_75t_L g798 ( 
.A1(n_696),
.A2(n_300),
.B1(n_567),
.B2(n_573),
.C(n_321),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_589),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_671),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_632),
.B(n_573),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_632),
.B(n_573),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_608),
.B(n_535),
.Y(n_803)
);

AOI22x1_ASAP7_75t_L g804 ( 
.A1(n_658),
.A2(n_540),
.B1(n_552),
.B2(n_535),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_616),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_616),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_683),
.Y(n_807)
);

INVxp33_ASAP7_75t_L g808 ( 
.A(n_692),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_632),
.B(n_558),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_608),
.B(n_540),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_639),
.B(n_682),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_683),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_723),
.A2(n_509),
.B1(n_556),
.B2(n_571),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_682),
.B(n_558),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_619),
.B(n_628),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_643),
.B(n_559),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_616),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_589),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_594),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_616),
.A2(n_559),
.B1(n_570),
.B2(n_509),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_630),
.B(n_433),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_625),
.A2(n_349),
.B1(n_243),
.B2(n_237),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_692),
.Y(n_823)
);

BUFx4f_ASAP7_75t_L g824 ( 
.A(n_659),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_606),
.B(n_214),
.C(n_212),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_712),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_659),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_687),
.A2(n_559),
.B(n_570),
.C(n_571),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_594),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_667),
.A2(n_556),
.B1(n_572),
.B2(n_574),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_658),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_708),
.B(n_572),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_SL g833 ( 
.A(n_625),
.B(n_447),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_687),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_664),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_596),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_581),
.B(n_220),
.C(n_214),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_636),
.B(n_449),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_642),
.B(n_455),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_690),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_598),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_715),
.B(n_572),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_614),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_681),
.A2(n_348),
.B1(n_231),
.B2(n_228),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_690),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_608),
.B(n_540),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_715),
.B(n_626),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_598),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_638),
.B(n_220),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_664),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_702),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_626),
.B(n_555),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_603),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_702),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_673),
.B(n_555),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_640),
.B(n_540),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_642),
.B(n_566),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_640),
.B(n_644),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_603),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_713),
.A2(n_552),
.B(n_540),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_722),
.A2(n_350),
.B1(n_222),
.B2(n_224),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_691),
.B(n_382),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_626),
.B(n_555),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_701),
.B(n_228),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_704),
.A2(n_234),
.B1(n_232),
.B2(n_230),
.Y(n_865)
);

BUFx8_ASAP7_75t_L g866 ( 
.A(n_699),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_649),
.B(n_231),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_681),
.B(n_574),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_645),
.B(n_574),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_618),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_618),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_697),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_713),
.A2(n_557),
.B(n_569),
.C(n_568),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_717),
.B(n_555),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_640),
.B(n_540),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_659),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_662),
.B(n_694),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_698),
.A2(n_234),
.B1(n_232),
.B2(n_230),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_719),
.A2(n_634),
.B1(n_623),
.B2(n_578),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_597),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_685),
.B(n_237),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_739),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_739),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_739),
.B(n_651),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_739),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_762),
.B(n_660),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_SL g887 ( 
.A(n_824),
.B(n_719),
.Y(n_887)
);

OAI21xp33_ASAP7_75t_SL g888 ( 
.A1(n_769),
.A2(n_718),
.B(n_670),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_762),
.B(n_640),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_761),
.B(n_640),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_816),
.A2(n_666),
.B(n_610),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_738),
.B(n_578),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_858),
.A2(n_666),
.B(n_672),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_877),
.A2(n_590),
.B(n_599),
.C(n_600),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_763),
.B(n_583),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_873),
.A2(n_782),
.B(n_860),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_858),
.A2(n_675),
.B(n_672),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_880),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_756),
.A2(n_679),
.B(n_675),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_764),
.B(n_583),
.Y(n_900)
);

AOI21xp33_ASAP7_75t_L g901 ( 
.A1(n_881),
.A2(n_590),
.B(n_587),
.Y(n_901)
);

O2A1O1Ixp5_ASAP7_75t_L g902 ( 
.A1(n_770),
.A2(n_623),
.B(n_634),
.C(n_611),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_811),
.A2(n_620),
.B1(n_621),
.B2(n_622),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_775),
.B(n_587),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_758),
.A2(n_635),
.B(n_599),
.C(n_600),
.Y(n_905)
);

BUFx12f_ASAP7_75t_L g906 ( 
.A(n_866),
.Y(n_906)
);

NOR2x1p5_ASAP7_75t_L g907 ( 
.A(n_733),
.B(n_243),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_734),
.A2(n_686),
.B(n_679),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_793),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_751),
.B(n_604),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_873),
.A2(n_611),
.B(n_604),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_868),
.B(n_792),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_734),
.A2(n_688),
.B(n_686),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_839),
.Y(n_914)
);

NAND2x1p5_ASAP7_75t_L g915 ( 
.A(n_806),
.B(n_597),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_735),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_740),
.A2(n_689),
.B(n_688),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_792),
.B(n_612),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_740),
.A2(n_700),
.B(n_689),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_761),
.B(n_644),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_737),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_872),
.B(n_612),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_880),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_741),
.A2(n_707),
.B(n_700),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_741),
.A2(n_710),
.B(n_707),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_824),
.B(n_644),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_880),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_783),
.A2(n_622),
.B1(n_633),
.B2(n_620),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_782),
.A2(n_627),
.B(n_621),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_824),
.B(n_644),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_742),
.A2(n_711),
.B(n_710),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_724),
.B(n_627),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_806),
.B(n_633),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_732),
.B(n_617),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_742),
.A2(n_874),
.B(n_778),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_806),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_786),
.A2(n_635),
.B(n_711),
.C(n_709),
.Y(n_937)
);

AOI21x1_ASAP7_75t_L g938 ( 
.A1(n_803),
.A2(n_557),
.B(n_566),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_791),
.B(n_644),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_736),
.B(n_669),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_777),
.A2(n_674),
.B(n_617),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_847),
.B(n_650),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_SL g943 ( 
.A1(n_777),
.A2(n_794),
.B(n_778),
.C(n_753),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_794),
.A2(n_674),
.B(n_617),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_783),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_796),
.A2(n_677),
.B(n_674),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_743),
.Y(n_947)
);

BUFx4f_ASAP7_75t_L g948 ( 
.A(n_783),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_787),
.A2(n_720),
.B(n_709),
.C(n_705),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_745),
.B(n_680),
.Y(n_950)
);

OAI321xp33_ASAP7_75t_L g951 ( 
.A1(n_731),
.A2(n_574),
.A3(n_568),
.B1(n_569),
.B2(n_556),
.C(n_326),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_727),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_SL g953 ( 
.A(n_817),
.B(n_224),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_869),
.B(n_680),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_817),
.B(n_650),
.Y(n_955)
);

AND2x6_ASAP7_75t_L g956 ( 
.A(n_820),
.B(n_650),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_748),
.A2(n_684),
.B(n_680),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_862),
.B(n_684),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_817),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_781),
.B(n_684),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_808),
.B(n_823),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_765),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_808),
.B(n_725),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_744),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_753),
.A2(n_703),
.B(n_650),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_779),
.B(n_759),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_864),
.A2(n_557),
.B(n_703),
.C(n_569),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_833),
.B(n_650),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_746),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_747),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_788),
.B(n_568),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_783),
.B(n_568),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_776),
.B(n_614),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_729),
.A2(n_676),
.B(n_566),
.Y(n_974)
);

NAND2x1p5_ASAP7_75t_L g975 ( 
.A(n_805),
.B(n_556),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_783),
.B(n_569),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_805),
.Y(n_977)
);

AO21x1_ASAP7_75t_L g978 ( 
.A1(n_726),
.A2(n_728),
.B(n_749),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_750),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_866),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_815),
.B(n_614),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_783),
.B(n_556),
.Y(n_982)
);

O2A1O1Ixp5_ASAP7_75t_L g983 ( 
.A1(n_832),
.A2(n_498),
.B(n_502),
.C(n_504),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_752),
.A2(n_293),
.B(n_360),
.C(n_302),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_821),
.B(n_678),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_880),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_826),
.B(n_225),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_768),
.A2(n_292),
.B(n_304),
.C(n_310),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_755),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_785),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_773),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_825),
.B(n_678),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_826),
.B(n_225),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_866),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_800),
.B(n_552),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_785),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_760),
.B(n_244),
.Y(n_997)
);

INVx8_ASAP7_75t_L g998 ( 
.A(n_857),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_797),
.A2(n_255),
.B(n_239),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_857),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_842),
.B(n_227),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_810),
.A2(n_552),
.B(n_502),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_807),
.A2(n_359),
.B1(n_343),
.B2(n_344),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_784),
.B(n_342),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_812),
.A2(n_279),
.B(n_297),
.C(n_257),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_834),
.Y(n_1006)
);

O2A1O1Ixp5_ASAP7_75t_L g1007 ( 
.A1(n_810),
.A2(n_498),
.B(n_502),
.C(n_504),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_766),
.Y(n_1008)
);

NOR2xp67_ASAP7_75t_L g1009 ( 
.A(n_838),
.B(n_556),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_784),
.B(n_342),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_867),
.B(n_244),
.Y(n_1011)
);

AND2x6_ASAP7_75t_L g1012 ( 
.A(n_840),
.B(n_300),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_843),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_843),
.Y(n_1014)
);

NOR2xp67_ASAP7_75t_L g1015 ( 
.A(n_849),
.B(n_556),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_827),
.A2(n_678),
.B1(n_364),
.B2(n_374),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_845),
.A2(n_267),
.B(n_324),
.C(n_346),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_814),
.B(n_678),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_851),
.A2(n_336),
.B(n_354),
.C(n_376),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_843),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_854),
.B(n_552),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_828),
.A2(n_399),
.B(n_383),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_784),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_878),
.B(n_350),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_852),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_831),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_831),
.A2(n_387),
.B(n_343),
.C(n_367),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_837),
.B(n_351),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_863),
.B(n_347),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_879),
.A2(n_506),
.B(n_505),
.Y(n_1030)
);

AOI33xp33_ASAP7_75t_L g1031 ( 
.A1(n_861),
.A2(n_347),
.A3(n_348),
.B1(n_349),
.B2(n_358),
.B3(n_359),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_855),
.B(n_358),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_876),
.B(n_361),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_772),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_827),
.B(n_366),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_857),
.B(n_366),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_822),
.B(n_372),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_876),
.B(n_398),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_831),
.A2(n_389),
.B(n_357),
.C(n_394),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_835),
.B(n_351),
.Y(n_1040)
);

NAND2x1_ASAP7_75t_L g1041 ( 
.A(n_835),
.B(n_502),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_865),
.B(n_357),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_771),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_754),
.A2(n_504),
.B(n_9),
.C(n_11),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_730),
.A2(n_364),
.B1(n_394),
.B2(n_393),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_857),
.B(n_374),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_835),
.B(n_385),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_767),
.B(n_385),
.Y(n_1048)
);

OR2x2_ASAP7_75t_SL g1049 ( 
.A(n_809),
.B(n_300),
.Y(n_1049)
);

INVx5_ASAP7_75t_L g1050 ( 
.A(n_850),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_850),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_850),
.B(n_389),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_790),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_813),
.A2(n_392),
.B1(n_393),
.B2(n_284),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_790),
.B(n_504),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_882),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_916),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_895),
.A2(n_754),
.B(n_726),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_961),
.B(n_728),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_914),
.B(n_757),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_895),
.A2(n_875),
.B(n_846),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_900),
.A2(n_875),
.B(n_856),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_900),
.A2(n_856),
.B(n_870),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_910),
.A2(n_904),
.B(n_935),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_946),
.A2(n_871),
.B(n_870),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_912),
.B(n_871),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_914),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_909),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1011),
.B(n_830),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_997),
.B(n_795),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_921),
.A2(n_798),
.B1(n_780),
.B2(n_789),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_963),
.A2(n_801),
.B1(n_802),
.B2(n_848),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_906),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_887),
.Y(n_1074)
);

AOI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_1045),
.A2(n_771),
.B(n_774),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_962),
.B(n_799),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_952),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_911),
.A2(n_804),
.B(n_780),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_947),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_964),
.Y(n_1080)
);

BUFx8_ASAP7_75t_L g1081 ( 
.A(n_980),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1025),
.B(n_799),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_985),
.B(n_818),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_1036),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_960),
.A2(n_1022),
.B(n_888),
.C(n_981),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_994),
.B(n_818),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_945),
.B(n_819),
.Y(n_1087)
);

BUFx4f_ASAP7_75t_L g1088 ( 
.A(n_998),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_966),
.B(n_819),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_945),
.A2(n_859),
.B1(n_853),
.B2(n_848),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_948),
.A2(n_836),
.B1(n_853),
.B2(n_841),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1036),
.B(n_829),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_948),
.A2(n_829),
.B1(n_789),
.B2(n_774),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_882),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_907),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_969),
.A2(n_979),
.B1(n_991),
.B2(n_970),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_953),
.A2(n_392),
.B1(n_337),
.B2(n_333),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_891),
.A2(n_329),
.B(n_328),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_968),
.B(n_246),
.Y(n_1099)
);

BUFx5_ASAP7_75t_L g1100 ( 
.A(n_956),
.Y(n_1100)
);

BUFx8_ASAP7_75t_L g1101 ( 
.A(n_1046),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_998),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_SL g1103 ( 
.A(n_953),
.B(n_252),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_882),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1006),
.A2(n_325),
.B1(n_317),
.B2(n_307),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_933),
.B(n_306),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_903),
.A2(n_301),
.B(n_253),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1024),
.A2(n_1022),
.B(n_1027),
.C(n_1001),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_885),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1000),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_885),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_892),
.B(n_8),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_885),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_933),
.B(n_254),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1034),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_977),
.Y(n_1116)
);

BUFx4f_ASAP7_75t_L g1117 ( 
.A(n_998),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1037),
.B(n_1003),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_934),
.B(n_990),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_1013),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_932),
.B(n_8),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_928),
.A2(n_269),
.B1(n_298),
.B2(n_296),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1003),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_990),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_990),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_903),
.A2(n_265),
.B1(n_295),
.B2(n_294),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_956),
.A2(n_263),
.B1(n_283),
.B2(n_282),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_973),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_899),
.A2(n_261),
.B(n_275),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1031),
.B(n_12),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_898),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_897),
.A2(n_266),
.B(n_262),
.Y(n_1132)
);

O2A1O1Ixp5_ASAP7_75t_L g1133 ( 
.A1(n_896),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_943),
.A2(n_259),
.B(n_258),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_887),
.B(n_956),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_987),
.B(n_256),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_989),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1008),
.Y(n_1138)
);

AND2x2_ASAP7_75t_SL g1139 ( 
.A(n_936),
.B(n_300),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_993),
.B(n_17),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1043),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_898),
.Y(n_1142)
);

OAI21xp33_ASAP7_75t_L g1143 ( 
.A1(n_1029),
.A2(n_18),
.B(n_19),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_893),
.A2(n_196),
.B(n_181),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_908),
.A2(n_178),
.B(n_170),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_918),
.B(n_22),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_886),
.B(n_24),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1023),
.B(n_26),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_922),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_SL g1150 ( 
.A(n_898),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1053),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_958),
.A2(n_29),
.B(n_30),
.C(n_33),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_R g1153 ( 
.A(n_936),
.B(n_164),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_923),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_SL g1155 ( 
.A1(n_896),
.A2(n_33),
.B(n_34),
.C(n_37),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1023),
.B(n_954),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_913),
.A2(n_157),
.B(n_152),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_956),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_1158)
);

NAND2x2_ASAP7_75t_L g1159 ( 
.A(n_1032),
.B(n_40),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_940),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_971),
.B(n_42),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_959),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_959),
.B(n_71),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_923),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1053),
.B(n_44),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_923),
.Y(n_1166)
);

BUFx12f_ASAP7_75t_L g1167 ( 
.A(n_927),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1045),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_975),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_940),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1033),
.B(n_46),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_995),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1035),
.B(n_48),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_894),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_1174)
);

OAI21xp33_ASAP7_75t_SL g1175 ( 
.A1(n_972),
.A2(n_55),
.B(n_57),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_883),
.B(n_61),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_917),
.A2(n_78),
.B(n_125),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1038),
.B(n_62),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_996),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_919),
.A2(n_75),
.B(n_118),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1009),
.B(n_62),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_996),
.B(n_63),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_927),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1050),
.B(n_65),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1042),
.A2(n_65),
.B(n_68),
.C(n_69),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_924),
.A2(n_72),
.B(n_73),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1048),
.B(n_1028),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1004),
.B(n_1010),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1026),
.B(n_84),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1044),
.A2(n_999),
.B(n_901),
.C(n_992),
.Y(n_1190)
);

CKINVDCx6p67_ASAP7_75t_R g1191 ( 
.A(n_1050),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1054),
.A2(n_999),
.B1(n_901),
.B2(n_976),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1054),
.A2(n_88),
.B1(n_89),
.B2(n_95),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_951),
.A2(n_104),
.B(n_150),
.C(n_974),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_984),
.A2(n_1005),
.B(n_1017),
.C(n_988),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1050),
.B(n_1026),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1016),
.A2(n_978),
.B1(n_884),
.B2(n_930),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_925),
.A2(n_931),
.B(n_911),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1055),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1026),
.B(n_1040),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_950),
.B(n_1050),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1047),
.B(n_1052),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1051),
.B(n_883),
.Y(n_1203)
);

O2A1O1Ixp5_ASAP7_75t_L g1204 ( 
.A1(n_939),
.A2(n_967),
.B(n_889),
.C(n_942),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1051),
.B(n_905),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_R g1206 ( 
.A(n_927),
.B(n_986),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1039),
.B(n_986),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_929),
.B(n_1018),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1057),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1085),
.A2(n_929),
.B(n_1021),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1078),
.A2(n_983),
.B(n_938),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1064),
.A2(n_949),
.B(n_937),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1081),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1208),
.A2(n_982),
.B(n_1015),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1178),
.A2(n_951),
.B(n_1019),
.C(n_974),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1149),
.B(n_986),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1108),
.A2(n_902),
.B(n_926),
.C(n_955),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1065),
.A2(n_1007),
.B(n_1002),
.Y(n_1218)
);

CKINVDCx8_ASAP7_75t_R g1219 ( 
.A(n_1115),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1190),
.A2(n_1055),
.A3(n_965),
.B(n_941),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1058),
.A2(n_944),
.B(n_957),
.Y(n_1221)
);

INVxp67_ASAP7_75t_SL g1222 ( 
.A(n_1067),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1202),
.A2(n_1195),
.B(n_1194),
.C(n_1147),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1102),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1061),
.A2(n_1030),
.B(n_890),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1128),
.B(n_975),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1068),
.B(n_920),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1079),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1081),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1205),
.A2(n_1020),
.B(n_1041),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1118),
.A2(n_1059),
.B(n_1140),
.C(n_1143),
.Y(n_1231)
);

CKINVDCx11_ASAP7_75t_R g1232 ( 
.A(n_1073),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1135),
.A2(n_1020),
.B(n_1014),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1126),
.A2(n_1014),
.B1(n_1049),
.B2(n_915),
.Y(n_1234)
);

NAND3x1_ASAP7_75t_L g1235 ( 
.A(n_1158),
.B(n_1030),
.C(n_1012),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1068),
.B(n_915),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1204),
.A2(n_1012),
.B(n_1063),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1077),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1166),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_SL g1240 ( 
.A1(n_1148),
.A2(n_1012),
.B(n_1121),
.C(n_1112),
.Y(n_1240)
);

INVxp67_ASAP7_75t_L g1241 ( 
.A(n_1116),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1090),
.A2(n_1012),
.A3(n_1093),
.B(n_1091),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1088),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1080),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1084),
.B(n_1110),
.Y(n_1245)
);

BUFx10_ASAP7_75t_L g1246 ( 
.A(n_1150),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1103),
.A2(n_1069),
.B1(n_1174),
.B2(n_1135),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_1150),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1062),
.A2(n_1201),
.B(n_1083),
.Y(n_1249)
);

BUFx12f_ASAP7_75t_L g1250 ( 
.A(n_1101),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1070),
.B(n_1092),
.Y(n_1251)
);

OAI21xp33_ASAP7_75t_L g1252 ( 
.A1(n_1168),
.A2(n_1103),
.B(n_1174),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1171),
.A2(n_1173),
.B(n_1188),
.C(n_1192),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1102),
.B(n_1124),
.Y(n_1254)
);

NAND3x1_ASAP7_75t_L g1255 ( 
.A(n_1086),
.B(n_1130),
.C(n_1187),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1096),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1161),
.A2(n_1112),
.B(n_1121),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1144),
.A2(n_1177),
.B(n_1186),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1145),
.A2(n_1180),
.B(n_1157),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1185),
.A2(n_1207),
.B(n_1200),
.C(n_1123),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1125),
.B(n_1131),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1167),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1138),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1172),
.A2(n_1170),
.B(n_1160),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1197),
.A2(n_1136),
.B(n_1139),
.C(n_1152),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1176),
.B(n_1095),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1089),
.A2(n_1161),
.B(n_1156),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1156),
.A2(n_1146),
.B(n_1075),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1075),
.A2(n_1066),
.B(n_1133),
.Y(n_1269)
);

AOI221x1_ASAP7_75t_L g1270 ( 
.A1(n_1126),
.A2(n_1181),
.B1(n_1146),
.B2(n_1122),
.C(n_1148),
.Y(n_1270)
);

AOI221x1_ASAP7_75t_L g1271 ( 
.A1(n_1122),
.A2(n_1182),
.B1(n_1165),
.B2(n_1096),
.C(n_1107),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1141),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1155),
.A2(n_1105),
.B(n_1175),
.C(n_1114),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1088),
.Y(n_1274)
);

AO22x1_ASAP7_75t_L g1275 ( 
.A1(n_1101),
.A2(n_1176),
.B1(n_1074),
.B2(n_1060),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1142),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1127),
.A2(n_1097),
.B(n_1193),
.C(n_1072),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1105),
.B(n_1117),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1199),
.A2(n_1119),
.B(n_1066),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1203),
.A2(n_1196),
.B(n_1082),
.Y(n_1280)
);

NOR2xp67_ASAP7_75t_L g1281 ( 
.A(n_1162),
.B(n_1120),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1087),
.A2(n_1162),
.B(n_1165),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1120),
.A2(n_1098),
.B(n_1184),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1117),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1076),
.B(n_1179),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1137),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1151),
.B(n_1106),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1159),
.A2(n_1169),
.B1(n_1191),
.B2(n_1163),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1134),
.A2(n_1129),
.B(n_1132),
.C(n_1189),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1164),
.B(n_1099),
.Y(n_1290)
);

NAND3xp33_ASAP7_75t_SL g1291 ( 
.A(n_1153),
.B(n_1071),
.C(n_1206),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1154),
.A2(n_1183),
.B(n_1094),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1154),
.Y(n_1293)
);

NOR2x1_ASAP7_75t_SL g1294 ( 
.A(n_1183),
.B(n_1056),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1056),
.A2(n_1094),
.B(n_1104),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1094),
.B(n_1104),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1104),
.A2(n_1109),
.B(n_1111),
.Y(n_1297)
);

BUFx10_ASAP7_75t_L g1298 ( 
.A(n_1109),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1100),
.A2(n_1109),
.B(n_1111),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1111),
.A2(n_641),
.B(n_595),
.C(n_1178),
.Y(n_1300)
);

OA21x2_ASAP7_75t_L g1301 ( 
.A1(n_1100),
.A2(n_1198),
.B(n_896),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1113),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1113),
.A2(n_1085),
.B(n_641),
.Y(n_1303)
);

BUFx10_ASAP7_75t_L g1304 ( 
.A(n_1100),
.Y(n_1304)
);

INVxp67_ASAP7_75t_L g1305 ( 
.A(n_1100),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1118),
.A2(n_877),
.B1(n_1103),
.B2(n_531),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1190),
.A2(n_967),
.A3(n_1194),
.B(n_1091),
.Y(n_1307)
);

AOI221xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1174),
.A2(n_1168),
.B1(n_1123),
.B2(n_1143),
.C(n_1185),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1102),
.B(n_998),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1067),
.B(n_579),
.Y(n_1310)
);

INVx4_ASAP7_75t_L g1311 ( 
.A(n_1167),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1149),
.B(n_585),
.Y(n_1312)
);

NAND3xp33_ASAP7_75t_L g1313 ( 
.A(n_1085),
.B(n_1168),
.C(n_881),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1118),
.A2(n_877),
.B1(n_1103),
.B2(n_531),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1085),
.A2(n_1064),
.B(n_948),
.Y(n_1315)
);

NOR4xp25_ASAP7_75t_L g1316 ( 
.A(n_1123),
.B(n_1143),
.C(n_1174),
.D(n_1168),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1198),
.A2(n_1078),
.B(n_1065),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1190),
.A2(n_967),
.A3(n_1194),
.B(n_1091),
.Y(n_1318)
);

NOR2x1_ASAP7_75t_SL g1319 ( 
.A(n_1162),
.B(n_1196),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1081),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_L g1321 ( 
.A1(n_1118),
.A2(n_844),
.B1(n_652),
.B2(n_696),
.C(n_1011),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1198),
.A2(n_1078),
.B(n_1065),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1178),
.A2(n_641),
.B(n_595),
.C(n_1108),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1198),
.A2(n_1078),
.B(n_1065),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1085),
.A2(n_948),
.B1(n_945),
.B2(n_595),
.Y(n_1325)
);

AND3x4_ASAP7_75t_L g1326 ( 
.A(n_1073),
.B(n_837),
.C(n_1036),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1085),
.A2(n_1064),
.B(n_948),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1085),
.A2(n_1064),
.B(n_948),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1085),
.A2(n_1064),
.B(n_948),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1073),
.Y(n_1330)
);

INVx4_ASAP7_75t_SL g1331 ( 
.A(n_1073),
.Y(n_1331)
);

OR2x6_ASAP7_75t_L g1332 ( 
.A(n_1102),
.B(n_998),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1118),
.B(n_585),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1077),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1118),
.B(n_585),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1102),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1085),
.A2(n_1064),
.B(n_948),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1149),
.B(n_585),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_L g1339 ( 
.A(n_1085),
.B(n_1168),
.C(n_881),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1198),
.A2(n_1078),
.B(n_1065),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1085),
.A2(n_1194),
.B(n_1190),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1198),
.A2(n_1078),
.B(n_1065),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1149),
.B(n_585),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1077),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1085),
.A2(n_948),
.B1(n_945),
.B2(n_595),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1085),
.A2(n_1064),
.B(n_948),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1190),
.A2(n_967),
.A3(n_1194),
.B(n_1091),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1190),
.A2(n_967),
.A3(n_1194),
.B(n_1091),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1198),
.A2(n_1078),
.B(n_1065),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1085),
.A2(n_948),
.B1(n_945),
.B2(n_595),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1085),
.A2(n_595),
.B(n_641),
.C(n_561),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1085),
.A2(n_1194),
.B(n_1190),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1178),
.A2(n_641),
.B(n_595),
.C(n_1108),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1077),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1085),
.A2(n_1064),
.B(n_948),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1198),
.A2(n_896),
.B(n_1078),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1085),
.A2(n_1194),
.B(n_1190),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_SL g1358 ( 
.A1(n_1085),
.A2(n_1194),
.B(n_1205),
.C(n_1148),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1085),
.A2(n_1064),
.B(n_948),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1190),
.A2(n_967),
.A3(n_1194),
.B(n_1091),
.Y(n_1360)
);

BUFx8_ASAP7_75t_SL g1361 ( 
.A(n_1320),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1238),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1252),
.A2(n_1306),
.B1(n_1314),
.B2(n_1321),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1333),
.B(n_1335),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1330),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1334),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1246),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1222),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1313),
.A2(n_1339),
.B1(n_1341),
.B2(n_1352),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1313),
.A2(n_1339),
.B1(n_1341),
.B2(n_1352),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1344),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1228),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1244),
.Y(n_1373)
);

OAI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1306),
.A2(n_1314),
.B1(n_1247),
.B2(n_1357),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1250),
.Y(n_1375)
);

INVx6_ASAP7_75t_L g1376 ( 
.A(n_1246),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1312),
.B(n_1338),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1243),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1343),
.B(n_1310),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1323),
.A2(n_1353),
.B1(n_1231),
.B2(n_1223),
.Y(n_1380)
);

BUFx4f_ASAP7_75t_SL g1381 ( 
.A(n_1274),
.Y(n_1381)
);

BUFx4f_ASAP7_75t_SL g1382 ( 
.A(n_1274),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1252),
.A2(n_1247),
.B1(n_1357),
.B2(n_1257),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1278),
.A2(n_1326),
.B1(n_1291),
.B2(n_1265),
.Y(n_1384)
);

AOI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1308),
.A2(n_1300),
.B1(n_1215),
.B2(n_1345),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_1213),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1256),
.A2(n_1270),
.B1(n_1325),
.B2(n_1350),
.Y(n_1387)
);

INVx4_ASAP7_75t_L g1388 ( 
.A(n_1243),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1219),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1351),
.A2(n_1253),
.B(n_1277),
.Y(n_1390)
);

BUFx12f_ASAP7_75t_L g1391 ( 
.A(n_1248),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1248),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1276),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1257),
.A2(n_1251),
.B1(n_1286),
.B2(n_1303),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1331),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1271),
.A2(n_1285),
.B1(n_1241),
.B2(n_1210),
.Y(n_1396)
);

INVx4_ASAP7_75t_SL g1397 ( 
.A(n_1309),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1268),
.A2(n_1263),
.B1(n_1272),
.B2(n_1287),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1216),
.Y(n_1399)
);

BUFx8_ASAP7_75t_L g1400 ( 
.A(n_1229),
.Y(n_1400)
);

AOI22x1_ASAP7_75t_L g1401 ( 
.A1(n_1283),
.A2(n_1327),
.B1(n_1359),
.B2(n_1315),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1260),
.A2(n_1354),
.B1(n_1227),
.B2(n_1273),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1331),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1293),
.Y(n_1404)
);

BUFx4f_ASAP7_75t_SL g1405 ( 
.A(n_1284),
.Y(n_1405)
);

BUFx2_ASAP7_75t_SL g1406 ( 
.A(n_1311),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1239),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1236),
.Y(n_1408)
);

INVxp67_ASAP7_75t_SL g1409 ( 
.A(n_1301),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1316),
.A2(n_1234),
.B1(n_1308),
.B2(n_1268),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1267),
.A2(n_1245),
.B1(n_1269),
.B2(n_1316),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1269),
.A2(n_1264),
.B1(n_1266),
.B2(n_1301),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1309),
.B(n_1332),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1262),
.Y(n_1414)
);

BUFx8_ASAP7_75t_SL g1415 ( 
.A(n_1284),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1279),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1255),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1284),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1311),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1296),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1288),
.A2(n_1290),
.B1(n_1226),
.B2(n_1329),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1235),
.A2(n_1328),
.B1(n_1337),
.B2(n_1355),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1346),
.A2(n_1261),
.B1(n_1332),
.B2(n_1309),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1261),
.A2(n_1332),
.B1(n_1225),
.B2(n_1254),
.Y(n_1424)
);

CKINVDCx11_ASAP7_75t_R g1425 ( 
.A(n_1298),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1275),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1225),
.A2(n_1358),
.B1(n_1360),
.B2(n_1307),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1254),
.Y(n_1428)
);

BUFx12f_ASAP7_75t_L g1429 ( 
.A(n_1298),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1302),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1299),
.Y(n_1431)
);

INVx6_ASAP7_75t_L g1432 ( 
.A(n_1304),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1294),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1214),
.A2(n_1356),
.B1(n_1280),
.B2(n_1249),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1224),
.A2(n_1336),
.B1(n_1281),
.B2(n_1217),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1336),
.Y(n_1436)
);

INVx6_ASAP7_75t_L g1437 ( 
.A(n_1304),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1292),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1319),
.Y(n_1439)
);

BUFx12f_ASAP7_75t_L g1440 ( 
.A(n_1295),
.Y(n_1440)
);

CKINVDCx6p67_ASAP7_75t_R g1441 ( 
.A(n_1297),
.Y(n_1441)
);

BUFx12f_ASAP7_75t_L g1442 ( 
.A(n_1281),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1282),
.A2(n_1289),
.B1(n_1233),
.B2(n_1230),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1220),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1307),
.B(n_1360),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1220),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1212),
.A2(n_1305),
.B1(n_1356),
.B2(n_1221),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1258),
.A2(n_1259),
.B(n_1240),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1307),
.A2(n_1318),
.B1(n_1348),
.B2(n_1347),
.Y(n_1449)
);

INVx6_ASAP7_75t_L g1450 ( 
.A(n_1242),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1237),
.A2(n_1360),
.B1(n_1348),
.B2(n_1347),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1318),
.A2(n_1348),
.B1(n_1347),
.B2(n_1242),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1211),
.A2(n_1218),
.B1(n_1317),
.B2(n_1322),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1324),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1349),
.A2(n_1306),
.B1(n_1314),
.B2(n_1323),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1340),
.A2(n_1252),
.B1(n_1118),
.B2(n_1306),
.Y(n_1456)
);

CKINVDCx11_ASAP7_75t_R g1457 ( 
.A(n_1342),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1238),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1306),
.A2(n_1314),
.B1(n_1247),
.B2(n_1103),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1313),
.A2(n_1118),
.B1(n_531),
.B2(n_1339),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1219),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1252),
.A2(n_1118),
.B1(n_1314),
.B2(n_1306),
.Y(n_1462)
);

NAND2x1p5_ASAP7_75t_L g1463 ( 
.A(n_1274),
.B(n_1088),
.Y(n_1463)
);

INVx6_ASAP7_75t_L g1464 ( 
.A(n_1246),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1232),
.Y(n_1465)
);

OAI21xp33_ASAP7_75t_L g1466 ( 
.A1(n_1323),
.A2(n_1353),
.B(n_1253),
.Y(n_1466)
);

CKINVDCx11_ASAP7_75t_R g1467 ( 
.A(n_1219),
.Y(n_1467)
);

INVx6_ASAP7_75t_L g1468 ( 
.A(n_1246),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1209),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1306),
.A2(n_1314),
.B1(n_1247),
.B2(n_1103),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1252),
.A2(n_1118),
.B1(n_1314),
.B2(n_1306),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1320),
.Y(n_1472)
);

CKINVDCx11_ASAP7_75t_R g1473 ( 
.A(n_1219),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1320),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1306),
.A2(n_1314),
.B1(n_1247),
.B2(n_1103),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1320),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1243),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1252),
.A2(n_1118),
.B1(n_1314),
.B2(n_1306),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1333),
.B(n_1335),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1209),
.Y(n_1480)
);

INVx8_ASAP7_75t_L g1481 ( 
.A(n_1320),
.Y(n_1481)
);

CKINVDCx11_ASAP7_75t_R g1482 ( 
.A(n_1219),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1243),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1243),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1222),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1306),
.A2(n_1314),
.B1(n_1247),
.B2(n_1103),
.Y(n_1486)
);

BUFx12f_ASAP7_75t_L g1487 ( 
.A(n_1232),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1232),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1320),
.Y(n_1489)
);

AO22x1_ASAP7_75t_L g1490 ( 
.A1(n_1326),
.A2(n_582),
.B1(n_1118),
.B2(n_530),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1209),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1333),
.B(n_1335),
.Y(n_1492)
);

OAI22x1_ASAP7_75t_L g1493 ( 
.A1(n_1306),
.A2(n_1314),
.B1(n_1247),
.B2(n_1326),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1209),
.Y(n_1494)
);

INVxp33_ASAP7_75t_SL g1495 ( 
.A(n_1232),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1209),
.Y(n_1496)
);

CKINVDCx11_ASAP7_75t_R g1497 ( 
.A(n_1219),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1429),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1416),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1479),
.B(n_1492),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1368),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1445),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1397),
.B(n_1413),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1444),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1383),
.A2(n_1363),
.B1(n_1385),
.B2(n_1384),
.Y(n_1505)
);

INVx4_ASAP7_75t_SL g1506 ( 
.A(n_1450),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1449),
.B(n_1456),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1372),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1459),
.A2(n_1475),
.B(n_1470),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1393),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1373),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1485),
.Y(n_1512)
);

AO32x2_ASAP7_75t_L g1513 ( 
.A1(n_1455),
.A2(n_1380),
.A3(n_1447),
.B1(n_1402),
.B2(n_1422),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1490),
.B(n_1389),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1457),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1469),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1480),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1448),
.A2(n_1434),
.B(n_1409),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1449),
.B(n_1456),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1491),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1494),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1466),
.A2(n_1390),
.B(n_1459),
.C(n_1486),
.Y(n_1522)
);

CKINVDCx6p67_ASAP7_75t_R g1523 ( 
.A(n_1395),
.Y(n_1523)
);

AO31x2_ASAP7_75t_L g1524 ( 
.A1(n_1493),
.A2(n_1446),
.A3(n_1443),
.B(n_1448),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1379),
.B(n_1364),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1432),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1362),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1496),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1452),
.B(n_1383),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1431),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1451),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1397),
.B(n_1413),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1401),
.A2(n_1434),
.B(n_1454),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1431),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1414),
.Y(n_1535)
);

AND2x2_ASAP7_75t_SL g1536 ( 
.A(n_1363),
.B(n_1462),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1397),
.B(n_1423),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1452),
.A2(n_1411),
.B(n_1412),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1408),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1423),
.B(n_1412),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1399),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1460),
.A2(n_1475),
.B1(n_1486),
.B2(n_1470),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1411),
.A2(n_1435),
.B(n_1417),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1404),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1439),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1374),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1471),
.A2(n_1478),
.B(n_1398),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1374),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1365),
.Y(n_1549)
);

OA21x2_ASAP7_75t_L g1550 ( 
.A1(n_1471),
.A2(n_1478),
.B(n_1398),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1420),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1427),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1410),
.B(n_1369),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1369),
.A2(n_1370),
.B(n_1387),
.Y(n_1554)
);

OA21x2_ASAP7_75t_L g1555 ( 
.A1(n_1394),
.A2(n_1424),
.B(n_1421),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1396),
.A2(n_1387),
.B(n_1377),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1410),
.B(n_1370),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1427),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1394),
.B(n_1424),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1396),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1453),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1441),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1366),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1460),
.A2(n_1426),
.B1(n_1421),
.B2(n_1438),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1440),
.A2(n_1433),
.B1(n_1407),
.B2(n_1428),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1436),
.Y(n_1566)
);

INVx4_ASAP7_75t_L g1567 ( 
.A(n_1437),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1437),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1371),
.B(n_1458),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1461),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1418),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1367),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1442),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1430),
.B(n_1418),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1378),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1378),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_1381),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1477),
.Y(n_1578)
);

NAND4xp25_ASAP7_75t_L g1579 ( 
.A(n_1419),
.B(n_1495),
.C(n_1388),
.D(n_1483),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1484),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1425),
.B(n_1392),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1376),
.Y(n_1582)
);

INVxp67_ASAP7_75t_SL g1583 ( 
.A(n_1463),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1392),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1464),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1464),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1381),
.A2(n_1382),
.B1(n_1406),
.B2(n_1419),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1465),
.A2(n_1403),
.B1(n_1474),
.B2(n_1472),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1468),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1468),
.B(n_1386),
.Y(n_1590)
);

INVx3_ASAP7_75t_L g1591 ( 
.A(n_1468),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1481),
.B(n_1489),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1382),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1386),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1405),
.Y(n_1595)
);

AOI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1405),
.A2(n_1391),
.B(n_1415),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1481),
.A2(n_1476),
.B(n_1400),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1500),
.B(n_1473),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1512),
.B(n_1400),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1500),
.B(n_1497),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1563),
.B(n_1467),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1554),
.A2(n_1481),
.B(n_1482),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1527),
.B(n_1488),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1522),
.A2(n_1375),
.B(n_1361),
.C(n_1487),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1553),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1543),
.A2(n_1533),
.B(n_1561),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1501),
.B(n_1512),
.Y(n_1607)
);

AO32x1_ASAP7_75t_L g1608 ( 
.A1(n_1553),
.A2(n_1557),
.A3(n_1505),
.B1(n_1560),
.B2(n_1558),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1515),
.B(n_1569),
.Y(n_1609)
);

INVx5_ASAP7_75t_SL g1610 ( 
.A(n_1523),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1508),
.Y(n_1611)
);

NOR2x1_ASAP7_75t_SL g1612 ( 
.A(n_1509),
.B(n_1562),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1557),
.B(n_1556),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1508),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1536),
.A2(n_1509),
.B1(n_1542),
.B2(n_1559),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1515),
.B(n_1566),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1549),
.A2(n_1514),
.B1(n_1570),
.B2(n_1559),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1581),
.A2(n_1555),
.B1(n_1573),
.B2(n_1597),
.Y(n_1618)
);

AOI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1560),
.A2(n_1548),
.B1(n_1546),
.B2(n_1552),
.C(n_1558),
.Y(n_1619)
);

AO32x2_ASAP7_75t_L g1620 ( 
.A1(n_1572),
.A2(n_1526),
.A3(n_1567),
.B1(n_1587),
.B2(n_1577),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1546),
.B(n_1548),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1545),
.B(n_1581),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1545),
.B(n_1578),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1511),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1511),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1536),
.A2(n_1529),
.B1(n_1555),
.B2(n_1564),
.Y(n_1626)
);

AOI221xp5_ASAP7_75t_L g1627 ( 
.A1(n_1552),
.A2(n_1529),
.B1(n_1531),
.B2(n_1525),
.C(n_1519),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1536),
.A2(n_1550),
.B1(n_1547),
.B2(n_1555),
.Y(n_1628)
);

OR2x6_ASAP7_75t_L g1629 ( 
.A(n_1537),
.B(n_1540),
.Y(n_1629)
);

OAI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1555),
.A2(n_1550),
.B(n_1547),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1540),
.A2(n_1519),
.B(n_1507),
.C(n_1531),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1499),
.B(n_1502),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1547),
.A2(n_1550),
.B1(n_1538),
.B2(n_1537),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1518),
.A2(n_1499),
.B(n_1513),
.Y(n_1634)
);

AO21x1_ASAP7_75t_L g1635 ( 
.A1(n_1544),
.A2(n_1517),
.B(n_1516),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_R g1636 ( 
.A(n_1596),
.B(n_1523),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1517),
.A2(n_1528),
.B1(n_1521),
.B2(n_1520),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1506),
.B(n_1503),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1538),
.A2(n_1513),
.B(n_1502),
.Y(n_1639)
);

OR2x6_ASAP7_75t_L g1640 ( 
.A(n_1503),
.B(n_1532),
.Y(n_1640)
);

OAI211xp5_ASAP7_75t_L g1641 ( 
.A1(n_1513),
.A2(n_1579),
.B(n_1518),
.C(n_1594),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1565),
.A2(n_1513),
.B(n_1583),
.C(n_1510),
.Y(n_1642)
);

O2A1O1Ixp33_ASAP7_75t_L g1643 ( 
.A1(n_1595),
.A2(n_1513),
.B(n_1589),
.C(n_1585),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_R g1644 ( 
.A(n_1596),
.B(n_1593),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1503),
.B(n_1532),
.Y(n_1645)
);

AOI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1521),
.A2(n_1528),
.B1(n_1544),
.B2(n_1541),
.C(n_1539),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1590),
.B(n_1582),
.Y(n_1647)
);

AO32x2_ASAP7_75t_L g1648 ( 
.A1(n_1577),
.A2(n_1538),
.A3(n_1541),
.B1(n_1551),
.B2(n_1539),
.Y(n_1648)
);

O2A1O1Ixp33_ASAP7_75t_SL g1649 ( 
.A1(n_1592),
.A2(n_1595),
.B(n_1593),
.C(n_1535),
.Y(n_1649)
);

AO21x1_ASAP7_75t_L g1650 ( 
.A1(n_1575),
.A2(n_1580),
.B(n_1576),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1538),
.A2(n_1518),
.B(n_1571),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_SL g1652 ( 
.A(n_1640),
.B(n_1568),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1651),
.B(n_1518),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1651),
.B(n_1524),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1635),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1648),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1648),
.B(n_1524),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1648),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1637),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1637),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1611),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1640),
.B(n_1645),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1614),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1624),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1625),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1634),
.B(n_1524),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1641),
.B(n_1585),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1613),
.A2(n_1627),
.B1(n_1626),
.B2(n_1628),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1607),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1634),
.B(n_1524),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1615),
.A2(n_1593),
.B1(n_1591),
.B2(n_1586),
.Y(n_1671)
);

CKINVDCx20_ASAP7_75t_R g1672 ( 
.A(n_1610),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1639),
.B(n_1504),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1606),
.B(n_1534),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1606),
.B(n_1534),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1620),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1633),
.B(n_1530),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1612),
.Y(n_1678)
);

OAI221xp5_ASAP7_75t_SL g1679 ( 
.A1(n_1619),
.A2(n_1592),
.B1(n_1573),
.B2(n_1574),
.C(n_1498),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1632),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1650),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1620),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1620),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1646),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1682),
.B(n_1653),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1676),
.B(n_1641),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1657),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1676),
.B(n_1630),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1684),
.B(n_1642),
.C(n_1602),
.Y(n_1689)
);

NOR2x1_ASAP7_75t_L g1690 ( 
.A(n_1681),
.B(n_1599),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1661),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1672),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1657),
.Y(n_1693)
);

AOI33xp33_ASAP7_75t_L g1694 ( 
.A1(n_1684),
.A2(n_1628),
.A3(n_1619),
.B1(n_1633),
.B2(n_1616),
.B3(n_1643),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1653),
.B(n_1647),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1659),
.B(n_1623),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1652),
.B(n_1645),
.Y(n_1697)
);

OAI21xp33_ASAP7_75t_L g1698 ( 
.A1(n_1667),
.A2(n_1602),
.B(n_1631),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1653),
.B(n_1622),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1678),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1662),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1676),
.B(n_1683),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1668),
.A2(n_1617),
.B1(n_1618),
.B2(n_1599),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1676),
.B(n_1630),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1678),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1661),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1663),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1663),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1664),
.Y(n_1709)
);

OAI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1679),
.A2(n_1605),
.B1(n_1604),
.B2(n_1621),
.C(n_1643),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1652),
.B(n_1638),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1664),
.Y(n_1712)
);

NOR3xp33_ASAP7_75t_L g1713 ( 
.A(n_1679),
.B(n_1582),
.C(n_1589),
.Y(n_1713)
);

AND2x2_ASAP7_75t_SL g1714 ( 
.A(n_1662),
.B(n_1676),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1676),
.B(n_1621),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1683),
.B(n_1677),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1662),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1665),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1677),
.B(n_1656),
.Y(n_1719)
);

INVx5_ASAP7_75t_L g1720 ( 
.A(n_1681),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1681),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1667),
.A2(n_1608),
.B1(n_1629),
.B2(n_1636),
.Y(n_1722)
);

AOI33xp33_ASAP7_75t_L g1723 ( 
.A1(n_1655),
.A2(n_1609),
.A3(n_1649),
.B1(n_1598),
.B2(n_1600),
.B3(n_1603),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1687),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1702),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1691),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1720),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1685),
.B(n_1674),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1721),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1691),
.B(n_1660),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1685),
.B(n_1674),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1706),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1706),
.B(n_1660),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1707),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1707),
.B(n_1680),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1720),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1703),
.A2(n_1655),
.B1(n_1658),
.B2(n_1656),
.C(n_1666),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1708),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1702),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1708),
.B(n_1680),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1690),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1720),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1720),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1687),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1690),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1709),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1720),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1714),
.B(n_1675),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1709),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1714),
.B(n_1675),
.Y(n_1750)
);

NOR4xp25_ASAP7_75t_SL g1751 ( 
.A(n_1698),
.B(n_1636),
.C(n_1644),
.D(n_1610),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1712),
.B(n_1658),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1702),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1714),
.B(n_1675),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1719),
.B(n_1658),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1712),
.B(n_1673),
.Y(n_1756)
);

AND2x4_ASAP7_75t_SL g1757 ( 
.A(n_1711),
.B(n_1697),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1719),
.B(n_1669),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1718),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1719),
.B(n_1669),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1699),
.B(n_1666),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1715),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1718),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1693),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1726),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1758),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1757),
.B(n_1717),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1757),
.B(n_1717),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1729),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1757),
.B(n_1699),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1726),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1757),
.B(n_1720),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1758),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1758),
.B(n_1694),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1760),
.B(n_1723),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1760),
.B(n_1695),
.Y(n_1776)
);

INVxp67_ASAP7_75t_L g1777 ( 
.A(n_1729),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1726),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1737),
.A2(n_1698),
.B1(n_1689),
.B2(n_1703),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1760),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1732),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1730),
.B(n_1695),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1732),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1727),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1732),
.Y(n_1785)
);

NOR2x1p5_ASAP7_75t_L g1786 ( 
.A(n_1727),
.B(n_1692),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1730),
.B(n_1715),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1734),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1733),
.B(n_1695),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1733),
.B(n_1699),
.Y(n_1790)
);

NAND2x2_ASAP7_75t_L g1791 ( 
.A(n_1727),
.B(n_1692),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1737),
.A2(n_1689),
.B(n_1720),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1756),
.B(n_1715),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1762),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1734),
.Y(n_1795)
);

OAI21xp33_ASAP7_75t_SL g1796 ( 
.A1(n_1761),
.A2(n_1686),
.B(n_1716),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1727),
.B(n_1720),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1724),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1762),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1734),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1741),
.B(n_1721),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1741),
.B(n_1721),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1738),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1724),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1738),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1738),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1745),
.B(n_1696),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1745),
.B(n_1696),
.Y(n_1808)
);

INVx1_ASAP7_75t_SL g1809 ( 
.A(n_1736),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1761),
.B(n_1700),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1777),
.Y(n_1811)
);

INVxp67_ASAP7_75t_SL g1812 ( 
.A(n_1792),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1769),
.B(n_1761),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1774),
.B(n_1716),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1810),
.B(n_1748),
.Y(n_1815)
);

NAND4xp25_ASAP7_75t_L g1816 ( 
.A(n_1779),
.B(n_1686),
.C(n_1736),
.D(n_1692),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1810),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1786),
.B(n_1736),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1775),
.B(n_1716),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1782),
.B(n_1756),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1807),
.B(n_1686),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1770),
.B(n_1748),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1789),
.B(n_1752),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1784),
.Y(n_1824)
);

NOR2x1_ASAP7_75t_SL g1825 ( 
.A(n_1767),
.B(n_1742),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1798),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1798),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1765),
.Y(n_1828)
);

OR2x6_ASAP7_75t_L g1829 ( 
.A(n_1797),
.B(n_1742),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1808),
.B(n_1688),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_SL g1831 ( 
.A1(n_1796),
.A2(n_1666),
.B1(n_1710),
.B2(n_1654),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1765),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1809),
.B(n_1610),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1794),
.B(n_1688),
.Y(n_1834)
);

OAI21xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1772),
.A2(n_1743),
.B(n_1742),
.Y(n_1835)
);

INVxp33_ASAP7_75t_L g1836 ( 
.A(n_1767),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1799),
.B(n_1790),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1778),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1770),
.B(n_1748),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1804),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1766),
.B(n_1752),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1766),
.B(n_1688),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1778),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1772),
.B(n_1750),
.Y(n_1844)
);

INVx1_ASAP7_75t_SL g1845 ( 
.A(n_1801),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1784),
.B(n_1588),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1773),
.B(n_1704),
.Y(n_1847)
);

AOI21xp33_ASAP7_75t_L g1848 ( 
.A1(n_1812),
.A2(n_1802),
.B(n_1795),
.Y(n_1848)
);

INVxp67_ASAP7_75t_SL g1849 ( 
.A(n_1811),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1825),
.B(n_1772),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1828),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1828),
.Y(n_1852)
);

NAND2x1p5_ASAP7_75t_L g1853 ( 
.A(n_1824),
.B(n_1736),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1817),
.Y(n_1854)
);

NAND2xp33_ASAP7_75t_SL g1855 ( 
.A(n_1836),
.B(n_1751),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1845),
.B(n_1773),
.Y(n_1856)
);

OAI211xp5_ASAP7_75t_L g1857 ( 
.A1(n_1816),
.A2(n_1751),
.B(n_1743),
.C(n_1742),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1816),
.B(n_1846),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1825),
.B(n_1768),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1832),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1814),
.B(n_1780),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1817),
.Y(n_1862)
);

NOR4xp25_ASAP7_75t_SL g1863 ( 
.A(n_1835),
.B(n_1700),
.C(n_1705),
.D(n_1791),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1832),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1819),
.B(n_1780),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1831),
.A2(n_1791),
.B1(n_1776),
.B2(n_1710),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1820),
.B(n_1787),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1845),
.B(n_1755),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1815),
.B(n_1768),
.Y(n_1869)
);

AOI321xp33_ASAP7_75t_L g1870 ( 
.A1(n_1821),
.A2(n_1722),
.A3(n_1713),
.B1(n_1671),
.B2(n_1654),
.C(n_1670),
.Y(n_1870)
);

OAI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1813),
.A2(n_1722),
.B1(n_1704),
.B2(n_1701),
.Y(n_1871)
);

OAI322xp33_ASAP7_75t_L g1872 ( 
.A1(n_1837),
.A2(n_1787),
.A3(n_1704),
.B1(n_1793),
.B2(n_1803),
.C1(n_1800),
.C2(n_1795),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1815),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1818),
.B(n_1797),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1849),
.B(n_1824),
.Y(n_1875)
);

OAI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1870),
.A2(n_1835),
.B1(n_1830),
.B2(n_1834),
.C(n_1842),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1854),
.B(n_1862),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1873),
.B(n_1820),
.Y(n_1878)
);

OAI32xp33_ASAP7_75t_L g1879 ( 
.A1(n_1858),
.A2(n_1841),
.A3(n_1847),
.B1(n_1823),
.B2(n_1844),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1869),
.B(n_1833),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1869),
.B(n_1844),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1873),
.B(n_1823),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1852),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1852),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1854),
.B(n_1822),
.Y(n_1885)
);

OAI211xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1848),
.A2(n_1843),
.B(n_1838),
.C(n_1747),
.Y(n_1886)
);

AOI21xp33_ASAP7_75t_L g1887 ( 
.A1(n_1864),
.A2(n_1843),
.B(n_1838),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1864),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1862),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1871),
.A2(n_1840),
.B1(n_1826),
.B2(n_1827),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1866),
.A2(n_1818),
.B(n_1797),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1874),
.Y(n_1892)
);

AOI32xp33_ASAP7_75t_L g1893 ( 
.A1(n_1855),
.A2(n_1868),
.A3(n_1856),
.B1(n_1859),
.B2(n_1850),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1874),
.B(n_1822),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1855),
.A2(n_1857),
.B(n_1853),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1881),
.B(n_1859),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1892),
.B(n_1867),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1895),
.B(n_1818),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1875),
.B(n_1867),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1885),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1894),
.B(n_1861),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1877),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1878),
.B(n_1861),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1882),
.Y(n_1904)
);

AOI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1876),
.A2(n_1826),
.B1(n_1827),
.B2(n_1840),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1889),
.B(n_1880),
.Y(n_1906)
);

A2O1A1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1893),
.A2(n_1850),
.B(n_1860),
.C(n_1851),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1877),
.B(n_1865),
.Y(n_1908)
);

AOI32xp33_ASAP7_75t_L g1909 ( 
.A1(n_1899),
.A2(n_1886),
.A3(n_1883),
.B1(n_1884),
.B2(n_1888),
.Y(n_1909)
);

AOI32xp33_ASAP7_75t_L g1910 ( 
.A1(n_1904),
.A2(n_1895),
.A3(n_1879),
.B1(n_1818),
.B2(n_1865),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1898),
.A2(n_1863),
.B(n_1887),
.Y(n_1911)
);

NOR3xp33_ASAP7_75t_L g1912 ( 
.A(n_1902),
.B(n_1891),
.C(n_1887),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1903),
.Y(n_1913)
);

O2A1O1Ixp5_ASAP7_75t_L g1914 ( 
.A1(n_1907),
.A2(n_1872),
.B(n_1839),
.C(n_1853),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1896),
.B(n_1890),
.Y(n_1915)
);

INVxp67_ASAP7_75t_SL g1916 ( 
.A(n_1897),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1901),
.B(n_1853),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_SL g1918 ( 
.A1(n_1906),
.A2(n_1498),
.B(n_1829),
.Y(n_1918)
);

NOR2x1_ASAP7_75t_L g1919 ( 
.A(n_1908),
.B(n_1829),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1916),
.B(n_1902),
.Y(n_1920)
);

AOI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1914),
.A2(n_1905),
.B1(n_1900),
.B2(n_1804),
.C(n_1841),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1911),
.A2(n_1755),
.B1(n_1805),
.B2(n_1803),
.C(n_1800),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1913),
.Y(n_1923)
);

AOI222xp33_ASAP7_75t_L g1924 ( 
.A1(n_1915),
.A2(n_1919),
.B1(n_1917),
.B2(n_1912),
.C1(n_1910),
.C2(n_1909),
.Y(n_1924)
);

OAI22xp33_ASAP7_75t_L g1925 ( 
.A1(n_1918),
.A2(n_1829),
.B1(n_1743),
.B2(n_1747),
.Y(n_1925)
);

AOI211x1_ASAP7_75t_SL g1926 ( 
.A1(n_1911),
.A2(n_1829),
.B(n_1740),
.C(n_1735),
.Y(n_1926)
);

BUFx10_ASAP7_75t_L g1927 ( 
.A(n_1923),
.Y(n_1927)
);

O2A1O1Ixp33_ASAP7_75t_L g1928 ( 
.A1(n_1924),
.A2(n_1829),
.B(n_1839),
.C(n_1743),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1920),
.Y(n_1929)
);

OA22x2_ASAP7_75t_L g1930 ( 
.A1(n_1926),
.A2(n_1747),
.B1(n_1601),
.B2(n_1788),
.Y(n_1930)
);

AOI21xp33_ASAP7_75t_L g1931 ( 
.A1(n_1922),
.A2(n_1747),
.B(n_1788),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1921),
.A2(n_1805),
.B1(n_1705),
.B2(n_1806),
.C(n_1771),
.Y(n_1932)
);

OAI211xp5_ASAP7_75t_L g1933 ( 
.A1(n_1925),
.A2(n_1725),
.B(n_1753),
.C(n_1739),
.Y(n_1933)
);

AOI211xp5_ASAP7_75t_L g1934 ( 
.A1(n_1921),
.A2(n_1750),
.B(n_1754),
.C(n_1644),
.Y(n_1934)
);

AOI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1922),
.A2(n_1755),
.B1(n_1785),
.B2(n_1783),
.C(n_1781),
.Y(n_1935)
);

NAND4xp75_ASAP7_75t_L g1936 ( 
.A(n_1929),
.B(n_1750),
.C(n_1754),
.D(n_1728),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1927),
.Y(n_1937)
);

NAND4xp75_ASAP7_75t_L g1938 ( 
.A(n_1932),
.B(n_1931),
.C(n_1935),
.D(n_1928),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1930),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1933),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1934),
.B(n_1725),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1937),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1939),
.A2(n_1713),
.B1(n_1744),
.B2(n_1764),
.Y(n_1943)
);

OR3x1_ASAP7_75t_L g1944 ( 
.A(n_1937),
.B(n_1749),
.C(n_1746),
.Y(n_1944)
);

A2O1A1Ixp33_ASAP7_75t_L g1945 ( 
.A1(n_1942),
.A2(n_1940),
.B(n_1941),
.C(n_1938),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_SL g1946 ( 
.A1(n_1945),
.A2(n_1944),
.B1(n_1943),
.B2(n_1936),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1946),
.Y(n_1947)
);

INVxp33_ASAP7_75t_SL g1948 ( 
.A(n_1946),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1947),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1948),
.Y(n_1950)
);

OAI21xp33_ASAP7_75t_L g1951 ( 
.A1(n_1950),
.A2(n_1753),
.B(n_1739),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1949),
.B(n_1793),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1952),
.Y(n_1953)
);

OAI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1953),
.A2(n_1951),
.B(n_1731),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1954),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1955),
.A2(n_1746),
.B1(n_1749),
.B2(n_1763),
.C(n_1759),
.Y(n_1956)
);

AOI211xp5_ASAP7_75t_L g1957 ( 
.A1(n_1956),
.A2(n_1584),
.B(n_1591),
.C(n_1586),
.Y(n_1957)
);


endmodule