module fake_jpeg_8380_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_48),
.Y(n_57)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_18),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_37),
.A2(n_24),
.B1(n_19),
.B2(n_31),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_19),
.B1(n_43),
.B2(n_49),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_78),
.Y(n_128)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_80),
.B(n_81),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_83),
.Y(n_120)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_31),
.B(n_39),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_97),
.B(n_29),
.Y(n_126)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_87),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_108),
.B1(n_114),
.B2(n_69),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_91),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_93),
.B(n_44),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_94),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_44),
.C(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_57),
.B(n_50),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_44),
.C(n_42),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_49),
.A2(n_19),
.B1(n_30),
.B2(n_17),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_105),
.B1(n_116),
.B2(n_35),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_57),
.B(n_60),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_106),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_59),
.A2(n_30),
.B1(n_35),
.B2(n_21),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_59),
.Y(n_106)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_33),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_18),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_16),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_28),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_68),
.A2(n_17),
.B1(n_21),
.B2(n_28),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_26),
.A3(n_18),
.B1(n_20),
.B2(n_42),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_125),
.B1(n_130),
.B2(n_114),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_104),
.B(n_32),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_138),
.B(n_92),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_131),
.B(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_36),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_137),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_86),
.A2(n_36),
.B(n_69),
.C(n_29),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_116),
.B(n_93),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_36),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_32),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_71),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_147),
.B(n_150),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_107),
.B1(n_108),
.B2(n_113),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_151),
.B1(n_157),
.B2(n_163),
.Y(n_186)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_107),
.B1(n_76),
.B2(n_79),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_152),
.B(n_153),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_115),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_155),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_156),
.A2(n_161),
.B(n_170),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_91),
.B1(n_87),
.B2(n_98),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_93),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_139),
.B(n_124),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_84),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_165),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_127),
.B1(n_137),
.B2(n_126),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_110),
.B(n_90),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_122),
.B(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_167),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_78),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_172),
.B(n_175),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_85),
.B1(n_82),
.B2(n_80),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_177),
.B1(n_144),
.B2(n_120),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_122),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_20),
.Y(n_173)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_125),
.A2(n_45),
.B1(n_94),
.B2(n_20),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_124),
.B(n_18),
.Y(n_178)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_45),
.C(n_99),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_143),
.C(n_141),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_190),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_183),
.B(n_7),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_203),
.C(n_204),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_121),
.B1(n_141),
.B2(n_143),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_187),
.A2(n_188),
.B1(n_206),
.B2(n_7),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_120),
.B1(n_144),
.B2(n_136),
.Y(n_188)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_205),
.B1(n_152),
.B2(n_159),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_168),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_198),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_195),
.B(n_197),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_135),
.B(n_20),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_154),
.B(n_136),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_0),
.B(n_1),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_211),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_118),
.C(n_1),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_118),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_179),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_1),
.C(n_4),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_177),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_212),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_196),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_214),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_174),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_148),
.B(n_150),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_220),
.B(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_147),
.B1(n_156),
.B2(n_151),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_232),
.B1(n_206),
.B2(n_187),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_210),
.A2(n_172),
.B1(n_171),
.B2(n_164),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_166),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_6),
.Y(n_229)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_186),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_235),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_180),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_238),
.B(n_240),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_207),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_239),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_11),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_189),
.C(n_184),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_248),
.C(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_204),
.C(n_208),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_197),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_252),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_195),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_251),
.B(n_263),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_191),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_181),
.C(n_193),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_181),
.C(n_193),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_260),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_219),
.A2(n_188),
.B1(n_183),
.B2(n_201),
.Y(n_259)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_211),
.C(n_12),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_11),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_228),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_264),
.Y(n_292)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_252),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_265),
.B(n_236),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_242),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_231),
.B1(n_238),
.B2(n_232),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_213),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_247),
.B(n_257),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_276),
.B(n_280),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_216),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_278),
.Y(n_296)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_279),
.A2(n_281),
.B1(n_261),
.B2(n_229),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_237),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_222),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_282),
.A2(n_253),
.B1(n_226),
.B2(n_258),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_283),
.B(n_260),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_284),
.B(n_289),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_241),
.B(n_216),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_288),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_264),
.B(n_265),
.C(n_241),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_287),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_259),
.B(n_245),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_243),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_297),
.C(n_275),
.Y(n_302)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_215),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_248),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_295),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_263),
.C(n_236),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_266),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_297),
.C(n_272),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_299),
.C(n_300),
.Y(n_319)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_267),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_307),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_270),
.Y(n_305)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_308),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_275),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_11),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_289),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_287),
.B1(n_295),
.B2(n_285),
.Y(n_311)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_314),
.C(n_319),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_310),
.A2(n_286),
.B(n_290),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_298),
.Y(n_320)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_320),
.Y(n_327)
);

NOR2x1_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_304),
.Y(n_321)
);

NOR4xp25_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_316),
.C(n_317),
.D(n_313),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_298),
.C(n_299),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_272),
.C(n_14),
.Y(n_325)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_322),
.B(n_323),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_329),
.Y(n_332)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_330),
.B(n_327),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_15),
.B(n_12),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_14),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_15),
.Y(n_336)
);


endmodule