module fake_netlist_1_8602_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_10;
wire n_7;
AND2x4_ASAP7_75t_L g3 ( .A(n_1), .B(n_0), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
NOR2xp33_ASAP7_75t_L g5 ( .A(n_2), .B(n_1), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
NOR2x1_ASAP7_75t_SL g7 ( .A(n_4), .B(n_0), .Y(n_7) );
OA21x2_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_0), .B(n_2), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
OR2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_3), .Y(n_11) );
AOI221xp5_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_5), .B1(n_6), .B2(n_7), .C(n_0), .Y(n_12) );
O2A1O1Ixp33_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_9), .B(n_8), .C(n_7), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
AOI222xp33_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_2), .B1(n_8), .B2(n_9), .C1(n_11), .C2(n_12), .Y(n_15) );
endmodule