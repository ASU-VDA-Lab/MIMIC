module fake_netlist_1_12581_n_709 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_709);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_709;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_83), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_23), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_97), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_67), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_15), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_68), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_85), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_36), .Y(n_105) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_80), .B(n_62), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_55), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_93), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_17), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_3), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_74), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_21), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_89), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_69), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_92), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_78), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_48), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_56), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_66), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_1), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_61), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_3), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
BUFx10_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_38), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_27), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_86), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_54), .Y(n_130) );
BUFx3_ASAP7_75t_L g131 ( .A(n_17), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_37), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_70), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_84), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_4), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_16), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_52), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_95), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_71), .Y(n_139) );
INVxp67_ASAP7_75t_L g140 ( .A(n_47), .Y(n_140) );
INVx1_ASAP7_75t_SL g141 ( .A(n_82), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_28), .Y(n_142) );
BUFx8_ASAP7_75t_SL g143 ( .A(n_53), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_104), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g145 ( .A1(n_102), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_109), .B(n_0), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_108), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_131), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_108), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_128), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_131), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_128), .Y(n_152) );
INVx5_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_133), .A2(n_43), .B(n_94), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_109), .B(n_2), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_125), .B(n_4), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_104), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_136), .B(n_5), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_118), .B(n_5), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_163), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_163), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_163), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_153), .B(n_100), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_153), .B(n_112), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_163), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_156), .A2(n_123), .B1(n_102), .B2(n_101), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_163), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_153), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_163), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_147), .B(n_116), .Y(n_176) );
AND2x2_ASAP7_75t_L g177 ( .A(n_148), .B(n_135), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_147), .A2(n_135), .B1(n_111), .B2(n_136), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_158), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_158), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_153), .B(n_117), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
INVx5_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_149), .A2(n_127), .B1(n_142), .B2(n_132), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_189), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_184), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_177), .B(n_153), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_177), .B(n_153), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_184), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_177), .B(n_157), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_190), .A2(n_159), .B1(n_156), .B2(n_150), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_186), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_186), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_180), .A2(n_150), .B1(n_149), .B2(n_152), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_190), .A2(n_159), .B1(n_152), .B2(n_148), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_170), .A2(n_151), .B1(n_123), .B2(n_157), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_181), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_170), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_176), .B(n_157), .Y(n_205) );
NAND2xp33_ASAP7_75t_L g206 ( .A(n_188), .B(n_157), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_174), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_181), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_189), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_180), .A2(n_145), .B1(n_103), .B2(n_126), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_176), .B(n_151), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_174), .B(n_162), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_181), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_182), .Y(n_214) );
AO22x1_ASAP7_75t_L g215 ( .A1(n_185), .A2(n_114), .B1(n_105), .B2(n_107), .Y(n_215) );
INVxp67_ASAP7_75t_SL g216 ( .A(n_172), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_182), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_174), .B(n_146), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_167), .B(n_105), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_182), .Y(n_220) );
AOI221xp5_ASAP7_75t_L g221 ( .A1(n_174), .A2(n_145), .B1(n_155), .B2(n_146), .C(n_121), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_165), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_174), .A2(n_155), .B(n_161), .C(n_160), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_165), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_167), .B(n_124), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_208), .B(n_188), .Y(n_226) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_206), .A2(n_185), .B(n_168), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_202), .A2(n_98), .B1(n_137), .B2(n_168), .Y(n_228) );
AOI21x1_ASAP7_75t_L g229 ( .A1(n_215), .A2(n_185), .B(n_183), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_204), .B(n_175), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_196), .B(n_183), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_218), .A2(n_185), .B(n_154), .Y(n_232) );
OR2x6_ASAP7_75t_SL g233 ( .A(n_210), .B(n_107), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_218), .A2(n_188), .B(n_154), .Y(n_234) );
AO32x2_ASAP7_75t_L g235 ( .A1(n_200), .A2(n_188), .A3(n_160), .B1(n_175), .B2(n_179), .Y(n_235) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_222), .A2(n_178), .B(n_175), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_197), .B(n_175), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_192), .Y(n_238) );
INVx4_ASAP7_75t_L g239 ( .A(n_191), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_201), .A2(n_175), .B1(n_178), .B2(n_187), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_208), .B(n_188), .Y(n_241) );
BUFx12f_ASAP7_75t_L g242 ( .A(n_191), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_211), .B(n_172), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_205), .A2(n_188), .B(n_172), .Y(n_244) );
BUFx2_ASAP7_75t_L g245 ( .A(n_193), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_193), .B(n_178), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_205), .A2(n_188), .B(n_172), .Y(n_248) );
OAI21xp33_ASAP7_75t_L g249 ( .A1(n_194), .A2(n_113), .B(n_110), .Y(n_249) );
NAND3xp33_ASAP7_75t_L g250 ( .A(n_221), .B(n_188), .C(n_172), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_192), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_208), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_220), .B(n_189), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_194), .B(n_178), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_219), .B(n_178), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_213), .A2(n_166), .B(n_173), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_238), .A2(n_203), .B(n_214), .C(n_217), .Y(n_257) );
NOR2x1_ASAP7_75t_SL g258 ( .A(n_242), .B(n_200), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_237), .A2(n_210), .B(n_223), .C(n_221), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_242), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_226), .A2(n_213), .B(n_216), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_228), .B(n_212), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_226), .A2(n_214), .B(n_203), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_234), .A2(n_198), .B(n_199), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_233), .A2(n_198), .B1(n_195), .B2(n_199), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_251), .B(n_195), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_230), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_241), .A2(n_217), .B(n_199), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_241), .A2(n_198), .B(n_195), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_236), .A2(n_212), .B(n_220), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_245), .B(n_207), .Y(n_271) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_244), .A2(n_248), .A3(n_235), .B(n_240), .Y(n_272) );
INVxp67_ASAP7_75t_SL g273 ( .A(n_246), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_249), .B(n_225), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_232), .A2(n_220), .B(n_215), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_239), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_250), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_252), .B(n_207), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_227), .A2(n_222), .B(n_224), .Y(n_279) );
NAND2x1p5_ASAP7_75t_L g280 ( .A(n_239), .B(n_207), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_246), .B(n_207), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_266), .Y(n_282) );
AO31x2_ASAP7_75t_L g283 ( .A1(n_277), .A2(n_235), .A3(n_252), .B(n_231), .Y(n_283) );
AO221x1_ASAP7_75t_L g284 ( .A1(n_265), .A2(n_140), .B1(n_130), .B2(n_235), .C(n_120), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g285 ( .A(n_281), .B(n_253), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_259), .B(n_231), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_275), .A2(n_229), .B(n_235), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_264), .A2(n_256), .B(n_247), .Y(n_289) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_264), .A2(n_254), .B(n_139), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_280), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_279), .A2(n_253), .B(n_169), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_267), .B(n_243), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_265), .A2(n_243), .B1(n_255), .B2(n_179), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_279), .A2(n_119), .B(n_122), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_270), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_272), .Y(n_297) );
AO31x2_ASAP7_75t_L g298 ( .A1(n_258), .A2(n_255), .A3(n_165), .B(n_169), .Y(n_298) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_269), .A2(n_165), .B(n_169), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_262), .B(n_179), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g301 ( .A1(n_274), .A2(n_187), .B(n_179), .C(n_106), .Y(n_301) );
NAND4xp25_ASAP7_75t_L g302 ( .A(n_271), .B(n_179), .C(n_187), .D(n_141), .Y(n_302) );
AO31x2_ASAP7_75t_L g303 ( .A1(n_268), .A2(n_169), .A3(n_166), .B(n_171), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_288), .B(n_260), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_288), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_282), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_284), .A2(n_257), .B(n_263), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_296), .Y(n_311) );
OR2x6_ASAP7_75t_L g312 ( .A(n_291), .B(n_280), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_290), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_291), .B(n_278), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_291), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_290), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_290), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_291), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_297), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_299), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_302), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_283), .Y(n_327) );
AOI21x1_ASAP7_75t_L g328 ( .A1(n_287), .A2(n_261), .B(n_173), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
OA21x2_ASAP7_75t_L g330 ( .A1(n_292), .A2(n_273), .B(n_171), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_309), .B(n_283), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_322), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_309), .B(n_283), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_307), .B(n_286), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_316), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_319), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_319), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_322), .B(n_298), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_313), .B(n_283), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_320), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_307), .B(n_286), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_323), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_324), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_320), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_316), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_308), .B(n_283), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_316), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_323), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_308), .B(n_283), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_313), .B(n_302), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_315), .B(n_287), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
NAND2x1p5_ASAP7_75t_SL g353 ( .A(n_314), .B(n_284), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_327), .B(n_287), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_324), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_327), .B(n_287), .Y(n_356) );
NOR2x1p5_ASAP7_75t_L g357 ( .A(n_305), .B(n_300), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_305), .Y(n_358) );
INVx2_ASAP7_75t_R g359 ( .A(n_328), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_306), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_306), .B(n_287), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_326), .B(n_300), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_311), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_325), .B(n_295), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_311), .B(n_295), .Y(n_365) );
BUFx12f_ASAP7_75t_L g366 ( .A(n_312), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_311), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_304), .A2(n_293), .B1(n_294), .B2(n_295), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_317), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_321), .B(n_293), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_317), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_312), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_325), .B(n_295), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_352), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_337), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_338), .B(n_329), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_337), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_362), .B(n_314), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_358), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_331), .B(n_318), .Y(n_381) );
NOR2x1_ASAP7_75t_SL g382 ( .A(n_366), .B(n_312), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_340), .B(n_318), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_332), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_331), .B(n_318), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_331), .B(n_329), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_332), .Y(n_388) );
INVxp33_ASAP7_75t_L g389 ( .A(n_370), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_362), .B(n_295), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_342), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_338), .B(n_301), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_342), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_366), .B(n_143), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_366), .B(n_6), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_352), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_338), .B(n_298), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_333), .B(n_330), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_333), .B(n_330), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_352), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_348), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_348), .Y(n_402) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_335), .B(n_330), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_352), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_333), .B(n_330), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g406 ( .A(n_350), .B(n_187), .C(n_271), .D(n_281), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_358), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_336), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_354), .B(n_328), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_370), .B(n_298), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_354), .B(n_298), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_338), .B(n_298), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_355), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_354), .B(n_310), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_360), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_340), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_356), .B(n_310), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_338), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_344), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_356), .B(n_310), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_336), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_356), .B(n_303), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_334), .B(n_312), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_344), .B(n_303), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_336), .B(n_312), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_351), .B(n_303), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_344), .B(n_303), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_357), .A2(n_285), .B1(n_276), .B2(n_289), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_334), .B(n_272), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_341), .B(n_272), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_351), .B(n_303), .Y(n_432) );
NOR2xp33_ASAP7_75t_SL g433 ( .A(n_335), .B(n_285), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_360), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_335), .B(n_292), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_351), .B(n_303), .Y(n_436) );
OR2x6_ASAP7_75t_L g437 ( .A(n_373), .B(n_345), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_369), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_363), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_369), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_376), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_389), .B(n_345), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_426), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_384), .B(n_346), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_386), .B(n_345), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_378), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_384), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_388), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_419), .B(n_347), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_386), .B(n_350), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_381), .B(n_347), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_395), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_381), .B(n_347), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_388), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_379), .B(n_350), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_394), .B(n_6), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_419), .B(n_373), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_420), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_420), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_385), .B(n_339), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_391), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_391), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_383), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_383), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_385), .B(n_339), .Y(n_466) );
OAI332xp33_ASAP7_75t_L g467 ( .A1(n_411), .A2(n_341), .A3(n_349), .B1(n_346), .B2(n_339), .B3(n_365), .C1(n_12), .C2(n_13), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_419), .B(n_373), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_393), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_393), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_401), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_398), .B(n_349), .Y(n_472) );
AND3x2_ASAP7_75t_L g473 ( .A(n_433), .B(n_374), .C(n_364), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_401), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_426), .B(n_361), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_423), .B(n_361), .Y(n_476) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_403), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_439), .Y(n_478) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_403), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_402), .B(n_361), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_398), .B(n_343), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_399), .B(n_343), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_402), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_399), .B(n_343), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_405), .B(n_365), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_377), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_423), .B(n_364), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_427), .B(n_364), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_427), .B(n_374), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_407), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_405), .B(n_365), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_407), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_377), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_380), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_410), .B(n_374), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_410), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_426), .B(n_357), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_415), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_432), .B(n_363), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_432), .B(n_363), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_409), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_382), .B(n_367), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_436), .B(n_367), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_436), .B(n_367), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_408), .B(n_414), .Y(n_506) );
BUFx3_ASAP7_75t_L g507 ( .A(n_437), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_406), .A2(n_368), .B(n_372), .C(n_371), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_408), .B(n_371), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_414), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_416), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_382), .B(n_371), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_412), .B(n_372), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_412), .B(n_372), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_434), .B(n_368), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_438), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_377), .B(n_359), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_424), .B(n_7), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_425), .B(n_353), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_409), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_438), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_415), .B(n_359), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_441), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_445), .B(n_397), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_441), .B(n_418), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_506), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_476), .B(n_397), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_472), .B(n_418), .Y(n_528) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_503), .B(n_404), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_497), .B(n_421), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_508), .A2(n_479), .B(n_477), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_486), .B(n_425), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_497), .B(n_421), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_482), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_518), .A2(n_397), .B1(n_413), .B2(n_392), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_519), .A2(n_413), .B1(n_435), .B2(n_429), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_492), .B(n_428), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_465), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_455), .B(n_430), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_451), .B(n_413), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_456), .A2(n_431), .B1(n_390), .B2(n_437), .C(n_404), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_483), .Y(n_542) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_503), .B(n_440), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_496), .B(n_440), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_515), .B(n_422), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_498), .A2(n_435), .B1(n_422), .B2(n_375), .Y(n_547) );
O2A1O1Ixp5_ASAP7_75t_L g548 ( .A1(n_512), .A2(n_387), .B(n_375), .C(n_400), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_453), .B(n_435), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_495), .Y(n_550) );
INVxp33_ASAP7_75t_L g551 ( .A(n_442), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_460), .B(n_387), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_488), .B(n_396), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_489), .B(n_396), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_446), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_515), .B(n_400), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_485), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_490), .B(n_403), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_466), .B(n_359), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_502), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_458), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_496), .B(n_359), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_512), .B(n_353), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_447), .Y(n_564) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_507), .A2(n_353), .B1(n_285), .B2(n_299), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_463), .B(n_292), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_452), .B(n_7), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_450), .B(n_8), .Y(n_568) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_459), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_502), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_458), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_473), .B(n_289), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_463), .B(n_299), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_448), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_464), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_520), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_444), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_464), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_454), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_501), .B(n_9), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_475), .B(n_299), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_501), .B(n_9), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_449), .Y(n_583) );
NAND2xp33_ASAP7_75t_SL g584 ( .A(n_498), .B(n_115), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_505), .B(n_10), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_444), .B(n_10), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_461), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_505), .B(n_11), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_443), .A2(n_468), .B1(n_457), .B2(n_499), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_459), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_462), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_480), .B(n_11), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_469), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_470), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_480), .B(n_12), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_471), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_499), .B(n_115), .C(n_129), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_516), .B(n_13), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_541), .A2(n_467), .B1(n_484), .B2(n_491), .C(n_493), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_577), .B(n_500), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_523), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_531), .A2(n_509), .B(n_449), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_578), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_538), .B(n_504), .Y(n_604) );
OAI21xp33_ASAP7_75t_L g605 ( .A1(n_536), .A2(n_522), .B(n_475), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_567), .B(n_510), .C(n_511), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_527), .B(n_513), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_551), .B(n_457), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_526), .B(n_514), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_578), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_543), .A2(n_517), .B(n_521), .Y(n_611) );
AND3x1_ASAP7_75t_L g612 ( .A(n_563), .B(n_473), .C(n_494), .Y(n_612) );
OAI21xp33_ASAP7_75t_SL g613 ( .A1(n_531), .A2(n_509), .B(n_474), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_583), .B(n_487), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_590), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_572), .A2(n_481), .B(n_478), .Y(n_616) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_589), .A2(n_138), .B(n_134), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_572), .A2(n_289), .B(n_138), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_548), .B(n_129), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_535), .A2(n_134), .B1(n_187), .B2(n_164), .Y(n_620) );
AOI21xp33_ASAP7_75t_SL g621 ( .A1(n_529), .A2(n_14), .B(n_15), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_544), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_569), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_550), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_568), .B(n_14), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_539), .A2(n_164), .B1(n_18), .B2(n_19), .Y(n_626) );
OAI21xp33_ASAP7_75t_SL g627 ( .A1(n_558), .A2(n_16), .B(n_18), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_553), .B(n_19), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_554), .B(n_20), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_565), .A2(n_20), .B(n_21), .Y(n_630) );
BUFx2_ASAP7_75t_L g631 ( .A(n_576), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_545), .B(n_22), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_560), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_529), .A2(n_164), .B1(n_25), .B2(n_26), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_545), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_525), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_525), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_530), .A2(n_164), .B1(n_224), .B2(n_222), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_555), .B(n_24), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_564), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_584), .A2(n_164), .B1(n_30), .B2(n_31), .C(n_32), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_574), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_570), .Y(n_643) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_532), .A2(n_164), .B1(n_33), .B2(n_34), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_530), .A2(n_224), .B1(n_35), .B2(n_39), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_573), .A2(n_29), .B(n_40), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_635), .B(n_546), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_636), .B(n_556), .Y(n_648) );
AOI221x1_ASAP7_75t_SL g649 ( .A1(n_605), .A2(n_595), .B1(n_592), .B2(n_586), .C(n_598), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_613), .A2(n_533), .B1(n_592), .B2(n_595), .C(n_528), .Y(n_650) );
AOI32xp33_ASAP7_75t_L g651 ( .A1(n_612), .A2(n_540), .A3(n_524), .B1(n_549), .B2(n_575), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_637), .B(n_528), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_608), .B(n_557), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_633), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_606), .A2(n_533), .B1(n_547), .B2(n_562), .Y(n_655) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_623), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_602), .A2(n_537), .B1(n_580), .B2(n_582), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_599), .B(n_588), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_602), .B(n_571), .Y(n_659) );
AOI332xp33_ASAP7_75t_L g660 ( .A1(n_622), .A2(n_593), .A3(n_587), .B1(n_596), .B2(n_594), .B3(n_579), .C1(n_591), .C2(n_542), .Y(n_660) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_619), .Y(n_661) );
NAND3xp33_ASAP7_75t_SL g662 ( .A(n_621), .B(n_585), .C(n_597), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_627), .A2(n_534), .B1(n_581), .B2(n_561), .Y(n_663) );
OAI21xp33_ASAP7_75t_SL g664 ( .A1(n_611), .A2(n_598), .B(n_559), .Y(n_664) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_599), .A2(n_566), .B1(n_552), .B2(n_44), .C1(n_45), .C2(n_46), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_640), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_603), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_631), .A2(n_41), .B1(n_42), .B2(n_49), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_625), .A2(n_50), .B1(n_51), .B2(n_57), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_610), .Y(n_670) );
OAI22xp5_ASAP7_75t_SL g671 ( .A1(n_615), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_671) );
OAI222xp33_ASAP7_75t_L g672 ( .A1(n_616), .A2(n_63), .B1(n_64), .B2(n_65), .C1(n_72), .C2(n_73), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g673 ( .A1(n_617), .A2(n_76), .B(n_79), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g674 ( .A1(n_618), .A2(n_87), .B(n_88), .C(n_90), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_630), .B(n_91), .C(n_96), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_630), .A2(n_209), .B(n_189), .C(n_191), .Y(n_676) );
AOI21xp33_ASAP7_75t_SL g677 ( .A1(n_634), .A2(n_189), .B(n_209), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_601), .B(n_189), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_L g679 ( .A1(n_628), .A2(n_189), .B(n_629), .C(n_643), .Y(n_679) );
AOI221x1_ASAP7_75t_SL g680 ( .A1(n_604), .A2(n_189), .B1(n_624), .B2(n_600), .C(n_609), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_646), .A2(n_644), .B(n_641), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_642), .A2(n_632), .B1(n_626), .B2(n_614), .C(n_646), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_639), .A2(n_620), .B(n_607), .Y(n_683) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_638), .B(n_599), .C(n_602), .D(n_630), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_645), .B(n_631), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_665), .B(n_684), .C(n_650), .Y(n_686) );
NOR3x1_ASAP7_75t_L g687 ( .A(n_658), .B(n_661), .C(n_656), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_667), .B(n_670), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_666), .Y(n_689) );
AOI211xp5_ASAP7_75t_SL g690 ( .A1(n_681), .A2(n_662), .B(n_685), .C(n_671), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_659), .A2(n_667), .B(n_677), .C(n_664), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_679), .A2(n_651), .B(n_676), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_686), .B(n_668), .C(n_672), .Y(n_693) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_691), .B(n_675), .C(n_674), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_692), .B(n_678), .C(n_673), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_688), .B(n_653), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_696), .B(n_689), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_693), .B(n_690), .Y(n_698) );
OAI22x1_ASAP7_75t_L g699 ( .A1(n_694), .A2(n_687), .B1(n_663), .B2(n_669), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_697), .Y(n_700) );
XNOR2xp5_ASAP7_75t_L g701 ( .A(n_698), .B(n_695), .Y(n_701) );
OA21x2_ASAP7_75t_L g702 ( .A1(n_701), .A2(n_699), .B(n_682), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_700), .Y(n_703) );
OA22x2_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_655), .B1(n_654), .B2(n_657), .Y(n_704) );
OAI22x1_ASAP7_75t_L g705 ( .A1(n_702), .A2(n_680), .B1(n_649), .B2(n_652), .Y(n_705) );
AOI222xp33_ASAP7_75t_L g706 ( .A1(n_705), .A2(n_702), .B1(n_647), .B2(n_648), .C1(n_649), .C2(n_660), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_706), .B(n_702), .Y(n_707) );
OR2x6_ASAP7_75t_L g708 ( .A(n_707), .B(n_704), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_702), .B(n_683), .Y(n_709) );
endmodule