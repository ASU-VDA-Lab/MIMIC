module real_aes_7200_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g180 ( .A1(n_0), .A2(n_181), .B(n_184), .C(n_188), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_1), .B(n_172), .Y(n_191) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_3), .B(n_182), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_4), .A2(n_141), .B(n_511), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_5), .A2(n_146), .B(n_149), .C(n_538), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_6), .A2(n_141), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_7), .B(n_172), .Y(n_517) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_8), .A2(n_174), .B(n_249), .Y(n_248) );
AND2x6_ASAP7_75t_L g146 ( .A(n_9), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_10), .A2(n_146), .B(n_149), .C(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g551 ( .A(n_11), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_12), .B(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_12), .B(n_43), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_13), .B(n_187), .Y(n_540) );
INVx1_ASAP7_75t_L g167 ( .A(n_14), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_15), .B(n_182), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_16), .A2(n_183), .B(n_571), .C(n_573), .Y(n_570) );
XOR2xp5_ASAP7_75t_L g124 ( .A(n_17), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_17), .B(n_172), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_18), .B(n_455), .Y(n_454) );
AOI222xp33_ASAP7_75t_SL g457 ( .A1(n_19), .A2(n_458), .B1(n_459), .B2(n_468), .C1(n_735), .C2(n_736), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_20), .B(n_161), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_21), .A2(n_149), .B(n_152), .C(n_160), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_22), .A2(n_186), .B(n_242), .C(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_23), .B(n_187), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_24), .A2(n_42), .B1(n_465), .B2(n_466), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_24), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_25), .B(n_187), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g485 ( .A(n_26), .Y(n_485) );
INVx1_ASAP7_75t_L g524 ( .A(n_27), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_28), .A2(n_149), .B(n_160), .C(n_252), .Y(n_251) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_29), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_30), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_31), .A2(n_79), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_31), .Y(n_130) );
INVx1_ASAP7_75t_L g502 ( .A(n_32), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_33), .A2(n_141), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g144 ( .A(n_34), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_35), .A2(n_200), .B(n_201), .C(n_205), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_36), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_37), .A2(n_186), .B(n_514), .C(n_516), .Y(n_513) );
INVxp67_ASAP7_75t_L g503 ( .A(n_38), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_39), .B(n_254), .Y(n_253) );
CKINVDCx14_ASAP7_75t_R g512 ( .A(n_40), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_41), .A2(n_149), .B(n_160), .C(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_42), .Y(n_465) );
INVx1_ASAP7_75t_L g117 ( .A(n_43), .Y(n_117) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_44), .A2(n_188), .B(n_549), .C(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_45), .B(n_140), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_46), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_47), .B(n_182), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_48), .B(n_141), .Y(n_250) );
OAI22xp5_ASAP7_75t_SL g459 ( .A1(n_49), .A2(n_460), .B1(n_461), .B2(n_467), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_49), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_50), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_51), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_52), .A2(n_200), .B(n_205), .C(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g185 ( .A(n_53), .Y(n_185) );
INVx1_ASAP7_75t_L g228 ( .A(n_54), .Y(n_228) );
INVx1_ASAP7_75t_L g557 ( .A(n_55), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_56), .B(n_141), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_57), .Y(n_169) );
CKINVDCx14_ASAP7_75t_R g547 ( .A(n_58), .Y(n_547) );
INVx1_ASAP7_75t_L g147 ( .A(n_59), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_60), .B(n_141), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_61), .B(n_172), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_62), .A2(n_159), .B(n_215), .C(n_217), .Y(n_214) );
INVx1_ASAP7_75t_L g166 ( .A(n_63), .Y(n_166) );
INVx1_ASAP7_75t_SL g515 ( .A(n_64), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_65), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_66), .B(n_182), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_67), .B(n_172), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_68), .B(n_183), .Y(n_239) );
INVx1_ASAP7_75t_L g488 ( .A(n_69), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_70), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_71), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_72), .A2(n_149), .B(n_205), .C(n_268), .Y(n_267) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_73), .Y(n_213) );
INVx1_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_75), .A2(n_141), .B(n_546), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_76), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_77), .A2(n_141), .B(n_568), .Y(n_567) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_78), .A2(n_127), .B1(n_128), .B2(n_131), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_78), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_79), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_80), .A2(n_140), .B(n_498), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_81), .Y(n_521) );
INVx1_ASAP7_75t_L g569 ( .A(n_82), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_83), .B(n_157), .Y(n_156) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_84), .A2(n_462), .B1(n_463), .B2(n_464), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_84), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_85), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_86), .A2(n_141), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g572 ( .A(n_87), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_88), .A2(n_105), .B1(n_106), .B2(n_118), .Y(n_104) );
INVx2_ASAP7_75t_L g164 ( .A(n_89), .Y(n_164) );
INVx1_ASAP7_75t_L g539 ( .A(n_90), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_91), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_92), .B(n_187), .Y(n_240) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_93), .B(n_111), .C(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g450 ( .A(n_93), .B(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g471 ( .A(n_93), .B(n_452), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_93), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_94), .A2(n_149), .B(n_205), .C(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_95), .B(n_141), .Y(n_198) );
INVx1_ASAP7_75t_L g202 ( .A(n_96), .Y(n_202) );
INVxp67_ASAP7_75t_L g218 ( .A(n_97), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_98), .B(n_174), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_99), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g235 ( .A(n_100), .Y(n_235) );
INVx1_ASAP7_75t_L g269 ( .A(n_101), .Y(n_269) );
INVx2_ASAP7_75t_L g560 ( .A(n_102), .Y(n_560) );
AND2x2_ASAP7_75t_L g230 ( .A(n_103), .B(n_163), .Y(n_230) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
BUFx4f_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_115), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g452 ( .A(n_111), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVxp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B(n_456), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g741 ( .A(n_122), .Y(n_741) );
OAI21xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_447), .B(n_454), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_132), .B1(n_445), .B2(n_446), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_126), .Y(n_445) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g446 ( .A(n_132), .Y(n_446) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_132), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_381), .Y(n_132) );
NOR5xp2_ASAP7_75t_L g133 ( .A(n_134), .B(n_312), .C(n_341), .D(n_361), .E(n_368), .Y(n_133) );
OAI211xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_192), .B(n_256), .C(n_299), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_136), .A2(n_384), .B1(n_386), .B2(n_387), .Y(n_383) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_171), .Y(n_136) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_137), .Y(n_259) );
AND2x4_ASAP7_75t_L g292 ( .A(n_137), .B(n_293), .Y(n_292) );
INVx5_ASAP7_75t_L g310 ( .A(n_137), .Y(n_310) );
AND2x2_ASAP7_75t_L g319 ( .A(n_137), .B(n_311), .Y(n_319) );
AND2x2_ASAP7_75t_L g331 ( .A(n_137), .B(n_196), .Y(n_331) );
AND2x2_ASAP7_75t_L g427 ( .A(n_137), .B(n_295), .Y(n_427) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_168), .Y(n_137) );
AOI21xp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_148), .B(n_161), .Y(n_138) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_142), .B(n_146), .Y(n_236) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g159 ( .A(n_143), .Y(n_159) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
INVx1_ASAP7_75t_L g243 ( .A(n_144), .Y(n_243) );
INVx1_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_145), .Y(n_155) );
INVx3_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx1_ASAP7_75t_L g254 ( .A(n_145), .Y(n_254) );
BUFx3_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
INVx4_ASAP7_75t_SL g190 ( .A(n_146), .Y(n_190) );
INVx5_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx3_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_150), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_156), .B(n_158), .Y(n_152) );
INVx2_ASAP7_75t_L g157 ( .A(n_154), .Y(n_157) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx4_ASAP7_75t_L g216 ( .A(n_155), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_157), .A2(n_202), .B(n_203), .C(n_204), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_157), .A2(n_204), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_157), .A2(n_488), .B(n_489), .C(n_490), .Y(n_487) );
O2A1O1Ixp5_ASAP7_75t_L g538 ( .A1(n_157), .A2(n_490), .B(n_539), .C(n_540), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_158), .A2(n_182), .B(n_524), .C(n_525), .Y(n_523) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_159), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_162), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g170 ( .A(n_163), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_163), .A2(n_198), .B(n_199), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_163), .A2(n_225), .B(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_163), .A2(n_236), .B(n_521), .C(n_522), .Y(n_520) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_163), .A2(n_545), .B(n_552), .Y(n_544) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_164), .B(n_165), .Y(n_163) );
AND2x2_ASAP7_75t_L g175 ( .A(n_164), .B(n_165), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_170), .A2(n_535), .B(n_541), .Y(n_534) );
INVx2_ASAP7_75t_L g293 ( .A(n_171), .Y(n_293) );
AND2x2_ASAP7_75t_L g311 ( .A(n_171), .B(n_265), .Y(n_311) );
AND2x2_ASAP7_75t_L g330 ( .A(n_171), .B(n_264), .Y(n_330) );
AND2x2_ASAP7_75t_L g370 ( .A(n_171), .B(n_310), .Y(n_370) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_176), .B(n_191), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_173), .B(n_207), .Y(n_206) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_173), .A2(n_234), .B(n_244), .Y(n_233) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_173), .A2(n_266), .B(n_274), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_173), .B(n_275), .Y(n_274) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_173), .A2(n_484), .B(n_491), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_173), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_173), .B(n_542), .Y(n_541) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_174), .A2(n_250), .B(n_251), .Y(n_249) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g246 ( .A(n_175), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_179), .B(n_180), .C(n_190), .Y(n_177) );
INVx2_ASAP7_75t_L g200 ( .A(n_179), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_179), .A2(n_190), .B(n_213), .C(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_179), .A2(n_190), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_179), .A2(n_190), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_SL g546 ( .A1(n_179), .A2(n_190), .B(n_547), .C(n_548), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_SL g556 ( .A1(n_179), .A2(n_190), .B(n_557), .C(n_558), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_SL g568 ( .A1(n_179), .A2(n_190), .B(n_569), .C(n_570), .Y(n_568) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_182), .B(n_218), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g501 ( .A1(n_182), .A2(n_216), .B1(n_502), .B2(n_503), .Y(n_501) );
INVx5_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_183), .B(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_186), .B(n_515), .Y(n_514) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g549 ( .A(n_187), .Y(n_549) );
INVx2_ASAP7_75t_L g490 ( .A(n_188), .Y(n_490) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_189), .Y(n_204) );
INVx1_ASAP7_75t_L g573 ( .A(n_189), .Y(n_573) );
INVx1_ASAP7_75t_L g205 ( .A(n_190), .Y(n_205) );
INVxp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_220), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI322xp5_ASAP7_75t_L g429 ( .A1(n_195), .A2(n_231), .A3(n_284), .B1(n_292), .B2(n_346), .C1(n_430), .C2(n_433), .Y(n_429) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_208), .Y(n_195) );
INVx5_ASAP7_75t_L g261 ( .A(n_196), .Y(n_261) );
AND2x2_ASAP7_75t_L g278 ( .A(n_196), .B(n_263), .Y(n_278) );
BUFx2_ASAP7_75t_L g356 ( .A(n_196), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_196), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g433 ( .A(n_196), .B(n_340), .Y(n_433) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_206), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_208), .B(n_222), .Y(n_287) );
INVx1_ASAP7_75t_L g314 ( .A(n_208), .Y(n_314) );
AND2x2_ASAP7_75t_L g327 ( .A(n_208), .B(n_247), .Y(n_327) );
AND2x2_ASAP7_75t_L g428 ( .A(n_208), .B(n_346), .Y(n_428) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g282 ( .A(n_209), .B(n_222), .Y(n_282) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_209), .Y(n_290) );
OR2x2_ASAP7_75t_L g297 ( .A(n_209), .B(n_247), .Y(n_297) );
AND2x2_ASAP7_75t_L g307 ( .A(n_209), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_209), .B(n_233), .Y(n_336) );
INVxp67_ASAP7_75t_L g360 ( .A(n_209), .Y(n_360) );
AND2x2_ASAP7_75t_L g367 ( .A(n_209), .B(n_231), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_209), .B(n_247), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_209), .B(n_232), .Y(n_393) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_219), .Y(n_209) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_210), .A2(n_510), .B(n_517), .Y(n_509) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_210), .A2(n_555), .B(n_561), .Y(n_554) );
OA21x2_ASAP7_75t_L g566 ( .A1(n_210), .A2(n_567), .B(n_574), .Y(n_566) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_215), .A2(n_269), .B(n_270), .C(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_216), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_216), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_231), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_222), .B(n_248), .Y(n_337) );
OR2x2_ASAP7_75t_L g359 ( .A(n_222), .B(n_232), .Y(n_359) );
AND2x2_ASAP7_75t_L g372 ( .A(n_222), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_222), .B(n_327), .Y(n_378) );
OAI211xp5_ASAP7_75t_SL g382 ( .A1(n_222), .A2(n_383), .B(n_388), .C(n_397), .Y(n_382) );
AND2x2_ASAP7_75t_L g443 ( .A(n_222), .B(n_247), .Y(n_443) );
INVx5_ASAP7_75t_SL g222 ( .A(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g296 ( .A(n_223), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_223), .B(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_223), .B(n_291), .Y(n_303) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_223), .Y(n_305) );
OR2x2_ASAP7_75t_L g316 ( .A(n_223), .B(n_232), .Y(n_316) );
AND2x2_ASAP7_75t_SL g321 ( .A(n_223), .B(n_307), .Y(n_321) );
AND2x2_ASAP7_75t_L g346 ( .A(n_223), .B(n_232), .Y(n_346) );
AND2x2_ASAP7_75t_L g366 ( .A(n_223), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g404 ( .A(n_223), .B(n_231), .Y(n_404) );
OR2x2_ASAP7_75t_L g407 ( .A(n_223), .B(n_393), .Y(n_407) );
OR2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_230), .Y(n_223) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_247), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_232), .A2(n_351), .B(n_354), .C(n_360), .Y(n_350) );
INVx5_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_233), .B(n_247), .Y(n_281) );
AND2x2_ASAP7_75t_L g285 ( .A(n_233), .B(n_248), .Y(n_285) );
OR2x2_ASAP7_75t_L g291 ( .A(n_233), .B(n_247), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_237), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_236), .A2(n_485), .B(n_486), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_236), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_241), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_241), .A2(n_253), .B(n_255), .Y(n_252) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g495 ( .A(n_246), .Y(n_495) );
INVx1_ASAP7_75t_SL g308 ( .A(n_247), .Y(n_308) );
OR2x2_ASAP7_75t_L g436 ( .A(n_247), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_276), .B(n_279), .C(n_288), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AOI31xp33_ASAP7_75t_L g361 ( .A1(n_258), .A2(n_362), .A3(n_364), .B(n_365), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_259), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_260), .B(n_292), .Y(n_298) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_261), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g318 ( .A(n_261), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g323 ( .A(n_261), .B(n_293), .Y(n_323) );
AND2x2_ASAP7_75t_L g333 ( .A(n_261), .B(n_292), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_261), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g353 ( .A(n_261), .B(n_310), .Y(n_353) );
AND2x2_ASAP7_75t_L g358 ( .A(n_261), .B(n_330), .Y(n_358) );
OR2x2_ASAP7_75t_L g377 ( .A(n_261), .B(n_263), .Y(n_377) );
OR2x2_ASAP7_75t_L g379 ( .A(n_261), .B(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_261), .Y(n_426) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g326 ( .A(n_263), .B(n_293), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_263), .B(n_310), .Y(n_349) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
BUFx2_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_273), .Y(n_266) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx3_ASAP7_75t_L g516 ( .A(n_272), .Y(n_516) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g386 ( .A(n_278), .B(n_310), .Y(n_386) );
AOI322xp5_ASAP7_75t_L g388 ( .A1(n_278), .A2(n_292), .A3(n_330), .B1(n_389), .B2(n_390), .C1(n_391), .C2(n_394), .Y(n_388) );
INVx1_ASAP7_75t_L g396 ( .A(n_278), .Y(n_396) );
NAND2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_SL g390 ( .A(n_280), .Y(n_390) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
OR2x2_ASAP7_75t_L g342 ( .A(n_281), .B(n_287), .Y(n_342) );
INVx1_ASAP7_75t_L g373 ( .A(n_281), .Y(n_373) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI32xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_292), .A3(n_294), .B1(n_296), .B2(n_298), .Y(n_288) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AOI21xp33_ASAP7_75t_SL g328 ( .A1(n_291), .A2(n_306), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g343 ( .A(n_292), .Y(n_343) );
AND2x4_ASAP7_75t_L g340 ( .A(n_293), .B(n_310), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_293), .B(n_376), .Y(n_375) );
AOI322xp5_ASAP7_75t_L g405 ( .A1(n_294), .A2(n_321), .A3(n_340), .B1(n_373), .B2(n_406), .C1(n_408), .C2(n_409), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_294), .A2(n_371), .B1(n_435), .B2(n_436), .C(n_438), .Y(n_434) );
AND2x2_ASAP7_75t_L g322 ( .A(n_295), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g302 ( .A(n_297), .Y(n_302) );
OR2x2_ASAP7_75t_L g374 ( .A(n_297), .B(n_359), .Y(n_374) );
OAI31xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .A3(n_304), .B(n_309), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_300), .A2(n_333), .B1(n_334), .B2(n_338), .Y(n_332) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g345 ( .A(n_302), .B(n_346), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_304), .A2(n_345), .B1(n_398), .B2(n_401), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g387 ( .A(n_307), .B(n_356), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_307), .B(n_346), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_308), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g421 ( .A(n_308), .B(n_359), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_309), .A2(n_404), .B1(n_417), .B2(n_420), .Y(n_416) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g325 ( .A(n_310), .Y(n_325) );
AND2x2_ASAP7_75t_L g408 ( .A(n_310), .B(n_330), .Y(n_408) );
OR2x2_ASAP7_75t_L g410 ( .A(n_310), .B(n_377), .Y(n_410) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_310), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_311), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_311), .B(n_356), .Y(n_364) );
OAI211xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_317), .B(n_320), .C(n_332), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B1(n_324), .B2(n_327), .C(n_328), .Y(n_320) );
INVxp67_ASAP7_75t_L g432 ( .A(n_323), .Y(n_432) );
INVx1_ASAP7_75t_L g399 ( .A(n_324), .Y(n_399) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g363 ( .A(n_325), .B(n_330), .Y(n_363) );
INVx1_ASAP7_75t_L g380 ( .A(n_326), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_326), .B(n_353), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g395 ( .A(n_330), .Y(n_395) );
AND2x2_ASAP7_75t_L g401 ( .A(n_330), .B(n_356), .Y(n_401) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_SL g389 ( .A(n_337), .Y(n_389) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_340), .B(n_376), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_344), .B2(n_347), .C(n_350), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g437 ( .A(n_346), .Y(n_437) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g355 ( .A(n_349), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_353), .B(n_412), .Y(n_411) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B(n_359), .Y(n_354) );
OAI211xp5_ASAP7_75t_SL g402 ( .A1(n_357), .A2(n_403), .B(n_405), .C(n_411), .Y(n_402) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g414 ( .A(n_359), .Y(n_414) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI222xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B1(n_374), .B2(n_375), .C1(n_378), .C2(n_379), .Y(n_368) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g444 ( .A(n_375), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_376), .B(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_376), .A2(n_423), .B1(n_425), .B2(n_428), .Y(n_422) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
NOR4xp25_ASAP7_75t_L g381 ( .A(n_382), .B(n_402), .C(n_415), .D(n_434), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_384), .B(n_414), .Y(n_424) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g391 ( .A(n_389), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_392), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_422), .C(n_429), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx2_ASAP7_75t_L g431 ( .A(n_427), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_441), .B(n_444), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_446), .A2(n_469), .B1(n_472), .B2(n_474), .Y(n_468) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g455 ( .A(n_450), .Y(n_455) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_451), .B(n_473), .Y(n_735) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g472 ( .A(n_452), .B(n_473), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_454), .B(n_457), .C(n_741), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g737 ( .A(n_470), .Y(n_737) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g740 ( .A(n_472), .Y(n_740) );
INVx2_ASAP7_75t_L g738 ( .A(n_474), .Y(n_738) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_669), .Y(n_474) );
NAND5xp2_ASAP7_75t_L g475 ( .A(n_476), .B(n_598), .C(n_628), .D(n_649), .E(n_655), .Y(n_475) );
AOI221xp5_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_531), .B1(n_562), .B2(n_564), .C(n_575), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_528), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_506), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_SL g649 ( .A1(n_481), .A2(n_518), .B(n_650), .C(n_653), .Y(n_649) );
AND2x2_ASAP7_75t_L g719 ( .A(n_481), .B(n_519), .Y(n_719) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_493), .Y(n_481) );
AND2x2_ASAP7_75t_L g577 ( .A(n_482), .B(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g581 ( .A(n_482), .B(n_578), .Y(n_581) );
OR2x2_ASAP7_75t_L g607 ( .A(n_482), .B(n_519), .Y(n_607) );
AND2x2_ASAP7_75t_L g609 ( .A(n_482), .B(n_509), .Y(n_609) );
AND2x2_ASAP7_75t_L g627 ( .A(n_482), .B(n_508), .Y(n_627) );
INVx1_ASAP7_75t_L g660 ( .A(n_482), .Y(n_660) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g530 ( .A(n_483), .Y(n_530) );
AND2x2_ASAP7_75t_L g563 ( .A(n_483), .B(n_509), .Y(n_563) );
AND2x2_ASAP7_75t_L g716 ( .A(n_483), .B(n_519), .Y(n_716) );
AND2x2_ASAP7_75t_L g597 ( .A(n_493), .B(n_507), .Y(n_597) );
OR2x2_ASAP7_75t_L g601 ( .A(n_493), .B(n_519), .Y(n_601) );
AND2x2_ASAP7_75t_L g626 ( .A(n_493), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g673 ( .A(n_493), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_493), .B(n_635), .Y(n_721) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B(n_504), .Y(n_493) );
INVx1_ASAP7_75t_L g579 ( .A(n_494), .Y(n_579) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OA21x2_ASAP7_75t_L g578 ( .A1(n_497), .A2(n_505), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OAI322xp33_ASAP7_75t_L g722 ( .A1(n_506), .A2(n_658), .A3(n_681), .B1(n_702), .B2(n_723), .C1(n_725), .C2(n_726), .Y(n_722) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_507), .B(n_578), .Y(n_725) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .Y(n_507) );
AND2x2_ASAP7_75t_L g529 ( .A(n_508), .B(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g594 ( .A(n_508), .B(n_519), .Y(n_594) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g635 ( .A(n_509), .B(n_519), .Y(n_635) );
AND2x2_ASAP7_75t_L g679 ( .A(n_509), .B(n_518), .Y(n_679) );
AND2x2_ASAP7_75t_L g562 ( .A(n_518), .B(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g580 ( .A(n_518), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_518), .B(n_609), .Y(n_733) );
INVx3_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g528 ( .A(n_519), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_519), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g647 ( .A(n_519), .B(n_578), .Y(n_647) );
AND2x2_ASAP7_75t_L g674 ( .A(n_519), .B(n_609), .Y(n_674) );
OR2x2_ASAP7_75t_L g730 ( .A(n_519), .B(n_581), .Y(n_730) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_526), .Y(n_519) );
INVx1_ASAP7_75t_SL g616 ( .A(n_528), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_529), .B(n_647), .Y(n_648) );
AND2x2_ASAP7_75t_L g682 ( .A(n_529), .B(n_672), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_529), .B(n_605), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_529), .B(n_727), .Y(n_726) );
OAI31xp33_ASAP7_75t_L g700 ( .A1(n_531), .A2(n_562), .A3(n_701), .B(n_703), .Y(n_700) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_543), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_532), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g683 ( .A(n_532), .B(n_618), .Y(n_683) );
OR2x2_ASAP7_75t_L g690 ( .A(n_532), .B(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g702 ( .A(n_532), .B(n_591), .Y(n_702) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g636 ( .A(n_533), .B(n_637), .Y(n_636) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g564 ( .A(n_534), .B(n_565), .Y(n_564) );
INVx4_ASAP7_75t_L g585 ( .A(n_534), .Y(n_585) );
AND2x2_ASAP7_75t_L g622 ( .A(n_534), .B(n_566), .Y(n_622) );
AND2x2_ASAP7_75t_L g621 ( .A(n_543), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g691 ( .A(n_543), .Y(n_691) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_553), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_544), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g591 ( .A(n_544), .B(n_554), .Y(n_591) );
INVx2_ASAP7_75t_L g611 ( .A(n_544), .Y(n_611) );
AND2x2_ASAP7_75t_L g625 ( .A(n_544), .B(n_554), .Y(n_625) );
AND2x2_ASAP7_75t_L g632 ( .A(n_544), .B(n_588), .Y(n_632) );
BUFx3_ASAP7_75t_L g642 ( .A(n_544), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_544), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g587 ( .A(n_553), .Y(n_587) );
AND2x2_ASAP7_75t_L g595 ( .A(n_553), .B(n_585), .Y(n_595) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g565 ( .A(n_554), .B(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_554), .Y(n_619) );
INVx2_ASAP7_75t_SL g602 ( .A(n_563), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_563), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_563), .B(n_672), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_564), .B(n_642), .Y(n_695) );
INVx1_ASAP7_75t_SL g729 ( .A(n_564), .Y(n_729) );
INVx1_ASAP7_75t_SL g637 ( .A(n_565), .Y(n_637) );
INVx1_ASAP7_75t_SL g588 ( .A(n_566), .Y(n_588) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_566), .Y(n_599) );
OR2x2_ASAP7_75t_L g610 ( .A(n_566), .B(n_585), .Y(n_610) );
AND2x2_ASAP7_75t_L g624 ( .A(n_566), .B(n_585), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_566), .B(n_614), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_580), .B(n_582), .C(n_593), .Y(n_575) );
AOI31xp33_ASAP7_75t_L g692 ( .A1(n_576), .A2(n_693), .A3(n_694), .B(n_695), .Y(n_692) );
AND2x2_ASAP7_75t_L g665 ( .A(n_577), .B(n_594), .Y(n_665) );
BUFx3_ASAP7_75t_L g605 ( .A(n_578), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_578), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g641 ( .A(n_578), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_578), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g596 ( .A(n_581), .Y(n_596) );
OAI222xp33_ASAP7_75t_L g705 ( .A1(n_581), .A2(n_706), .B1(n_709), .B2(n_710), .C1(n_711), .C2(n_712), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_589), .Y(n_582) );
INVx1_ASAP7_75t_L g711 ( .A(n_583), .Y(n_711) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_585), .B(n_588), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_585), .B(n_611), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_585), .B(n_586), .Y(n_681) );
INVx1_ASAP7_75t_L g732 ( .A(n_585), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_586), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g734 ( .A(n_586), .Y(n_734) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx2_ASAP7_75t_L g614 ( .A(n_587), .Y(n_614) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_588), .Y(n_657) );
AOI32xp33_ASAP7_75t_L g593 ( .A1(n_589), .A2(n_594), .A3(n_595), .B1(n_596), .B2(n_597), .Y(n_593) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_591), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g668 ( .A(n_591), .Y(n_668) );
OR2x2_ASAP7_75t_L g709 ( .A(n_591), .B(n_610), .Y(n_709) );
INVx1_ASAP7_75t_L g645 ( .A(n_592), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_594), .B(n_605), .Y(n_630) );
INVx3_ASAP7_75t_L g639 ( .A(n_594), .Y(n_639) );
AOI322xp5_ASAP7_75t_L g655 ( .A1(n_594), .A2(n_639), .A3(n_656), .B1(n_658), .B2(n_661), .C1(n_665), .C2(n_666), .Y(n_655) );
AND2x2_ASAP7_75t_L g631 ( .A(n_595), .B(n_632), .Y(n_631) );
INVxp67_ASAP7_75t_L g708 ( .A(n_595), .Y(n_708) );
A2O1A1O1Ixp25_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_603), .C(n_611), .D(n_612), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_599), .B(n_642), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_601), .A2(n_613), .B1(n_616), .B2(n_617), .C(n_620), .Y(n_612) );
INVx1_ASAP7_75t_SL g727 ( .A(n_601), .Y(n_727) );
AOI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .B(n_610), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_605), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI221xp5_ASAP7_75t_SL g697 ( .A1(n_607), .A2(n_691), .B1(n_698), .B2(n_699), .C(n_700), .Y(n_697) );
OAI222xp33_ASAP7_75t_L g728 ( .A1(n_608), .A2(n_729), .B1(n_730), .B2(n_731), .C1(n_733), .C2(n_734), .Y(n_728) );
AND2x2_ASAP7_75t_L g686 ( .A(n_609), .B(n_672), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_609), .A2(n_624), .B(n_671), .Y(n_698) );
INVx1_ASAP7_75t_L g712 ( .A(n_609), .Y(n_712) );
INVx2_ASAP7_75t_SL g615 ( .A(n_610), .Y(n_615) );
AND2x2_ASAP7_75t_L g618 ( .A(n_611), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_SL g652 ( .A(n_614), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_614), .B(n_624), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_615), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_615), .B(n_625), .Y(n_654) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_623), .B(n_626), .Y(n_620) );
INVx1_ASAP7_75t_SL g638 ( .A(n_622), .Y(n_638) );
AND2x2_ASAP7_75t_L g685 ( .A(n_622), .B(n_668), .Y(n_685) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g724 ( .A(n_624), .B(n_642), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_625), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g710 ( .A(n_626), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B1(n_633), .B2(n_640), .C(n_643), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_637), .A2(n_644), .B1(n_646), .B2(n_648), .Y(n_643) );
OR2x2_ASAP7_75t_L g714 ( .A(n_638), .B(n_642), .Y(n_714) );
OR2x2_ASAP7_75t_L g717 ( .A(n_638), .B(n_652), .Y(n_717) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_659), .A2(n_714), .B1(n_715), .B2(n_717), .C(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND3xp33_ASAP7_75t_SL g669 ( .A(n_670), .B(n_684), .C(n_696), .Y(n_669) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B1(n_677), .B2(n_680), .C1(n_682), .C2(n_683), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_672), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g694 ( .A(n_674), .Y(n_694) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_687), .B2(n_689), .C(n_692), .Y(n_684) );
INVx1_ASAP7_75t_L g699 ( .A(n_685), .Y(n_699) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI21xp33_ASAP7_75t_L g718 ( .A1(n_689), .A2(n_719), .B(n_720), .Y(n_718) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
NOR5xp2_ASAP7_75t_L g696 ( .A(n_697), .B(n_705), .C(n_713), .D(n_722), .E(n_728), .Y(n_696) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
endmodule