module fake_jpeg_17084_n_166 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_6),
.Y(n_24)
);

AOI21xp33_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_26),
.B(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_6),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_20),
.Y(n_28)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_18),
.B1(n_13),
.B2(n_20),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_41),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_23),
.A2(n_17),
.B1(n_11),
.B2(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_14),
.B1(n_19),
.B2(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_14),
.B1(n_19),
.B2(n_13),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_22),
.B1(n_28),
.B2(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_30),
.B1(n_22),
.B2(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_9),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_53),
.Y(n_56)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_38),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_35),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_61),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_62),
.B(n_68),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_2),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_49),
.B(n_47),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_80),
.B(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_62),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_55),
.B1(n_50),
.B2(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_50),
.B1(n_68),
.B2(n_35),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_54),
.B(n_42),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_28),
.C(n_29),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_72),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_52),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_57),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_73),
.B(n_82),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_81),
.C(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_61),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_62),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_80),
.B1(n_79),
.B2(n_70),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_107),
.C(n_102),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_82),
.B(n_68),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_102),
.B(n_20),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_104),
.B1(n_38),
.B2(n_39),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_74),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_109),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_115),
.C(n_117),
.Y(n_126)
);

XOR2x2_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_94),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_28),
.B(n_34),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_85),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_114),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_79),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_91),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_88),
.B1(n_65),
.B2(n_35),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_119),
.B1(n_121),
.B2(n_106),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_96),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_35),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_106),
.C(n_105),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_64),
.B1(n_66),
.B2(n_39),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_111),
.C(n_20),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_124),
.B1(n_115),
.B2(n_128),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_29),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_113),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_136),
.B1(n_29),
.B2(n_27),
.Y(n_145)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_127),
.C(n_126),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_66),
.B1(n_34),
.B2(n_2),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_34),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_143),
.C(n_146),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_127),
.B1(n_4),
.B2(n_5),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_29),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_29),
.C(n_27),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_3),
.Y(n_154)
);

NAND4xp25_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_139),
.C(n_138),
.D(n_134),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_151),
.B(n_144),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_27),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_10),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_158),
.A3(n_3),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_150),
.B(n_5),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_146),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.C(n_8),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_9),
.C(n_10),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_10),
.Y(n_166)
);


endmodule