module fake_jpeg_968_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_SL g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_0),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_16),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_5),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_10),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_7),
.B(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_3),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_15),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_24),
.B1(n_16),
.B2(n_17),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_32),
.B(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_26),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_23),
.B1(n_15),
.B2(n_20),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_32),
.C(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_40),
.Y(n_43)
);

AOI321xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_39),
.A3(n_35),
.B1(n_36),
.B2(n_28),
.C(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_29),
.B(n_19),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_6),
.C(n_19),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_8),
.B1(n_45),
.B2(n_14),
.Y(n_47)
);


endmodule