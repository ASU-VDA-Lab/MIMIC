module fake_jpeg_5697_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_29),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

OR2x2_ASAP7_75t_SL g52 ( 
.A(n_28),
.B(n_24),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_30),
.B(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_38),
.Y(n_56)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_47),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_50),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_57),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_13),
.B1(n_25),
.B2(n_23),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_55),
.B1(n_28),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_25),
.B1(n_23),
.B2(n_18),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_53),
.B(n_55),
.C(n_52),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_18),
.B1(n_17),
.B2(n_5),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_17),
.B1(n_4),
.B2(n_2),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_2),
.B1(n_7),
.B2(n_9),
.Y(n_74)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_67),
.B1(n_73),
.B2(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_35),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_70),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_27),
.B1(n_28),
.B2(n_8),
.Y(n_67)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_72),
.Y(n_81)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_11),
.B(n_42),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_90),
.B(n_91),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_85),
.B1(n_79),
.B2(n_68),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_47),
.B1(n_49),
.B2(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_46),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_57),
.A3(n_42),
.B1(n_11),
.B2(n_10),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_57),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_71),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_70),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_70),
.B1(n_68),
.B2(n_79),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_98),
.B1(n_80),
.B2(n_82),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_75),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_102),
.C(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_93),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_77),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_108),
.C(n_110),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_85),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_107),
.B(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_102),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_96),
.B(n_97),
.C(n_100),
.D(n_90),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_81),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_101),
.C(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_105),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_118),
.Y(n_120)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_117),
.B(n_111),
.C(n_118),
.D(n_112),
.Y(n_121)
);

OAI21x1_ASAP7_75t_SL g123 ( 
.A1(n_121),
.A2(n_122),
.B(n_77),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_114),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_123),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_122),
.B(n_71),
.Y(n_125)
);


endmodule