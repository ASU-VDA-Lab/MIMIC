module fake_jpeg_27252_n_145 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.C(n_41),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_26),
.C(n_19),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_29),
.B1(n_25),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_56),
.B1(n_33),
.B2(n_16),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_40),
.B1(n_29),
.B2(n_25),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_55),
.B1(n_28),
.B2(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_31),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_40),
.B1(n_34),
.B2(n_38),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_33),
.B1(n_35),
.B2(n_38),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_31),
.B1(n_17),
.B2(n_15),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_70),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_69),
.B1(n_53),
.B2(n_45),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_27),
.B1(n_30),
.B2(n_21),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_23),
.B1(n_17),
.B2(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_68),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_35),
.B1(n_41),
.B2(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NAND2xp67_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_0),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_42),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_60),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_44),
.A3(n_42),
.B1(n_54),
.B2(n_45),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_65),
.B1(n_53),
.B2(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_71),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_69),
.B(n_61),
.C(n_63),
.Y(n_93)
);

OAI22x1_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_78),
.B1(n_80),
.B2(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_96),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_67),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_57),
.B(n_45),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_85),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_89),
.B1(n_53),
.B2(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_82),
.B1(n_75),
.B2(n_78),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_102),
.A2(n_103),
.B1(n_96),
.B2(n_90),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_106),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_85),
.C(n_89),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_84),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_1),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_113),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_118),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_107),
.C(n_114),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_3),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_125),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_111),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_126),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_103),
.B(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_108),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_93),
.B(n_117),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_4),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_122),
.B(n_124),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_133),
.A2(n_6),
.B(n_7),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_124),
.C(n_126),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_135),
.B(n_131),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_136),
.A2(n_128),
.B1(n_129),
.B2(n_4),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_139),
.B(n_140),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_134),
.C(n_5),
.Y(n_142)
);

AOI21x1_ASAP7_75t_L g140 ( 
.A1(n_136),
.A2(n_9),
.B(n_13),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_9),
.B(n_5),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_143),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_141),
.Y(n_145)
);


endmodule