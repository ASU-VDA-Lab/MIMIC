module fake_jpeg_20812_n_259 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_259);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_259;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_17),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_27),
.Y(n_60)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_42),
.Y(n_69)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_31),
.Y(n_74)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx12f_ASAP7_75t_SL g47 ( 
.A(n_22),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_22),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_25),
.B1(n_21),
.B2(n_44),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_56),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_18),
.B1(n_29),
.B2(n_26),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_63),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_25),
.B1(n_23),
.B2(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_60),
.B(n_73),
.Y(n_112)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_76),
.B1(n_86),
.B2(n_2),
.Y(n_110)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_66),
.Y(n_96)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_70),
.Y(n_100)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_24),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_85),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_20),
.B1(n_32),
.B2(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_24),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_30),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx6p67_ASAP7_75t_R g82 ( 
.A(n_36),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_16),
.Y(n_97)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_28),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_36),
.A2(n_20),
.B1(n_28),
.B2(n_16),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_41),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_44),
.B1(n_46),
.B2(n_33),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_16),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_22),
.B(n_33),
.C(n_16),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_113),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_52),
.B(n_46),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_84),
.C(n_66),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_104),
.B1(n_105),
.B2(n_117),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_75),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_46),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_33),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_115),
.B1(n_5),
.B2(n_6),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_56),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_54),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_48),
.B(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_92),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_49),
.B(n_4),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_113),
.A2(n_76),
.B1(n_64),
.B2(n_82),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_124),
.B1(n_125),
.B2(n_139),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_127),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_100),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_122),
.B(n_129),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_72),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_97),
.B(n_105),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_82),
.B1(n_72),
.B2(n_59),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_53),
.B1(n_71),
.B2(n_48),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_134),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_112),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_14),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_57),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_51),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_172)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_89),
.A2(n_53),
.B1(n_71),
.B2(n_51),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_102),
.Y(n_162)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_143),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_111),
.B1(n_106),
.B2(n_99),
.Y(n_160)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_107),
.B1(n_111),
.B2(n_98),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

NOR4xp25_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_98),
.C(n_107),
.D(n_105),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_142),
.A2(n_117),
.B(n_91),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_150),
.A2(n_152),
.B(n_162),
.Y(n_196)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_176),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_168),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_159),
.B1(n_160),
.B2(n_131),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_106),
.B1(n_99),
.B2(n_97),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_118),
.A2(n_147),
.B(n_131),
.C(n_139),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_136),
.B(n_134),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_7),
.C(n_9),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_171),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_102),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_132),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_7),
.B(n_9),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_128),
.Y(n_182)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_124),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_188),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_182),
.A2(n_186),
.B(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_189),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_119),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_190),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_140),
.C(n_125),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_161),
.B(n_130),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_193),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_10),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_12),
.B(n_13),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_11),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_172),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_163),
.B(n_183),
.Y(n_217)
);

OAI322xp33_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_162),
.A3(n_159),
.B1(n_163),
.B2(n_166),
.C1(n_172),
.C2(n_155),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_203),
.B(n_206),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_156),
.B1(n_157),
.B2(n_163),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_209),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_211),
.Y(n_218)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_153),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_SL g211 ( 
.A1(n_192),
.A2(n_195),
.A3(n_196),
.B1(n_179),
.B2(n_168),
.C1(n_185),
.C2(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_196),
.B(n_179),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_213),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_188),
.C(n_186),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_224),
.C(n_206),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_204),
.B(n_203),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_222),
.B(n_226),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_189),
.C(n_153),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_231),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_234),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_220),
.A2(n_209),
.B1(n_208),
.B2(n_197),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_219),
.Y(n_239)
);

NAND4xp25_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_168),
.C(n_202),
.D(n_208),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_216),
.B(n_226),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_207),
.B(n_213),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_214),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_238),
.A2(n_234),
.B(n_223),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_215),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_234),
.C(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_231),
.B1(n_233),
.B2(n_228),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_245),
.A2(n_247),
.B(n_249),
.Y(n_252)
);

OAI221xp5_ASAP7_75t_L g247 ( 
.A1(n_243),
.A2(n_197),
.B1(n_230),
.B2(n_235),
.C(n_227),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_248),
.A2(n_243),
.B(n_223),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_250),
.A2(n_253),
.B(n_252),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_149),
.B(n_151),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_254),
.A2(n_176),
.B(n_13),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_251),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_256),
.B(n_149),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_244),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_258),
.CI(n_232),
.CON(n_259),
.SN(n_259)
);


endmodule