module real_jpeg_30574_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_0),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g376 ( 
.A(n_0),
.Y(n_376)
);

NAND2x1p5_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_1),
.Y(n_166)
);

NAND2xp33_ASAP7_75t_R g284 ( 
.A(n_1),
.B(n_285),
.Y(n_284)
);

NAND2x1_ASAP7_75t_L g290 ( 
.A(n_1),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_1),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_1),
.B(n_385),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_1),
.B(n_154),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_1),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_1),
.B(n_282),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

AND2x4_ASAP7_75t_L g64 ( 
.A(n_2),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_2),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_2),
.B(n_123),
.Y(n_122)
);

NAND2x1p5_ASAP7_75t_L g187 ( 
.A(n_2),
.B(n_106),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_2),
.B(n_246),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_2),
.B(n_468),
.Y(n_467)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_3),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_3),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_3),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_3),
.B(n_325),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_3),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_3),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_3),
.B(n_418),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_5),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_5),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_5),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_5),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_5),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_5),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_5),
.B(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_6),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_8),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_8),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_9),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_9),
.B(n_45),
.Y(n_52)
);

NAND2x1_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_9),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_9),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_9),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_9),
.B(n_282),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_9),
.B(n_476),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_9),
.B(n_499),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_11),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_37),
.Y(n_36)
);

AND2x4_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_59),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_12),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_12),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_12),
.B(n_34),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_12),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_12),
.B(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_14),
.B(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_14),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_14),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_14),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_14),
.B(n_471),
.Y(n_470)
);

NAND2x1_ASAP7_75t_SL g480 ( 
.A(n_14),
.B(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_14),
.B(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_16),
.Y(n_259)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_16),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_75),
.Y(n_74)
);

NAND2x1_ASAP7_75t_L g105 ( 
.A(n_17),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_17),
.B(n_120),
.Y(n_119)
);

AND2x4_ASAP7_75t_SL g174 ( 
.A(n_17),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_17),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_17),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_17),
.B(n_359),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_17),
.Y(n_374)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_234),
.B(n_458),
.C(n_551),
.D(n_568),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_337),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_272),
.B(n_333),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g337 ( 
.A(n_26),
.B(n_338),
.C(n_340),
.Y(n_337)
);

AOI22x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_190),
.B1(n_226),
.B2(n_268),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_28),
.B(n_191),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_114),
.Y(n_28)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_29),
.B(n_270),
.C(n_271),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_77),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_54),
.Y(n_30)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_31),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_43),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_32),
.A2(n_49),
.B(n_261),
.C(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.C(n_39),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_33),
.A2(n_36),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_33),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_33),
.A2(n_110),
.B1(n_203),
.B2(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_36),
.A2(n_111),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_36),
.B(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_36),
.B(n_358),
.Y(n_382)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_38),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_39),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_39),
.Y(n_497)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_41),
.Y(n_209)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_41),
.Y(n_242)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_41),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_44),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_44),
.B(n_53),
.Y(n_262)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_48),
.Y(n_331)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_49),
.A2(n_53),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_49),
.A2(n_53),
.B1(n_80),
.B2(n_488),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_L g568 ( 
.A(n_49),
.B(n_80),
.C(n_466),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_51),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_51),
.Y(n_246)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_51),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_53),
.B(n_252),
.C(n_518),
.Y(n_517)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_54),
.B(n_77),
.C(n_267),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_67),
.C(n_72),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_56),
.B(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.C(n_64),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_58),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_61),
.B(n_64),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_62),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_64),
.B(n_183),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g362 ( 
.A1(n_64),
.A2(n_182),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_64),
.B(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_68),
.A2(n_74),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_70),
.Y(n_387)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_71),
.Y(n_186)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_76),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_93),
.C(n_108),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_78),
.A2(n_79),
.B1(n_93),
.B2(n_94),
.Y(n_222)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

OAI22x1_ASAP7_75t_L g178 ( 
.A1(n_80),
.A2(n_90),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_80),
.A2(n_196),
.B1(n_198),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_80),
.Y(n_488)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2x1_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_86),
.B(n_90),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_88),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.C(n_105),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2x2_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_97),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_163)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_98),
.Y(n_434)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_101),
.B(n_241),
.C(n_490),
.Y(n_527)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_102),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_102),
.Y(n_247)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_108),
.Y(n_221)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_110),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_111),
.B(n_173),
.C(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_112),
.A2(n_493),
.B1(n_494),
.B2(n_497),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_169),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_144),
.C(n_149),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_116),
.B(n_144),
.C(n_149),
.Y(n_270)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_117),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_131),
.C(n_141),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_118),
.B(n_141),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.C(n_126),
.Y(n_118)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_119),
.B(n_171),
.Y(n_279)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_122),
.Y(n_253)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_125),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_126),
.B(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_129),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_131),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_137),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_132),
.B(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_135),
.B(n_137),
.Y(n_201)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_137),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_137),
.A2(n_196),
.B1(n_198),
.B2(n_465),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_137),
.A2(n_465),
.B1(n_524),
.B2(n_525),
.Y(n_523)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_139),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_140),
.Y(n_326)
);

BUFx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_145),
.B(n_150),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.C(n_163),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_151),
.A2(n_152),
.B1(n_156),
.B2(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_155),
.Y(n_215)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_163),
.A2(n_281),
.B(n_284),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_167),
.Y(n_285)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_168),
.Y(n_473)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_169),
.Y(n_271)
);

XOR2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_170),
.B(n_178),
.C(n_181),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_175),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_176),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_182),
.A2(n_183),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_188),
.C(n_189),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_183),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_183),
.B(n_213),
.C(n_234),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_187),
.B(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_189),
.B(n_196),
.C(n_465),
.Y(n_483)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_219),
.C(n_223),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_192),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.C(n_216),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_193),
.B(n_217),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g561 ( 
.A(n_196),
.B(n_488),
.C(n_489),
.Y(n_561)
);

XOR2x2_ASAP7_75t_SL g275 ( 
.A(n_199),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.C(n_205),
.Y(n_199)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_200),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_202),
.B(n_206),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_203),
.Y(n_318)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.C(n_213),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_207),
.A2(n_213),
.B1(n_214),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_207),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_210),
.B(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_214),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_213),
.A2(n_214),
.B1(n_466),
.B2(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_214),
.B(n_465),
.C(n_466),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_215),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_220),
.B(n_224),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_227),
.B(n_269),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_227),
.B(n_269),
.Y(n_336)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_266),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_249),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_229),
.Y(n_548)
);

XOR2x2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_230),
.B(n_238),
.C(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_248),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g512 ( 
.A(n_240),
.Y(n_512)
);

XNOR2x1_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_245),
.Y(n_490)
);

INVxp33_ASAP7_75t_SL g549 ( 
.A(n_249),
.Y(n_549)
);

OAI22x1_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_249)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_260),
.Y(n_250)
);

INVxp33_ASAP7_75t_SL g538 ( 
.A(n_251),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_256),
.Y(n_518)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g539 ( 
.A(n_260),
.Y(n_539)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_264),
.B(n_538),
.C(n_539),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_266),
.A2(n_547),
.B(n_550),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_300),
.B(n_332),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_339),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_298),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_298),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.C(n_295),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_295),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.C(n_286),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_286),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.C(n_290),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_288),
.B(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_289),
.B(n_290),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

XNOR2x2_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_303),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.C(n_311),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_312),
.Y(n_343)
);

XNOR2x1_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.C(n_319),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_313),
.B(n_347),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_316),
.A2(n_317),
.B1(n_319),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_324),
.C(n_327),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_320),
.A2(n_321),
.B1(n_327),
.B2(n_328),
.Y(n_448)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_323),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_324),
.B(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B(n_336),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_365),
.B(n_456),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_342),
.Y(n_457)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_345),
.B(n_457),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.C(n_352),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_346),
.B(n_452),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_349),
.A2(n_350),
.B1(n_352),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_352),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_356),
.C(n_362),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_353),
.A2(n_354),
.B1(n_362),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_356),
.B(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_362),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_450),
.B(n_455),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_439),
.B(n_449),
.Y(n_366)
);

AOI21x1_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_409),
.B(n_438),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_401),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_383),
.B1(n_399),
.B2(n_400),
.Y(n_369)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

AOI221xp5_ASAP7_75t_L g438 ( 
.A1(n_370),
.A2(n_383),
.B1(n_399),
.B2(n_400),
.C(n_401),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_381),
.B2(n_382),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_371),
.B(n_382),
.C(n_400),
.Y(n_440)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_377),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_377),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx6_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_383),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_388),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_384),
.B(n_389),
.C(n_393),
.Y(n_446)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_393),
.B1(n_397),
.B2(n_398),
.Y(n_388)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_389),
.Y(n_397)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_393),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.C(n_405),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_402),
.A2(n_403),
.B1(n_421),
.B2(n_422),
.Y(n_420)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_404),
.A2(n_405),
.B1(n_406),
.B2(n_423),
.Y(n_422)
);

CKINVDCx12_ASAP7_75t_R g423 ( 
.A(n_404),
.Y(n_423)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_424),
.B(n_437),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_420),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_420),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_417),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_417),
.Y(n_426)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx5_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_430),
.B(n_436),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_426),
.B(n_427),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_435),
.Y(n_430)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_441),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_445),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_446),
.C(n_447),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_SL g455 ( 
.A(n_451),
.B(n_454),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_529),
.Y(n_458)
);

OAI211xp5_ASAP7_75t_L g551 ( 
.A1(n_459),
.A2(n_552),
.B(n_555),
.C(n_556),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_509),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_460),
.B(n_509),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_491),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_478),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_462),
.B(n_478),
.C(n_491),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_469),
.C(n_474),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_464),
.B(n_507),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_466),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_466),
.A2(n_526),
.B1(n_563),
.B2(n_564),
.Y(n_562)
);

BUFx4f_ASAP7_75t_SL g466 ( 
.A(n_467),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_470),
.A2(n_474),
.B1(n_475),
.B2(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_470),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_486),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_480),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_480),
.Y(n_484)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_483),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_483),
.B(n_484),
.C(n_486),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_R g491 ( 
.A(n_492),
.B(n_503),
.C(n_506),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_504),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_497),
.C(n_498),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_498),
.Y(n_514)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_521),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_519),
.C(n_522),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_510),
.B(n_541),
.Y(n_540)
);

MAJx2_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_513),
.C(n_516),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_511),
.B(n_534),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_513),
.B(n_517),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_520),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_522),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_527),
.C(n_528),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_528),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_543),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_530),
.A2(n_553),
.B(n_554),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_540),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_531),
.B(n_540),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_535),
.C(n_537),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_533),
.B(n_545),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_535),
.B(n_537),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_544),
.B(n_546),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_544),
.B(n_546),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_549),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_548),
.B(n_549),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_557),
.B(n_560),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_567),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_566),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_560),
.A2(n_561),
.B1(n_562),
.B2(n_565),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_562),
.Y(n_565)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);


endmodule