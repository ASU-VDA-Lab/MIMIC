module fake_jpeg_19789_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_0),
.B(n_5),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_77),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_85),
.Y(n_98)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_49),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_66),
.B1(n_50),
.B2(n_59),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_55),
.B1(n_51),
.B2(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_45),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_67),
.B1(n_64),
.B2(n_61),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_86),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_93),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_99),
.B1(n_3),
.B2(n_6),
.Y(n_110)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_63),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_62),
.CI(n_48),
.CON(n_101),
.SN(n_101)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_24),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_57),
.A3(n_84),
.B1(n_60),
.B2(n_56),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_8),
.B(n_9),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_53),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_27),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_7),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_11),
.B1(n_15),
.B2(n_17),
.Y(n_117)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_10),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_18),
.B1(n_22),
.B2(n_23),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_120),
.C(n_121),
.Y(n_123)
);

OAI321xp33_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_112),
.A3(n_108),
.B1(n_100),
.B2(n_107),
.C(n_101),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_111),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_102),
.B(n_118),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_122),
.C(n_29),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_28),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_36),
.C(n_39),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_40),
.B(n_41),
.Y(n_136)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_136),
.Y(n_137)
);


endmodule