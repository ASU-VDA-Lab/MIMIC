module fake_jpeg_5195_n_337 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_44),
.Y(n_67)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_53),
.B1(n_17),
.B2(n_33),
.Y(n_72)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_0),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_62),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_49),
.B1(n_17),
.B2(n_47),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_61),
.A2(n_100),
.B1(n_104),
.B2(n_12),
.Y(n_128)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_78),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_29),
.B1(n_24),
.B2(n_19),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_73),
.A2(n_76),
.B1(n_88),
.B2(n_98),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_24),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_80),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_29),
.B1(n_33),
.B2(n_23),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_79),
.B1(n_86),
.B2(n_91),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_38),
.B1(n_42),
.B2(n_51),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_44),
.A2(n_36),
.B1(n_32),
.B2(n_31),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_89),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_25),
.B1(n_32),
.B2(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_36),
.B1(n_32),
.B2(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_95),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_25),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_13),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_97),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_36),
.B1(n_30),
.B2(n_28),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_101),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_30),
.B1(n_28),
.B2(n_22),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_43),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_43),
.A2(n_30),
.B1(n_28),
.B2(n_22),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_37),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_37),
.A3(n_22),
.B1(n_12),
.B2(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_117),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_0),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_88),
.B1(n_76),
.B2(n_100),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_131),
.B1(n_96),
.B2(n_95),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_71),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_72),
.B1(n_81),
.B2(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_129),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_57),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_94),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_165)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_61),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_4),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_84),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_68),
.B(n_80),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_6),
.Y(n_160)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_142),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_141),
.A2(n_165),
.B1(n_158),
.B2(n_140),
.Y(n_200)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_143),
.A2(n_154),
.B1(n_170),
.B2(n_171),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_66),
.C(n_93),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_145),
.C(n_161),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_103),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_104),
.B1(n_78),
.B2(n_89),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_146),
.A2(n_174),
.B1(n_169),
.B2(n_173),
.Y(n_214)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_151),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_102),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g207 ( 
.A1(n_150),
.A2(n_176),
.A3(n_126),
.B1(n_130),
.B2(n_137),
.Y(n_207)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_131),
.B(n_134),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_105),
.B(n_101),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_168),
.B(n_175),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_69),
.B1(n_87),
.B2(n_59),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_97),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_158),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_108),
.B(n_5),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_160),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_70),
.C(n_8),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_6),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_166),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_110),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_167),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_6),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_113),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_124),
.A2(n_10),
.B1(n_11),
.B2(n_125),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_106),
.A2(n_10),
.B1(n_11),
.B2(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_10),
.Y(n_172)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_173),
.A2(n_134),
.B1(n_137),
.B2(n_114),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_118),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_121),
.A2(n_111),
.B(n_122),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_108),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_121),
.B1(n_128),
.B2(n_138),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_179),
.A2(n_200),
.B1(n_212),
.B2(n_214),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_180),
.B(n_187),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_184),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_108),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_186),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_131),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_115),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_199),
.Y(n_225)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_196),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_115),
.C(n_114),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_210),
.C(n_168),
.Y(n_234)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_126),
.C(n_130),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_204),
.B(n_168),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_159),
.A2(n_162),
.B1(n_134),
.B2(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_160),
.Y(n_222)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_126),
.C(n_130),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_141),
.A2(n_155),
.B1(n_170),
.B2(n_175),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_230),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_229),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_152),
.B(n_155),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_235),
.B(n_189),
.Y(n_250)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_226),
.B(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_147),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_231),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_186),
.A2(n_154),
.B1(n_143),
.B2(n_163),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_195),
.B1(n_194),
.B2(n_191),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_172),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_234),
.C(n_197),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_198),
.A2(n_196),
.B(n_188),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_190),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_203),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_198),
.B(n_192),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_250),
.Y(n_282)
);

NOR4xp25_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_207),
.C(n_182),
.D(n_189),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_246),
.B(n_215),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_212),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_248),
.C(n_254),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_185),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_236),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_210),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_185),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_262),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_179),
.C(n_201),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_261),
.C(n_224),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_205),
.C(n_195),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_227),
.A2(n_194),
.B(n_209),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_217),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_191),
.B1(n_217),
.B2(n_213),
.Y(n_281)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_237),
.C(n_223),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_216),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_240),
.A2(n_221),
.B1(n_238),
.B2(n_224),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_232),
.B1(n_215),
.B2(n_220),
.Y(n_275)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_270),
.B(n_278),
.Y(n_295)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_252),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_216),
.Y(n_274)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_280),
.B1(n_250),
.B2(n_258),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_251),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_246),
.Y(n_293)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_244),
.B(n_230),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_281),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_228),
.B1(n_226),
.B2(n_218),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_262),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_218),
.B1(n_239),
.B2(n_208),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_284),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_239),
.C(n_254),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_252),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_291),
.B1(n_297),
.B2(n_258),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_275),
.A2(n_249),
.B1(n_271),
.B2(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_282),
.Y(n_302)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_299),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_268),
.A2(n_267),
.B1(n_257),
.B2(n_251),
.Y(n_297)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_256),
.B(n_277),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_300),
.A2(n_307),
.B(n_287),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_287),
.B1(n_296),
.B2(n_294),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_302),
.B(n_297),
.Y(n_317)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_247),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_310),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_269),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_269),
.C(n_288),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_256),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_282),
.B1(n_280),
.B2(n_276),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_294),
.B1(n_295),
.B2(n_298),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_291),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_255),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_263),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_316),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_320),
.B(n_308),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_318),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_272),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_305),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_313),
.A2(n_301),
.B1(n_319),
.B2(n_305),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_327),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_314),
.A2(n_245),
.B1(n_300),
.B2(n_307),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_317),
.C(n_261),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_326),
.B(n_315),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_312),
.A2(n_285),
.B(n_259),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_326),
.B1(n_324),
.B2(n_316),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_323),
.B(n_321),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_333),
.B(n_328),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_323),
.C(n_330),
.Y(n_335)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_325),
.B(n_306),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_300),
.Y(n_337)
);


endmodule