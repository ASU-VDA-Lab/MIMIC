module real_jpeg_23465_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_349, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_349;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_69),
.B1(n_70),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_1),
.A2(n_74),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_74),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_74),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_4),
.A2(n_12),
.B1(n_89),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_4),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_4),
.A2(n_69),
.B1(n_70),
.B2(n_99),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_99),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_99),
.Y(n_198)
);

INVx8_ASAP7_75t_SL g85 ( 
.A(n_5),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_6),
.A2(n_91),
.B(n_93),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_6),
.B(n_82),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_95),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_6),
.B(n_30),
.C(n_31),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_6),
.B(n_72),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_6),
.A2(n_46),
.B1(n_192),
.B2(n_198),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_7),
.A2(n_44),
.B1(n_69),
.B2(n_70),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_7),
.A2(n_44),
.B1(n_89),
.B2(n_107),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_52),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_8),
.A2(n_52),
.B1(n_69),
.B2(n_70),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_8),
.A2(n_52),
.B1(n_91),
.B2(n_235),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_9),
.A2(n_61),
.B1(n_69),
.B2(n_70),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_61),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_9),
.A2(n_61),
.B1(n_89),
.B2(n_96),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_11),
.A2(n_69),
.B1(n_70),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_11),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_76),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_76),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_11),
.A2(n_76),
.B1(n_91),
.B2(n_235),
.Y(n_234)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_14),
.A2(n_38),
.B1(n_69),
.B2(n_70),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_14),
.A2(n_38),
.B1(n_88),
.B2(n_301),
.Y(n_300)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_15),
.Y(n_128)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_15),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_342),
.C(n_346),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_340),
.B(n_345),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_330),
.B(n_339),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_295),
.A3(n_325),
.B1(n_328),
.B2(n_329),
.C(n_349),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_271),
.B(n_294),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_245),
.B(n_270),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_135),
.B(n_218),
.C(n_244),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_120),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_24),
.B(n_120),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_102),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_57),
.B1(n_100),
.B2(n_101),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_26),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_26),
.B(n_101),
.C(n_102),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_45),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_27),
.B(n_45),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_34),
.B(n_39),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_28),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_28),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_28),
.B(n_95),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_28),
.A2(n_164),
.B(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_29),
.B(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_34),
.Y(n_227)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_35),
.A2(n_36),
.B1(n_67),
.B2(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_35),
.B(n_67),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_36),
.A2(n_68),
.A3(n_70),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_36),
.B(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_39),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_60),
.B(n_62),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_40),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_40),
.A2(n_152),
.B(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_40),
.A2(n_151),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_40),
.A2(n_150),
.B1(n_151),
.B2(n_172),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_40),
.A2(n_151),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_40),
.A2(n_62),
.B(n_228),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_40),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_50),
.B(n_53),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_46),
.A2(n_53),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_46),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_46),
.A2(n_189),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_46),
.A2(n_146),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_47),
.B(n_54),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_47),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_49),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.C(n_78),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_58),
.A2(n_59),
.B1(n_63),
.B2(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_73),
.B1(n_75),
.B2(n_77),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_75),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_64),
.A2(n_73),
.B1(n_77),
.B2(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_64),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_64),
.A2(n_77),
.B1(n_265),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_65),
.A2(n_72),
.B1(n_134),
.B2(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_65),
.B(n_240),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_65),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_65),
.A2(n_72),
.B(n_112),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_70),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_84),
.B(n_94),
.C(n_115),
.Y(n_114)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_69),
.B(n_95),
.CON(n_143),
.SN(n_143)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_83),
.C(n_96),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_72),
.B(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_77),
.A2(n_265),
.B(n_266),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_78),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_90),
.B2(n_97),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_82),
.B1(n_98),
.B2(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_80),
.A2(n_82),
.B1(n_106),
.B2(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_80),
.A2(n_234),
.B(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_80),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_80),
.B(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_80),
.A2(n_82),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_80),
.A2(n_286),
.B(n_319),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_80),
.A2(n_82),
.B(n_285),
.Y(n_346)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_81),
.B(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_81),
.B(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_81),
.A2(n_300),
.B(n_302),
.Y(n_299)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_91),
.Y(n_235)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_95),
.B(n_128),
.Y(n_203)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_105),
.B(n_109),
.C(n_113),
.Y(n_242)
);

INVx8_ASAP7_75t_L g301 ( 
.A(n_107),
.Y(n_301)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_111),
.B(n_266),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_112),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_116),
.B1(n_117),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_128),
.B(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_126),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_121),
.B(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_124),
.B(n_126),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_132),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_128),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_129),
.B(n_183),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_213),
.B(n_217),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_166),
.B(n_212),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_153),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_140),
.B(n_153),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_148),
.C(n_149),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_141),
.B(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_148),
.B(n_149),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_161),
.C(n_165),
.Y(n_214)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_165),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_160),
.Y(n_165)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_163),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_207),
.B(n_211),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_185),
.B(n_206),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_169),
.B(n_175),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_173),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_180),
.C(n_181),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_194),
.B(n_205),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_193),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_200),
.B(n_204),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_196),
.B(n_197),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_208),
.B(n_209),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_220),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_242),
.B2(n_243),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_230),
.C(n_243),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_229),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_229),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_226),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_241),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_236),
.C(n_241),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_246),
.B(n_247),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_269),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_256),
.B1(n_267),
.B2(n_268),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_268),
.C(n_269),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_252),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_253),
.B1(n_284),
.B2(n_288),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_252),
.A2(n_288),
.B(n_289),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_260),
.C(n_263),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_261),
.Y(n_343)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_273),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_292),
.B2(n_293),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_282),
.B1(n_290),
.B2(n_291),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_276),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_291),
.C(n_293),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_279),
.B(n_281),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_279),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_280),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_297),
.C(n_313),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_281),
.B(n_297),
.CI(n_313),
.CON(n_327),
.SN(n_327)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_289),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_284),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_314),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_314),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_304),
.B2(n_305),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_299),
.B1(n_316),
.B2(n_323),
.Y(n_315)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_307),
.C(n_310),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_323),
.C(n_324),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_300),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_302),
.B(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_310),
.B2(n_311),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_311),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_317),
.C(n_321),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_324),
.Y(n_314)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_327),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_332),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_338),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_337),
.C(n_338),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_344),
.Y(n_345)
);


endmodule