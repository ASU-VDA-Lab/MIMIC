module fake_jpeg_13509_n_184 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_23),
.B(n_12),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

INVx11_ASAP7_75t_SL g77 ( 
.A(n_38),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_27),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_10),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_87),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_91),
.Y(n_97)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_81),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_20),
.B(n_48),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_72),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_62),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_71),
.Y(n_113)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_76),
.B1(n_78),
.B2(n_70),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_78),
.B1(n_63),
.B2(n_70),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_128),
.B1(n_58),
.B2(n_73),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_114),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_57),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_60),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_121),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_64),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_77),
.B(n_54),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_125),
.Y(n_143)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_69),
.Y(n_121)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_71),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_58),
.B1(n_76),
.B2(n_77),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_67),
.C(n_54),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_120),
.C(n_9),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_133),
.B(n_142),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_138),
.B(n_122),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_124),
.A2(n_55),
.B1(n_67),
.B2(n_6),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_4),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_4),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_147),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_5),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_5),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_149),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_6),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_67),
.B1(n_24),
.B2(n_29),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_119),
.B1(n_31),
.B2(n_50),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_152),
.B(n_155),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_163),
.B(n_165),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_7),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_159),
.C(n_160),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_21),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_22),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_162),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_34),
.C(n_46),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_32),
.C(n_44),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_166),
.A2(n_129),
.B(n_138),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_131),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_145),
.C(n_143),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_176),
.C(n_158),
.Y(n_177)
);

INVxp33_ASAP7_75t_SL g178 ( 
.A(n_175),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_151),
.A3(n_156),
.B1(n_141),
.B2(n_164),
.C1(n_157),
.C2(n_150),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_168),
.C(n_167),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_173),
.B1(n_178),
.B2(n_169),
.Y(n_180)
);

OAI222xp33_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_170),
.B1(n_129),
.B2(n_143),
.C1(n_151),
.C2(n_165),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_166),
.B(n_136),
.Y(n_182)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_19),
.B1(n_43),
.B2(n_42),
.C(n_41),
.Y(n_183)
);

AOI321xp33_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_17),
.A3(n_37),
.B1(n_18),
.B2(n_47),
.C(n_16),
.Y(n_184)
);


endmodule