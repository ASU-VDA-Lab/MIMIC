module fake_jpeg_15847_n_157 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_157);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx11_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_48),
.B1(n_23),
.B2(n_14),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_26),
.B1(n_16),
.B2(n_25),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_14),
.B1(n_19),
.B2(n_23),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_36),
.B(n_22),
.C(n_21),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_27),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_36),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_60),
.B(n_66),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_17),
.B(n_28),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_33),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_65),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_37),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_28),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_68),
.B1(n_45),
.B2(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_19),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_45),
.B1(n_42),
.B2(n_50),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_76),
.Y(n_92)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

BUFx2_ASAP7_75t_SL g75 ( 
.A(n_58),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_89),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVxp33_ASAP7_75t_SL g85 ( 
.A(n_62),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_70),
.B(n_31),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_59),
.C(n_60),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_100),
.C(n_105),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_96),
.B1(n_97),
.B2(n_103),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_67),
.B1(n_70),
.B2(n_65),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_70),
.B1(n_33),
.B2(n_0),
.Y(n_97)
);

CKINVDCx6p67_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_35),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_101),
.B(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_31),
.B1(n_35),
.B2(n_22),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_21),
.C(n_18),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_81),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_118),
.C(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_74),
.CI(n_73),
.CON(n_113),
.SN(n_113)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_76),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_114),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_121),
.C(n_126),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_93),
.C(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_113),
.B1(n_118),
.B2(n_97),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_71),
.B1(n_18),
.B2(n_6),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_113),
.B1(n_106),
.B2(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_99),
.C(n_5),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_133),
.B(n_2),
.C(n_5),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_134),
.B(n_126),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVxp33_ASAP7_75t_SL g140 ( 
.A(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_138),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_128),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_125),
.B(n_124),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_7),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_145),
.B(n_146),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_144),
.B(n_131),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_135),
.C(n_120),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_147),
.A2(n_149),
.B1(n_9),
.B2(n_12),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_135),
.B1(n_10),
.B2(n_12),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_148),
.A2(n_9),
.B(n_10),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_152),
.C(n_147),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_38),
.C(n_154),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_38),
.Y(n_157)
);


endmodule