module real_jpeg_8220_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_43;
wire n_8;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_50;
wire n_33;
wire n_29;
wire n_49;
wire n_52;
wire n_10;
wire n_9;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_48;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

OR2x2_ASAP7_75t_SL g21 ( 
.A(n_1),
.B(n_3),
.Y(n_21)
);

OR2x2_ASAP7_75t_SL g37 ( 
.A(n_1),
.B(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_2),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_2),
.B(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_2),
.A2(n_22),
.B1(n_50),
.B2(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_4),
.A2(n_5),
.B1(n_14),
.B2(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g12 ( 
.A1(n_5),
.A2(n_13),
.B(n_15),
.Y(n_12)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

OA21x2_ASAP7_75t_L g42 ( 
.A1(n_5),
.A2(n_43),
.B(n_45),
.Y(n_42)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_11),
.B(n_17),
.C(n_48),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_8),
.B(n_32),
.Y(n_52)
);

OR2x2_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_16),
.Y(n_11)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

OAI211xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B(n_25),
.C(n_38),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_22),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_32),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_34),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);


endmodule