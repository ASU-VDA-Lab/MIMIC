module fake_jpeg_15520_n_67 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_2),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_10),
.A2(n_0),
.B(n_3),
.C(n_4),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_20),
.B(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_34),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_5),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_36),
.C(n_41),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_44),
.C(n_34),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_38),
.B1(n_23),
.B2(n_27),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_32),
.B1(n_39),
.B2(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_56),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_47),
.B1(n_49),
.B2(n_39),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_59),
.C(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_21),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_32),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_63),
.B(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_11),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_65),
.B1(n_16),
.B2(n_12),
.Y(n_67)
);


endmodule