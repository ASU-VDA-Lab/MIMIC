module fake_jpeg_8209_n_335 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_57),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_33),
.B1(n_21),
.B2(n_32),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_28),
.B1(n_18),
.B2(n_45),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_21),
.B1(n_19),
.B2(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_45),
.B1(n_38),
.B2(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_33),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_32),
.B1(n_19),
.B2(n_43),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_43),
.B1(n_38),
.B2(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_31),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_19),
.B1(n_24),
.B2(n_34),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_34),
.B1(n_18),
.B2(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_17),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_61),
.B(n_52),
.C(n_69),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_65),
.B1(n_54),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_65),
.B1(n_60),
.B2(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_17),
.Y(n_106)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_60),
.B1(n_48),
.B2(n_20),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_83),
.B1(n_35),
.B2(n_27),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_40),
.B1(n_26),
.B2(n_22),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_94),
.B1(n_65),
.B2(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_88),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_26),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_93),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_16),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_0),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_40),
.B1(n_13),
.B2(n_14),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_46),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_36),
.C(n_41),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_123),
.Y(n_134)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_111),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_108),
.B1(n_89),
.B2(n_74),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_126),
.B1(n_93),
.B2(n_77),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_117),
.B1(n_73),
.B2(n_93),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_115),
.Y(n_150)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_48),
.B1(n_20),
.B2(n_27),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_81),
.B1(n_94),
.B2(n_85),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_48),
.B1(n_20),
.B2(n_36),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_122),
.B(n_72),
.Y(n_136)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_63),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_35),
.B(n_17),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_96),
.C(n_79),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_88),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_51),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_131),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_145),
.B1(n_147),
.B2(n_104),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_72),
.B1(n_86),
.B2(n_91),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_151),
.B1(n_105),
.B2(n_116),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_142),
.B1(n_103),
.B2(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_137),
.B(n_140),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_98),
.C(n_72),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_98),
.C(n_87),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_93),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_154),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_73),
.B1(n_20),
.B2(n_41),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_160),
.Y(n_195)
);

AOI32xp33_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_118),
.A3(n_128),
.B1(n_106),
.B2(n_123),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_163),
.B(n_46),
.Y(n_211)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_162),
.B1(n_168),
.B2(n_170),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_99),
.B(n_111),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_173),
.B1(n_153),
.B2(n_148),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_108),
.B1(n_99),
.B2(n_126),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_163),
.B1(n_166),
.B2(n_170),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_99),
.B1(n_127),
.B2(n_109),
.Y(n_168)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_99),
.B1(n_107),
.B2(n_124),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_153),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_114),
.B1(n_109),
.B2(n_107),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_100),
.B1(n_107),
.B2(n_121),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_182),
.B1(n_135),
.B2(n_129),
.Y(n_203)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_136),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_107),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_180),
.C(n_132),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_179),
.B(n_147),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_100),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_136),
.A2(n_131),
.B1(n_141),
.B2(n_144),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_197),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_133),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_186),
.A2(n_190),
.B(n_84),
.Y(n_237)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_192),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_133),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_204),
.B1(n_174),
.B2(n_162),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_146),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_199),
.C(n_206),
.Y(n_215)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_156),
.B1(n_175),
.B2(n_51),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_155),
.C(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_41),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_1),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_209),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_46),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_212),
.C(n_180),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_16),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_46),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_216),
.A2(n_221),
.B1(n_230),
.B2(n_233),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_171),
.Y(n_217)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_178),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_219),
.C(n_238),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_170),
.B(n_173),
.C(n_156),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_190),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_201),
.B1(n_188),
.B2(n_186),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_175),
.B1(n_155),
.B2(n_84),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_229),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_84),
.B1(n_78),
.B2(n_3),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_210),
.Y(n_243)
);

OAI22x1_ASAP7_75t_L g233 ( 
.A1(n_186),
.A2(n_190),
.B1(n_191),
.B2(n_211),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_234),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_191),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_236),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_78),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_203),
.C(n_212),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_240),
.B(n_221),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_187),
.B(n_200),
.C(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_198),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_224),
.B(n_223),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_188),
.B1(n_206),
.B2(n_205),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_248),
.A2(n_255),
.B1(n_236),
.B2(n_228),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_237),
.B(n_230),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_1),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_238),
.C(n_219),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_256),
.C(n_257),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_78),
.B1(n_5),
.B2(n_6),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_4),
.C(n_5),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_4),
.C(n_5),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_213),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_260),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_4),
.Y(n_260)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_242),
.B(n_239),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_272),
.B(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_268),
.B(n_251),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_270),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_274),
.B1(n_278),
.B2(n_249),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_242),
.A2(n_221),
.B(n_235),
.Y(n_272)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_231),
.B1(n_214),
.B2(n_7),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_247),
.B(n_239),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_214),
.C(n_6),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_260),
.C(n_257),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_241),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_256),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_291),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_SL g286 ( 
.A(n_265),
.B(n_240),
.C(n_243),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_272),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_246),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_270),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_246),
.C(n_258),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_293),
.C(n_263),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_255),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_261),
.B1(n_264),
.B2(n_273),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_253),
.C(n_8),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_296),
.A2(n_7),
.B(n_8),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_283),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_276),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_303),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_302),
.B(n_274),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_282),
.B(n_274),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_SL g305 ( 
.A1(n_285),
.A2(n_268),
.B(n_263),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_7),
.Y(n_315)
);

OAI321xp33_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_274),
.A3(n_271),
.B1(n_266),
.B2(n_253),
.C(n_11),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_306),
.A2(n_279),
.B(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_311),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_300),
.A2(n_286),
.B1(n_283),
.B2(n_287),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_297),
.C(n_301),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_302),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_8),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_319),
.A2(n_321),
.B(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_295),
.C(n_303),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_310),
.Y(n_323)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_323),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_315),
.B(n_9),
.C(n_10),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_SL g331 ( 
.A1(n_325),
.A2(n_326),
.B(n_328),
.C(n_329),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_8),
.C(n_9),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_9),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_317),
.B(n_320),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_331),
.Y(n_333)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_320),
.B(n_11),
.Y(n_334)
);

OAI321xp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_11),
.A3(n_12),
.B1(n_324),
.B2(n_309),
.C(n_328),
.Y(n_335)
);


endmodule