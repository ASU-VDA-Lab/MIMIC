module fake_jpeg_15359_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_8),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_30),
.B1(n_35),
.B2(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_54),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_47),
.A2(n_41),
.B1(n_45),
.B2(n_17),
.Y(n_88)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_34),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_18),
.B1(n_34),
.B2(n_21),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_44),
.B1(n_18),
.B2(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp67_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_17),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_62),
.A2(n_55),
.B1(n_46),
.B2(n_67),
.Y(n_103)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_21),
.B1(n_18),
.B2(n_30),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_92)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_37),
.Y(n_73)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_90),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_44),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_0),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_41),
.B1(n_38),
.B2(n_19),
.Y(n_82)
);

OAI22x1_ASAP7_75t_L g130 ( 
.A1(n_82),
.A2(n_106),
.B1(n_92),
.B2(n_81),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_39),
.B(n_23),
.C(n_24),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_49),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_102),
.C(n_103),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_107),
.B1(n_0),
.B2(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_31),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_28),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_16),
.B(n_31),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_29),
.C(n_28),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_105),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_33),
.B1(n_48),
.B2(n_47),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_64),
.A2(n_29),
.B1(n_28),
.B2(n_16),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_109),
.A2(n_122),
.B(n_27),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_79),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_83),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_10),
.B1(n_11),
.B2(n_9),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_80),
.C(n_81),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_121),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_27),
.C(n_26),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_99),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_80),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_146),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_140),
.B(n_143),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_107),
.B1(n_96),
.B2(n_97),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_151),
.B1(n_154),
.B2(n_141),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_72),
.B(n_90),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_144),
.A2(n_13),
.B(n_4),
.Y(n_203)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_68),
.B1(n_101),
.B2(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_69),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_74),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_87),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_104),
.B1(n_98),
.B2(n_86),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_75),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_112),
.B(n_85),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_124),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_160),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_159),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_133),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_22),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_78),
.C(n_7),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_26),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_117),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_126),
.B1(n_136),
.B2(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_71),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_166),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_120),
.B(n_129),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_71),
.Y(n_168)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_170),
.A2(n_189),
.B1(n_145),
.B2(n_157),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_178),
.B(n_186),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_131),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_143),
.B(n_125),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_188),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_120),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_198),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_142),
.B(n_155),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_113),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_126),
.B1(n_136),
.B2(n_137),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_78),
.B1(n_10),
.B2(n_12),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_153),
.B1(n_152),
.B2(n_163),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_22),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_203),
.Y(n_221)
);

AOI22x1_ASAP7_75t_R g194 ( 
.A1(n_161),
.A2(n_22),
.B1(n_12),
.B2(n_15),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_196),
.Y(n_209)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_14),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_15),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_140),
.B(n_7),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_139),
.A2(n_2),
.B(n_3),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_2),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_167),
.C(n_151),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_204),
.B(n_205),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_166),
.C(n_160),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_154),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_211),
.A2(n_193),
.B(n_221),
.C(n_203),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_212),
.A2(n_216),
.B1(n_217),
.B2(n_220),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_170),
.A2(n_145),
.B1(n_164),
.B2(n_169),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_190),
.A2(n_169),
.B1(n_5),
.B2(n_6),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_223),
.B1(n_202),
.B2(n_191),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_195),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_232),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_178),
.A2(n_174),
.B1(n_190),
.B2(n_197),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_3),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_225),
.B(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_3),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_230),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_5),
.C(n_186),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_231),
.B(n_196),
.Y(n_254)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_253),
.B1(n_220),
.B2(n_201),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_236),
.A2(n_238),
.B1(n_175),
.B2(n_198),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_250),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_179),
.B1(n_197),
.B2(n_183),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_211),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_185),
.B(n_182),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_221),
.B1(n_231),
.B2(n_207),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_180),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_180),
.Y(n_245)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_188),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_246),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_171),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_188),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_238),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_228),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_258),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_215),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_259),
.A2(n_260),
.B1(n_236),
.B2(n_240),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_224),
.B1(n_204),
.B2(n_208),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_245),
.B(n_206),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_273),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_205),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_264),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_223),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_209),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_268),
.C(n_254),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_219),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_276),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_233),
.B(n_173),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_257),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_287),
.C(n_289),
.Y(n_293)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_267),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_281),
.B(n_282),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_263),
.B(n_243),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_244),
.B1(n_234),
.B2(n_246),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_283),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_265),
.B1(n_260),
.B2(n_259),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_253),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_289),
.C(n_277),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_269),
.B(n_250),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_292),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_294),
.B(n_284),
.Y(n_311)
);

NOR3xp33_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_199),
.C(n_209),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_300),
.Y(n_315)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_266),
.C(n_258),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_262),
.C(n_249),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_247),
.C(n_256),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_302),
.C(n_173),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_252),
.C(n_225),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_208),
.B(n_193),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_278),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_308),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_285),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_313),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_314),
.Y(n_323)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_283),
.B(n_287),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_280),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_298),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_293),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_310),
.B(n_304),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_307),
.A2(n_305),
.B(n_296),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_315),
.B(n_312),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_327),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_316),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_318),
.B(n_317),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_329),
.C(n_323),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_326),
.B(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_313),
.Y(n_333)
);


endmodule