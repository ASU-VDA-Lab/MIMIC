module fake_jpeg_25338_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_55),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_46),
.Y(n_52)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_56),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_41),
.B1(n_39),
.B2(n_45),
.Y(n_60)
);

HAxp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_0),
.CON(n_55),
.SN(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_15),
.B1(n_33),
.B2(n_32),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_65),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_49),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_79),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_49),
.B1(n_14),
.B2(n_16),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_80),
.B1(n_81),
.B2(n_6),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_2),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_13),
.B1(n_31),
.B2(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_3),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_12),
.C(n_24),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_4),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_5),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_92),
.B1(n_77),
.B2(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_6),
.Y(n_89)
);

OA21x2_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_7),
.B(n_9),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_94),
.C(n_95),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_100),
.B(n_7),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_83),
.C(n_10),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_99),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_21),
.C(n_11),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_92),
.B1(n_88),
.B2(n_90),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_98),
.B(n_20),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_17),
.Y(n_106)
);

AOI31xp67_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_22),
.A3(n_23),
.B(n_36),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_102),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_105),
.Y(n_110)
);


endmodule