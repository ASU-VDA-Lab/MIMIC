module fake_jpeg_30336_n_96 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_1),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_50),
.Y(n_56)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_55),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_40),
.B1(n_37),
.B2(n_41),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_10),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_71),
.B1(n_32),
.B2(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_63),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_11),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_12),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_73),
.B(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_19),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_64),
.B1(n_29),
.B2(n_30),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_23),
.Y(n_78)
);

NOR4xp25_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_28),
.C(n_31),
.D(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_81),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_84),
.C(n_81),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_80),
.C(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_80),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_82),
.C(n_86),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_87),
.Y(n_95)
);

BUFx24_ASAP7_75t_SL g96 ( 
.A(n_95),
.Y(n_96)
);


endmodule