module fake_jpeg_27012_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_50),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_31),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

BUFx2_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_34),
.Y(n_89)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_17),
.B1(n_28),
.B2(n_21),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_62),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_66),
.Y(n_95)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_40),
.B1(n_33),
.B2(n_37),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_48),
.B1(n_39),
.B2(n_41),
.Y(n_101)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_70),
.B(n_78),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_34),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_73),
.A2(n_39),
.B(n_38),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_46),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_40),
.B1(n_33),
.B2(n_57),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_103),
.B1(n_73),
.B2(n_84),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_48),
.B1(n_16),
.B2(n_18),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_108),
.B1(n_110),
.B2(n_30),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_0),
.B(n_1),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_58),
.B1(n_66),
.B2(n_81),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_48),
.B1(n_41),
.B2(n_27),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_18),
.B1(n_20),
.B2(n_26),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_26),
.B1(n_30),
.B2(n_20),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_13),
.C(n_14),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_12),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_14),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_15),
.C(n_32),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_116),
.B(n_46),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_102),
.B(n_115),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_27),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_122),
.B(n_130),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_89),
.B1(n_88),
.B2(n_82),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_124),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_69),
.B1(n_76),
.B2(n_80),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_112),
.B1(n_103),
.B2(n_104),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_132),
.B1(n_135),
.B2(n_144),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_90),
.B(n_73),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_69),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_134),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_117),
.B1(n_95),
.B2(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_93),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_64),
.B1(n_68),
.B2(n_58),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_100),
.B(n_64),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_139),
.Y(n_159)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_74),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_34),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_92),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_34),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_19),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_86),
.B1(n_85),
.B2(n_83),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_29),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_29),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_109),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_155),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_156),
.B(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_115),
.B1(n_102),
.B2(n_111),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_160),
.B1(n_125),
.B2(n_137),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_15),
.B(n_32),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_38),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_157),
.B(n_158),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_111),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_98),
.B1(n_107),
.B2(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_23),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_120),
.A2(n_98),
.B(n_19),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_97),
.C(n_109),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_0),
.C(n_1),
.Y(n_198)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_176),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_109),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_27),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_173),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_136),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_139),
.A2(n_25),
.B(n_1),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_175),
.A2(n_180),
.B(n_146),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_127),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_133),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_179),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_119),
.A2(n_25),
.B(n_83),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_119),
.B(n_147),
.C(n_142),
.D(n_121),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_192),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_180),
.B(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_145),
.B1(n_125),
.B2(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_188),
.A2(n_196),
.B1(n_199),
.B2(n_159),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_195),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_25),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_27),
.B1(n_23),
.B2(n_7),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_193),
.A2(n_205),
.B1(n_176),
.B2(n_174),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_198),
.C(n_202),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_171),
.B(n_11),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_23),
.B1(n_11),
.B2(n_10),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_153),
.B(n_10),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_197),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_149),
.A2(n_9),
.B1(n_8),
.B2(n_2),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_8),
.C(n_1),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_148),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_150),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_168),
.Y(n_223)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_224),
.B(n_185),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_162),
.B1(n_150),
.B2(n_172),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_186),
.B1(n_184),
.B2(n_164),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_158),
.C(n_152),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_229),
.C(n_192),
.Y(n_237)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_225),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_223),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_154),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_172),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_230),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_159),
.C(n_165),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_231),
.B(n_193),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_230),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_240),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_242),
.B1(n_219),
.B2(n_212),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_245),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_205),
.B1(n_189),
.B2(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_227),
.B(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_241),
.B(n_214),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_194),
.C(n_185),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_224),
.C(n_166),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_223),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_246),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_183),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_216),
.B(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_215),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_198),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_250),
.B(n_217),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_251),
.B(n_264),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

INVx11_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_255),
.B1(n_224),
.B2(n_211),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_211),
.B1(n_226),
.B2(n_222),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_229),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_247),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_245),
.B(n_218),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_266),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_237),
.C(n_232),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_272),
.C(n_273),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_275),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_236),
.C(n_241),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_236),
.C(n_244),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_210),
.B1(n_246),
.B2(n_233),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_239),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_240),
.B1(n_206),
.B2(n_213),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_277),
.A2(n_220),
.B1(n_255),
.B2(n_206),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_181),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_242),
.C(n_247),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_203),
.C(n_161),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_252),
.B(n_261),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_285),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_265),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_286),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_220),
.B(n_177),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_288),
.B(n_269),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_279),
.C(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_267),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_293),
.B(n_294),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_269),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_282),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_296),
.B(n_281),
.Y(n_301)
);

AND3x1_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_283),
.C(n_289),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_268),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_302),
.C(n_297),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_268),
.B(n_163),
.Y(n_302)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_304),
.C(n_299),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_298),
.C(n_163),
.Y(n_306)
);

OAI321xp33_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_307)
);

AOI31xp67_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_3),
.A3(n_4),
.B(n_5),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_4),
.B1(n_5),
.B2(n_227),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_309),
.Y(n_310)
);


endmodule