module real_jpeg_5186_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_2),
.B(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_2),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_2),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_2),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_2),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_2),
.B(n_273),
.Y(n_415)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_4),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_4),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_5),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_5),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_5),
.B(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_5),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_5),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_5),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_5),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_5),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_6),
.B(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_6),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_6),
.B(n_260),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_6),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_6),
.B(n_429),
.Y(n_428)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_7),
.Y(n_96)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_7),
.Y(n_215)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_9),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_9),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_9),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_9),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_9),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_9),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_10),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_10),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_10),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_10),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_10),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_11),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_11),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_11),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_11),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_11),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_11),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_11),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_11),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_12),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_12),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_12),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_12),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_12),
.B(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_13),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_14),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_15),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_15),
.B(n_169),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_15),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_15),
.B(n_74),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_15),
.B(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_15),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_15),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_15),
.B(n_375),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_183),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_181),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_158),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_19),
.B(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_100),
.C(n_118),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g473 ( 
.A(n_20),
.B(n_100),
.CI(n_118),
.CON(n_473),
.SN(n_473)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_58),
.B1(n_98),
.B2(n_99),
.Y(n_20)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_42),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_22),
.B(n_42),
.C(n_99),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.C(n_37),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_23),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.C(n_31),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_24),
.B(n_49),
.C(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_24),
.A2(n_31),
.B1(n_68),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_24),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_24),
.A2(n_127),
.B1(n_133),
.B2(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_24),
.A2(n_133),
.B1(n_381),
.B2(n_382),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_66),
.Y(n_65)
);

OR2x2_ASAP7_75t_SL g143 ( 
.A(n_25),
.B(n_144),
.Y(n_143)
);

OR2x2_ASAP7_75t_SL g176 ( 
.A(n_25),
.B(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_27),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_27),
.Y(n_131)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_29),
.B(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_30),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_31),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_31),
.B(n_60),
.C(n_65),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_31),
.B(n_317),
.C(n_321),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_31),
.A2(n_68),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_32),
.Y(n_239)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_32),
.Y(n_431)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_33),
.Y(n_408)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_33),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_35),
.A2(n_37),
.B1(n_38),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_35),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_37),
.A2(n_38),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_37),
.A2(n_38),
.B1(n_150),
.B2(n_151),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_38),
.B(n_136),
.C(n_150),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_40),
.Y(n_145)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_40),
.Y(n_257)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_43),
.B(n_49),
.C(n_52),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_52),
.B2(n_56),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_48),
.A2(n_49),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_51),
.Y(n_246)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_69),
.C(n_81),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_59),
.B(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_62),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_65),
.B1(n_109),
.B2(n_113),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_64),
.B(n_103),
.C(n_109),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_64),
.A2(n_65),
.B1(n_127),
.B2(n_292),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_65),
.B(n_127),
.C(n_204),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_67),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_69),
.B(n_81),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.C(n_76),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_70),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_70),
.A2(n_123),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_70),
.B(n_109),
.C(n_245),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_73),
.B(n_76),
.Y(n_124)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_80),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_80),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_97),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_92),
.C(n_93),
.Y(n_117)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g383 ( 
.A(n_86),
.Y(n_383)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_87),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_88),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_88),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_88),
.B(n_272),
.C(n_275),
.Y(n_284)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_114),
.B2(n_115),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_116),
.C(n_117),
.Y(n_160)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_109),
.A2(n_113),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_109),
.A2(n_113),
.B1(n_244),
.B2(n_248),
.Y(n_243)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_112),
.Y(n_372)
);

INVx5_ASAP7_75t_L g389 ( 
.A(n_112),
.Y(n_389)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_135),
.C(n_155),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_119),
.A2(n_120),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.C(n_130),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_126),
.Y(n_336)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_127),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g367 ( 
.A(n_129),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_130),
.B(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_133),
.B(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_135),
.B(n_155),
.Y(n_353)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_137),
.B(n_343),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.C(n_146),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_139),
.B(n_147),
.Y(n_287)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_143),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_143),
.Y(n_286)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_145),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_149),
.Y(n_274)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g475 ( 
.A(n_158),
.Y(n_475)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.CI(n_161),
.CON(n_158),
.SN(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_171),
.B2(n_180),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_176),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_176),
.B(n_220),
.C(n_225),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_471),
.B(n_474),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_346),
.B(n_355),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_330),
.B(n_345),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_307),
.B(n_329),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_188),
.B(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_279),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_189),
.B(n_279),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_242),
.C(n_267),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_190),
.B(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_216),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_191),
.B(n_217),
.C(n_228),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_203),
.C(n_207),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_192),
.B(n_325),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g476 ( 
.A(n_192),
.Y(n_476)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.CI(n_199),
.CON(n_192),
.SN(n_192)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_193),
.B(n_195),
.C(n_199),
.Y(n_278)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_198),
.Y(n_412)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_203),
.A2(n_207),
.B1(n_208),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_203),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_204),
.B(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_323)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_228),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_219)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_220),
.A2(n_227),
.B1(n_254),
.B2(n_255),
.Y(n_390)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_230),
.B(n_231),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_229),
.B(n_236),
.C(n_240),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_234),
.B(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_241),
.B(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_241),
.B(n_386),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_241),
.B(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_242),
.B(n_267),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_249),
.C(n_251),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_243),
.A2(n_249),
.B1(n_250),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_243),
.Y(n_312)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_251),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.C(n_263),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_252),
.A2(n_253),
.B1(n_458),
.B2(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_258),
.A2(n_259),
.B1(n_263),
.B2(n_264),
.Y(n_459)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_278),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_270),
.C(n_278),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_275),
.Y(n_270)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_282),
.C(n_306),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_293),
.B1(n_305),
.B2(n_306),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_289),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_285),
.C(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_294),
.B(n_296),
.C(n_297),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_300),
.B(n_302),
.C(n_341),
.Y(n_340)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_327),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_308),
.B(n_327),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.C(n_324),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_309),
.A2(n_310),
.B1(n_464),
.B2(n_465),
.Y(n_463)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_313),
.B(n_324),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.C(n_323),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_314),
.B(n_451),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_316),
.B(n_323),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_317),
.A2(n_318),
.B1(n_321),
.B2(n_322),
.Y(n_378)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_320),
.Y(n_375)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_331),
.B(n_346),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_333),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_347),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_333),
.B(n_347),
.Y(n_470)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_337),
.CI(n_344),
.CON(n_333),
.SN(n_333)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_340),
.C(n_342),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_348),
.B(n_350),
.C(n_352),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

OAI31xp33_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_467),
.A3(n_468),
.B(n_470),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_461),
.B(n_466),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_446),
.B(n_460),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_403),
.B(n_445),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_391),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_360),
.B(n_391),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_379),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_376),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_362),
.B(n_376),
.C(n_379),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_368),
.C(n_373),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_364),
.B1(n_368),
.B2(n_369),
.Y(n_393)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx8_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_373),
.B(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_384),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_380),
.B(n_455),
.C(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_390),
.Y(n_384)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.C(n_402),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_392),
.B(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_394),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_394),
.A2(n_402),
.B1(n_437),
.B2(n_443),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_399),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_398),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_402),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_439),
.B(n_444),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_424),
.B(n_438),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_413),
.B(n_423),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_421),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_421),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_416),
.B(n_420),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_415),
.B(n_416),
.Y(n_420)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_420),
.A2(n_426),
.B1(n_432),
.B2(n_433),
.Y(n_425)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_420),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_434),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_434),
.Y(n_438)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_426),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_427),
.A2(n_428),
.B(n_432),
.Y(n_440)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_435),
.A2(n_436),
.B(n_437),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_440),
.B(n_441),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_448),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_452),
.B2(n_453),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_454),
.C(n_457),
.Y(n_462)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_457),
.Y(n_453)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_462),
.B(n_463),
.Y(n_466)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_464),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_472),
.B(n_473),
.Y(n_474)
);

BUFx24_ASAP7_75t_SL g478 ( 
.A(n_473),
.Y(n_478)
);


endmodule