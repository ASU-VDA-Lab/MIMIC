module fake_jpeg_16879_n_333 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_41),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_1),
.Y(n_40)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_40),
.B(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_18),
.B(n_6),
.Y(n_41)
);

NAND2x1_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_6),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_43),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2x1_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_12),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_45),
.B(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_62),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_1),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_22),
.B1(n_32),
.B2(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_19),
.B(n_1),
.CON(n_56),
.SN(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_7),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_14),
.B(n_23),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_67),
.Y(n_96)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_27),
.B(n_3),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_24),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_76),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_77),
.B(n_98),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_78),
.A2(n_81),
.B1(n_102),
.B2(n_31),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_24),
.C(n_33),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_84),
.B(n_31),
.C(n_28),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_103),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_89),
.Y(n_154)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_18),
.Y(n_136)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_23),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_115),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_16),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_101),
.B(n_112),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_15),
.B1(n_32),
.B2(n_30),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

CKINVDCx9p33_ASAP7_75t_R g110 ( 
.A(n_42),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_43),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_25),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_40),
.B(n_25),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_116),
.B(n_11),
.Y(n_164)
);

CKINVDCx12_ASAP7_75t_R g117 ( 
.A(n_59),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_118),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_48),
.B1(n_50),
.B2(n_49),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_80),
.B1(n_87),
.B2(n_114),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_45),
.B1(n_16),
.B2(n_40),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_144),
.B1(n_149),
.B2(n_73),
.Y(n_167)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_38),
.B(n_35),
.C(n_17),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_161),
.B(n_104),
.Y(n_170)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_58),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_132),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_31),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_79),
.C(n_84),
.Y(n_174)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_74),
.B(n_33),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_148),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_136),
.B(n_164),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_38),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_156),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_35),
.B1(n_17),
.B2(n_11),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_146),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_151),
.B1(n_79),
.B2(n_75),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_9),
.B1(n_11),
.B2(n_7),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_91),
.A2(n_28),
.B1(n_31),
.B2(n_9),
.Y(n_151)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_153),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_70),
.B(n_28),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_90),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_94),
.B(n_3),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_9),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_104),
.A2(n_3),
.B(n_4),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_162),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_82),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_131),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_165),
.A2(n_167),
.B1(n_170),
.B2(n_186),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_166),
.A2(n_178),
.B1(n_199),
.B2(n_202),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_174),
.B(n_187),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_119),
.A2(n_80),
.B1(n_87),
.B2(n_106),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_176),
.A2(n_183),
.B1(n_192),
.B2(n_200),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_119),
.A2(n_105),
.B1(n_107),
.B2(n_97),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_73),
.B(n_107),
.C(n_85),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_141),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_193),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_97),
.B1(n_118),
.B2(n_4),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_171),
.B1(n_190),
.B2(n_181),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_132),
.A2(n_92),
.B1(n_71),
.B2(n_5),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_4),
.B(n_85),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_186),
.A2(n_195),
.B(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_129),
.A2(n_71),
.B1(n_121),
.B2(n_142),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_125),
.A2(n_121),
.B(n_126),
.Y(n_195)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_175),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_138),
.B(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_147),
.A2(n_152),
.B1(n_146),
.B2(n_130),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_127),
.A2(n_143),
.B1(n_124),
.B2(n_120),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_139),
.A2(n_150),
.B1(n_157),
.B2(n_159),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_203),
.A2(n_185),
.B(n_208),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_206),
.B1(n_215),
.B2(n_185),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_205),
.B(n_211),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_139),
.B1(n_157),
.B2(n_140),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_122),
.C(n_160),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_162),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_154),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_202),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_148),
.C(n_134),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_232),
.C(n_235),
.Y(n_238)
);

CKINVDCx10_ASAP7_75t_R g213 ( 
.A(n_201),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_137),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_214),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_217),
.A2(n_218),
.B(n_224),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_178),
.A2(n_166),
.B(n_179),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_226),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_170),
.A2(n_172),
.B(n_195),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_183),
.A2(n_176),
.B1(n_192),
.B2(n_165),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_191),
.B(n_168),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_222),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_169),
.B(n_175),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_232),
.C(n_199),
.Y(n_262)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_181),
.B(n_180),
.C(n_188),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_237),
.B(n_244),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_189),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_241),
.C(n_256),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_185),
.C(n_189),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_243),
.A2(n_259),
.B(n_260),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_225),
.B1(n_230),
.B2(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_231),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_251),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_203),
.B1(n_218),
.B2(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_204),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_206),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_261),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_235),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_213),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_238),
.C(n_248),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_209),
.A2(n_233),
.B(n_221),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_209),
.A2(n_216),
.B(n_234),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_273),
.C(n_276),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_245),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_264),
.B(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_252),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_240),
.C(n_262),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_269),
.B(n_250),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVxp33_ASAP7_75t_SL g274 ( 
.A(n_239),
.Y(n_274)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_242),
.C(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_245),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_278),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_253),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_251),
.C(n_257),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_280),
.C(n_283),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_243),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_258),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_282),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_241),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_239),
.B(n_246),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_260),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_254),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_250),
.B1(n_254),
.B2(n_259),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_288),
.A2(n_298),
.B1(n_296),
.B2(n_300),
.Y(n_310)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_271),
.C(n_276),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_294),
.C(n_266),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_279),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_SL g295 ( 
.A(n_267),
.B(n_280),
.C(n_269),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_270),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_270),
.A2(n_275),
.B(n_266),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_300),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_283),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_303),
.C(n_308),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_295),
.B(n_286),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_309),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_287),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_289),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_288),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_310),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_317),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_291),
.C(n_286),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_320),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_297),
.B(n_293),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_301),
.B(n_306),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_294),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_309),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_315),
.B(n_312),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_322),
.C(n_302),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_313),
.B(n_317),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_321),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);

AOI221xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_328),
.B1(n_313),
.B2(n_330),
.C(n_316),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_316),
.Y(n_333)
);


endmodule