module fake_jpeg_11805_n_392 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_392);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_392;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_49),
.Y(n_86)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_45),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_50),
.Y(n_129)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_61),
.Y(n_90)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_53),
.Y(n_128)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g104 ( 
.A(n_57),
.Y(n_104)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_69),
.Y(n_102)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_65),
.A2(n_81),
.B(n_82),
.Y(n_122)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_67),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_68),
.B(n_72),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_12),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_0),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_74),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_76),
.Y(n_117)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_40),
.Y(n_95)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_79),
.Y(n_119)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_84),
.Y(n_88)
);

BUFx24_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_28),
.B1(n_37),
.B2(n_18),
.Y(n_89)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_81),
.B(n_28),
.CON(n_85),
.SN(n_85)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_85),
.B(n_95),
.C(n_127),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_89),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_44),
.B(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_111),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_28),
.B1(n_41),
.B2(n_40),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_98),
.A2(n_99),
.B1(n_106),
.B2(n_114),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_34),
.B1(n_23),
.B2(n_31),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_34),
.B1(n_37),
.B2(n_30),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_115),
.B1(n_120),
.B2(n_130),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_34),
.B1(n_24),
.B2(n_30),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_105),
.B1(n_112),
.B2(n_131),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_42),
.B1(n_41),
.B2(n_20),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_23),
.B1(n_24),
.B2(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_42),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_36),
.B1(n_26),
.B2(n_20),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_47),
.A2(n_26),
.B1(n_24),
.B2(n_37),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_54),
.A2(n_37),
.B1(n_15),
.B2(n_29),
.Y(n_115)
);

NAND2x1_ASAP7_75t_L g118 ( 
.A(n_57),
.B(n_15),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_6),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_56),
.A2(n_37),
.B1(n_58),
.B2(n_67),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_1),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_127),
.A3(n_32),
.B1(n_29),
.B2(n_7),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_45),
.B(n_1),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_46),
.A2(n_32),
.B1(n_29),
.B2(n_3),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_65),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_82),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_150)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_136),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_85),
.A2(n_95),
.B1(n_128),
.B2(n_87),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_141),
.A2(n_173),
.B1(n_100),
.B2(n_93),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_118),
.Y(n_181)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_143),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_2),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_144),
.B(n_153),
.Y(n_194)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_174),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_6),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_160),
.C(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_107),
.B(n_7),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_156),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_116),
.B1(n_104),
.B2(n_108),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_151),
.Y(n_210)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_8),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_9),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_154),
.B(n_159),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_9),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_113),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_168),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_10),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_10),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_88),
.B(n_29),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_113),
.B(n_32),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_146),
.B(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_10),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_180),
.Y(n_200)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

AO22x1_ASAP7_75t_L g172 ( 
.A1(n_103),
.A2(n_32),
.B1(n_118),
.B2(n_87),
.Y(n_172)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_123),
.B1(n_100),
.B2(n_93),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_177),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_94),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_109),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_137),
.Y(n_217)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_179),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_104),
.B(n_32),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_181),
.A2(n_162),
.B1(n_134),
.B2(n_172),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_123),
.C(n_121),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_221),
.C(n_176),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_91),
.B1(n_116),
.B2(n_94),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_187),
.A2(n_201),
.B1(n_179),
.B2(n_135),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_188),
.A2(n_204),
.B1(n_176),
.B2(n_202),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_207),
.B1(n_214),
.B2(n_157),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_190),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_96),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_206),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_139),
.A2(n_121),
.B1(n_110),
.B2(n_108),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_110),
.B1(n_126),
.B2(n_133),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_126),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_152),
.A2(n_133),
.B1(n_138),
.B2(n_167),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_167),
.A2(n_165),
.B1(n_164),
.B2(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_217),
.B(n_183),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_147),
.A2(n_160),
.B(n_146),
.C(n_142),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_162),
.B(n_156),
.C(n_172),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_147),
.B(n_178),
.C(n_160),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_148),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_222),
.B(n_224),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_250),
.C(n_210),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_158),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_225),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_243),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_255),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_174),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_139),
.B1(n_157),
.B2(n_175),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_229),
.A2(n_231),
.B1(n_235),
.B2(n_212),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_177),
.B1(n_145),
.B2(n_171),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_252),
.B1(n_254),
.B2(n_210),
.Y(n_283)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_240),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_181),
.A2(n_143),
.B1(n_136),
.B2(n_151),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_176),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_236),
.Y(n_285)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

INVx11_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_242),
.C(n_245),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_185),
.B(n_186),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_190),
.A2(n_184),
.B(n_209),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_185),
.B(n_183),
.C(n_195),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_199),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_249),
.Y(n_258)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_209),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_219),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_203),
.A2(n_221),
.B(n_208),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_253),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_187),
.A2(n_201),
.B1(n_211),
.B2(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_197),
.A2(n_211),
.B1(n_208),
.B2(n_214),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_207),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_196),
.B(n_191),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_256),
.B(n_213),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_249),
.A2(n_191),
.B1(n_203),
.B2(n_193),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_257),
.A2(n_273),
.B1(n_270),
.B2(n_285),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_231),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_264),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_213),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_262),
.B(n_266),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_246),
.B(n_193),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_202),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_267),
.A2(n_270),
.B(n_283),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g270 ( 
.A1(n_227),
.A2(n_215),
.B(n_220),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_237),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_225),
.B(n_220),
.Y(n_275)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_245),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_282),
.B(n_253),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_226),
.B1(n_235),
.B2(n_248),
.Y(n_290)
);

NOR3xp33_ASAP7_75t_SL g284 ( 
.A(n_243),
.B(n_223),
.C(n_234),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_242),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_293),
.C(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_297),
.B1(n_273),
.B2(n_270),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_258),
.B(n_250),
.CI(n_230),
.CON(n_291),
.SN(n_291)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_268),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_241),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_294),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_230),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_264),
.A2(n_252),
.B1(n_232),
.B2(n_247),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_251),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_299),
.C(n_302),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_233),
.C(n_239),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_258),
.B(n_240),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_309),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_270),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_257),
.B(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_275),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_304),
.B(n_305),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_262),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_269),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_276),
.C(n_263),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_259),
.A2(n_260),
.B1(n_269),
.B2(n_261),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_308),
.A2(n_311),
.B1(n_276),
.B2(n_274),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_284),
.B(n_260),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_310),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_307),
.Y(n_312)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_321),
.Y(n_333)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_316),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_311),
.A2(n_267),
.B1(n_274),
.B2(n_265),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_318),
.A2(n_329),
.B1(n_297),
.B2(n_310),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_267),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_298),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_324),
.Y(n_344)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_323),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_265),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g349 ( 
.A1(n_327),
.A2(n_291),
.B(n_295),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_309),
.Y(n_340)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_332),
.Y(n_334)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_336),
.A2(n_342),
.B1(n_349),
.B2(n_315),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_268),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_337),
.B(n_339),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_320),
.B(n_287),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_314),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_325),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_324),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_318),
.A2(n_278),
.B1(n_286),
.B2(n_271),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_317),
.B(n_302),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_345),
.B(n_346),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_306),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_300),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_347),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_278),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_348),
.Y(n_355)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_344),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_338),
.A2(n_331),
.B1(n_316),
.B2(n_321),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_354),
.A2(n_333),
.B1(n_343),
.B2(n_313),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_314),
.C(n_322),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_357),
.B(n_358),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_326),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_362),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_360),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_338),
.B1(n_349),
.B2(n_348),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_333),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_291),
.B(n_313),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_334),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_368),
.Y(n_373)
);

OAI321xp33_ASAP7_75t_L g376 ( 
.A1(n_365),
.A2(n_350),
.A3(n_359),
.B1(n_355),
.B2(n_362),
.C(n_343),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_372),
.Y(n_379)
);

NOR2x1_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_340),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_361),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_281),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_350),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_375),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_366),
.A2(n_354),
.B1(n_355),
.B2(n_352),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_377),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_353),
.C(n_357),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_378),
.B(n_365),
.C(n_367),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_281),
.Y(n_380)
);

NOR2x1_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_371),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_385),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_R g382 ( 
.A(n_373),
.B(n_371),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_382),
.B(n_383),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_386),
.A2(n_387),
.B(n_368),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_384),
.B(n_377),
.C(n_379),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_388),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_389),
.A2(n_390),
.B(n_382),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_391),
.B(n_379),
.Y(n_392)
);


endmodule