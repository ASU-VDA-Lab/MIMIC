module fake_jpeg_8211_n_228 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_10),
.B(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_36),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_17),
.Y(n_50)
);

CKINVDCx9p33_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_27),
.B1(n_18),
.B2(n_15),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_48),
.B1(n_52),
.B2(n_21),
.Y(n_67)
);

AO22x1_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_29),
.B1(n_37),
.B2(n_31),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_30),
.B(n_26),
.C(n_24),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_31),
.B1(n_35),
.B2(n_39),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_27),
.B1(n_18),
.B2(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_16),
.B1(n_24),
.B2(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_14),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_18),
.B1(n_27),
.B2(n_20),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_75),
.B1(n_42),
.B2(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_65),
.B1(n_43),
.B2(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_36),
.B1(n_34),
.B2(n_33),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_57),
.B1(n_45),
.B2(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_33),
.B1(n_47),
.B2(n_51),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_47),
.B1(n_54),
.B2(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_30),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_43),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_81),
.B(n_92),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_86),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_47),
.B1(n_51),
.B2(n_56),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_67),
.B1(n_70),
.B2(n_60),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_58),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_56),
.B1(n_45),
.B2(n_25),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_21),
.B1(n_26),
.B2(n_22),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_91),
.B1(n_61),
.B2(n_65),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_46),
.B1(n_14),
.B2(n_19),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_60),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_76),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_112),
.B1(n_92),
.B2(n_76),
.Y(n_131)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_106),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_73),
.B(n_60),
.C(n_72),
.D(n_66),
.Y(n_99)
);

XOR2x2_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_60),
.B1(n_64),
.B2(n_62),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_108),
.B1(n_78),
.B2(n_86),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_107),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_60),
.B1(n_75),
.B2(n_16),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_92),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_91),
.B1(n_90),
.B2(n_85),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_17),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_89),
.C(n_80),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_121),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_123),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_105),
.B(n_108),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_127),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_89),
.C(n_87),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_126),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_79),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_101),
.B1(n_22),
.B2(n_41),
.C(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_110),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_96),
.B(n_99),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_120),
.B1(n_130),
.B2(n_115),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_128),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_103),
.B(n_97),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_123),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_120),
.Y(n_156)
);

OAI22x1_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_63),
.B1(n_41),
.B2(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_148),
.B(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_8),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_126),
.C(n_119),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_164),
.C(n_165),
.Y(n_172)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_139),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_138),
.B1(n_148),
.B2(n_141),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_144),
.B(n_147),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_166),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_129),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_167),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_117),
.C(n_127),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_117),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_41),
.C(n_63),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_178),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_140),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_132),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_134),
.B1(n_137),
.B2(n_9),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_182),
.B1(n_152),
.B2(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_184),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_164),
.B1(n_155),
.B2(n_151),
.Y(n_184)
);

NAND4xp25_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_41),
.C(n_156),
.D(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_0),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_0),
.C(n_1),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_190),
.C(n_185),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_0),
.C(n_1),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_193),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_6),
.CI(n_12),
.CON(n_193),
.SN(n_193)
);

XOR2x2_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_176),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_196),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_172),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_169),
.B(n_176),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_202),
.C(n_204),
.Y(n_208)
);

OAI21x1_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_169),
.B(n_6),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_10),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_9),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_193),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_5),
.C(n_12),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_194),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_211),
.B(n_200),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_4),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_187),
.C(n_189),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_212),
.C(n_204),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_193),
.C(n_5),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_4),
.C(n_11),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_3),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_3),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_217),
.A2(n_218),
.B(n_209),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_11),
.B(n_13),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_4),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.C(n_221),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_219),
.C(n_13),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_1),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_2),
.Y(n_228)
);


endmodule