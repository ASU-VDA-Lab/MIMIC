module fake_jpeg_29771_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_59),
.Y(n_69)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_14),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_13),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_27),
.B(n_0),
.C(n_1),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_12),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_19),
.B(n_23),
.C(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_66),
.B(n_111),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_39),
.B1(n_38),
.B2(n_35),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_67),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_134)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_94),
.B1(n_97),
.B2(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_82),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_87),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_32),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_88),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_41),
.A2(n_27),
.B1(n_39),
.B2(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_89),
.A2(n_100),
.B1(n_2),
.B2(n_4),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_30),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_90),
.Y(n_133)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_39),
.B(n_38),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_43),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_35),
.B1(n_36),
.B2(n_32),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_45),
.B(n_23),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_101),
.B(n_102),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_22),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_62),
.A2(n_35),
.B1(n_33),
.B2(n_31),
.Y(n_104)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_52),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_31),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_35),
.B1(n_25),
.B2(n_22),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_25),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_128),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_66),
.A2(n_21),
.B1(n_12),
.B2(n_11),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_127),
.B1(n_140),
.B2(n_89),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_21),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_21),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_136),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_104),
.B1(n_113),
.B2(n_79),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_21),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_1),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_7),
.B(n_8),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_147),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_150),
.A2(n_157),
.B1(n_160),
.B2(n_137),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_175),
.Y(n_188)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_153),
.B(n_154),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_69),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_114),
.A2(n_64),
.B1(n_72),
.B2(n_92),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_80),
.B1(n_105),
.B2(n_107),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_177),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_80),
.B1(n_105),
.B2(n_107),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_128),
.A2(n_97),
.B1(n_110),
.B2(n_72),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_70),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_173),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_70),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_172),
.C(n_177),
.Y(n_210)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_92),
.B(n_71),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_176),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_68),
.C(n_64),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_84),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_84),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_139),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_110),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_99),
.B1(n_68),
.B2(n_95),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_85),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_141),
.A2(n_85),
.B(n_95),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_98),
.B(n_116),
.C(n_7),
.Y(n_213)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_182),
.A2(n_191),
.B1(n_201),
.B2(n_204),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_192),
.B1(n_205),
.B2(n_211),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_141),
.B1(n_131),
.B2(n_119),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_150),
.A2(n_131),
.B1(n_103),
.B2(n_109),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_135),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_198),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_148),
.B(n_168),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_197),
.A2(n_213),
.B(n_146),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_121),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_121),
.B1(n_109),
.B2(n_142),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_145),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_115),
.B1(n_130),
.B2(n_120),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_157),
.A2(n_149),
.B1(n_172),
.B2(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_130),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_115),
.B1(n_120),
.B2(n_98),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_116),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_158),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_221),
.Y(n_250)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_202),
.A2(n_163),
.A3(n_170),
.B1(n_167),
.B2(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_187),
.A2(n_163),
.B(n_176),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_207),
.B(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_170),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_222),
.B(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_167),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_152),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_226),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_184),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_164),
.C(n_161),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_10),
.C(n_8),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_156),
.B(n_8),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_233),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_191),
.B(n_9),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_156),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

OAI321xp33_ASAP7_75t_L g236 ( 
.A1(n_188),
.A2(n_7),
.A3(n_8),
.B1(n_10),
.B2(n_197),
.C(n_205),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_192),
.B1(n_211),
.B2(n_189),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_244),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_241),
.A2(n_242),
.B1(n_237),
.B2(n_225),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_187),
.B1(n_207),
.B2(n_182),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_201),
.B1(n_210),
.B2(n_188),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_253),
.B1(n_229),
.B2(n_216),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_193),
.Y(n_244)
);

OAI322xp33_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_214),
.A3(n_212),
.B1(n_190),
.B2(n_194),
.C1(n_203),
.C2(n_200),
.Y(n_248)
);

AOI321xp33_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_217),
.A3(n_221),
.B1(n_236),
.B2(n_225),
.C(n_231),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_183),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_256),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_183),
.B1(n_196),
.B2(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_249),
.A2(n_238),
.B1(n_219),
.B2(n_215),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_259),
.B1(n_265),
.B2(n_266),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_252),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_240),
.B(n_220),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_264),
.Y(n_274)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_226),
.B(n_218),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_222),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_270),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_233),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_250),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_253),
.B1(n_245),
.B2(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_251),
.C(n_256),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_275),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_243),
.C(n_242),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_278),
.C(n_250),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_239),
.B(n_245),
.C(n_217),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_230),
.B(n_264),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_SL g283 ( 
.A(n_268),
.B(n_246),
.C(n_223),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_223),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_241),
.B1(n_254),
.B2(n_267),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_262),
.C(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_289),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_288),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_262),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_265),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_295),
.B1(n_278),
.B2(n_274),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_293),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_246),
.B1(n_254),
.B2(n_238),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

AOI31xp67_ASAP7_75t_SL g298 ( 
.A1(n_287),
.A2(n_283),
.A3(n_278),
.B(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_301),
.B1(n_297),
.B2(n_302),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_263),
.B(n_218),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_289),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_306),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_299),
.C(n_286),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_285),
.C(n_234),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_215),
.B1(n_232),
.B2(n_307),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_288),
.B1(n_232),
.B2(n_235),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_304),
.C(n_306),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_311),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_312),
.C(n_309),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_309),
.Y(n_315)
);


endmodule