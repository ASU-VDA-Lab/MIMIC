module fake_aes_9338_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
BUFx3_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
AND2x4_ASAP7_75t_L g5 ( .A(n_4), .B(n_0), .Y(n_5) );
NAND3xp33_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .C(n_1), .Y(n_6) );
OR2x2_ASAP7_75t_L g7 ( .A(n_5), .B(n_4), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
AOI221xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_3), .B1(n_4), .B2(n_6), .C(n_0), .Y(n_9) );
AOI21xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_3), .B(n_4), .Y(n_10) );
OAI222xp33_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_0), .B1(n_1), .B2(n_2), .C1(n_3), .C2(n_4), .Y(n_11) );
endmodule