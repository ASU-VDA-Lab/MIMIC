module fake_jpeg_24776_n_136 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_11),
.Y(n_38)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_13),
.B1(n_16),
.B2(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_38),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_16),
.B(n_21),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_14),
.B1(n_19),
.B2(n_17),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_46),
.B1(n_14),
.B2(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_13),
.B1(n_24),
.B2(n_30),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_50),
.B1(n_52),
.B2(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_16),
.B1(n_20),
.B2(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_11),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_51),
.Y(n_55)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_59),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_54),
.B(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_64),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_34),
.C(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_71),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_74),
.B(n_60),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_35),
.C(n_12),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_65),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_66),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_70),
.B1(n_67),
.B2(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_88),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_33),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_35),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_87),
.A2(n_79),
.B1(n_85),
.B2(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_50),
.B1(n_45),
.B2(n_35),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_89),
.B(n_9),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_7),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_45),
.CI(n_33),
.CON(n_105),
.SN(n_105)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_99),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_78),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_107),
.C(n_93),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_108),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_3),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_1),
.C(n_2),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_98),
.C(n_95),
.Y(n_116)
);

NAND4xp25_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_105),
.C(n_101),
.D(n_109),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_3),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_115),
.A2(n_107),
.B(n_102),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_4),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_124),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_126),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_4),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_118),
.C(n_4),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.C(n_128),
.Y(n_134)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_134),
.B(n_135),
.CI(n_5),
.CON(n_136),
.SN(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_130),
.C(n_5),
.Y(n_135)
);


endmodule