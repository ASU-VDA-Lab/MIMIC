module fake_jpeg_213_n_695 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_695);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_695;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_60),
.Y(n_171)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g217 ( 
.A(n_61),
.Y(n_217)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_64),
.Y(n_202)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_65),
.Y(n_139)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_67),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_68),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_70),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_71),
.B(n_80),
.Y(n_159)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_77),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_79),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_22),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_37),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_83),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_24),
.B(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_84),
.B(n_89),
.Y(n_170)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_19),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_108),
.Y(n_140)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_88),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_90),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_91),
.B(n_93),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_22),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_41),
.B(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_98),
.B(n_103),
.Y(n_201)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_100),
.Y(n_227)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_25),
.B(n_18),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_25),
.B(n_17),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_113),
.B(n_120),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_26),
.B(n_17),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_121),
.B(n_127),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_21),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_50),
.Y(n_129)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_129),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_49),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_131),
.B(n_31),
.Y(n_222)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_136),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_138),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_142),
.B(n_161),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_78),
.A2(n_30),
.B1(n_54),
.B2(n_47),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_149),
.A2(n_152),
.B1(n_167),
.B2(n_49),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_82),
.A2(n_30),
.B1(n_50),
.B2(n_54),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_158),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_74),
.A2(n_27),
.B1(n_56),
.B2(n_55),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_160),
.A2(n_193),
.B1(n_107),
.B2(n_21),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_96),
.A2(n_57),
.B1(n_47),
.B2(n_40),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_126),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_168),
.B(n_188),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_129),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_173),
.Y(n_292)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_177),
.Y(n_289)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_75),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_184),
.Y(n_306)
);

BUFx8_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

CKINVDCx6p67_ASAP7_75t_R g312 ( 
.A(n_185),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_66),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_119),
.A2(n_26),
.B1(n_56),
.B2(n_55),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_87),
.A2(n_57),
.B(n_32),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_196),
.B(n_224),
.Y(n_266)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_83),
.Y(n_199)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_SL g203 ( 
.A(n_81),
.B(n_36),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_203),
.B(n_2),
.Y(n_276)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_208),
.Y(n_304)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_92),
.B(n_36),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_214),
.B(n_110),
.Y(n_260)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_67),
.Y(n_216)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_69),
.Y(n_218)
);

BUFx8_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_94),
.A2(n_53),
.B1(n_27),
.B2(n_45),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_220),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_222),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_77),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_97),
.Y(n_226)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_101),
.Y(n_228)
);

INVx3_ASAP7_75t_SL g245 ( 
.A(n_228),
.Y(n_245)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_102),
.Y(n_229)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_39),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_231),
.B(n_273),
.Y(n_319)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_233),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_166),
.A2(n_40),
.B1(n_39),
.B2(n_35),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_234),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_195),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_237),
.B(n_256),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_53),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_240),
.B(n_241),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_45),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_242),
.A2(n_249),
.B1(n_271),
.B2(n_298),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_159),
.B(n_35),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_243),
.B(n_250),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_244),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_246),
.Y(n_344)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_247),
.Y(n_348)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_144),
.Y(n_248)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_248),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_195),
.A2(n_31),
.B1(n_29),
.B2(n_222),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_159),
.B(n_204),
.Y(n_250)
);

BUFx24_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

BUFx2_ASAP7_75t_SL g318 ( 
.A(n_251),
.Y(n_318)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_252),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_149),
.A2(n_116),
.B1(n_115),
.B2(n_114),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_254),
.A2(n_279),
.B1(n_217),
.B2(n_189),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_204),
.B(n_29),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_255),
.B(n_269),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_184),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_257),
.Y(n_329)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_260),
.B(n_263),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_17),
.Y(n_263)
);

CKINVDCx12_ASAP7_75t_R g264 ( 
.A(n_133),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_264),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_140),
.B(n_16),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_265),
.B(n_270),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_133),
.Y(n_267)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_197),
.Y(n_268)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_170),
.B(n_16),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_202),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_223),
.Y(n_272)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_272),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_170),
.B(n_0),
.Y(n_273)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_151),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_274),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_227),
.B(n_0),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_275),
.B(n_300),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_SL g369 ( 
.A(n_276),
.B(n_143),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_152),
.Y(n_278)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_167),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_151),
.B(n_138),
.Y(n_280)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_280),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_173),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_281),
.Y(n_349)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_139),
.Y(n_283)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_139),
.Y(n_284)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_178),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_285),
.A2(n_296),
.B1(n_301),
.B2(n_215),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_141),
.Y(n_291)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_147),
.Y(n_294)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_294),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_134),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_295)
);

NOR2x1_ASAP7_75t_L g376 ( 
.A(n_295),
.B(n_297),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_137),
.B(n_10),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_148),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_136),
.B(n_11),
.Y(n_299)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_299),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_153),
.B(n_14),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_200),
.A2(n_14),
.B1(n_15),
.B2(n_191),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_206),
.Y(n_302)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_155),
.Y(n_303)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_303),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_171),
.B(n_15),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_305),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_156),
.B(n_15),
.Y(n_307)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_186),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_313),
.Y(n_357)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_210),
.Y(n_310)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_310),
.Y(n_375)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_175),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_215),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_175),
.Y(n_314)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_316),
.A2(n_306),
.B1(n_293),
.B2(n_284),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_266),
.A2(n_221),
.B1(n_135),
.B2(n_145),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_317),
.A2(n_325),
.B1(n_330),
.B2(n_333),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_231),
.A2(n_150),
.B1(n_181),
.B2(n_205),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_270),
.A2(n_186),
.B1(n_164),
.B2(n_163),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_278),
.A2(n_221),
.B1(n_213),
.B2(n_211),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_273),
.B(n_308),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_371),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_296),
.A2(n_174),
.B1(n_213),
.B2(n_211),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_341),
.A2(n_342),
.B1(n_362),
.B2(n_258),
.Y(n_411)
);

OA22x2_ASAP7_75t_L g345 ( 
.A1(n_276),
.A2(n_176),
.B1(n_192),
.B2(n_154),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_283),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_254),
.A2(n_225),
.B1(n_198),
.B2(n_217),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_347),
.Y(n_410)
);

AOI32xp33_ASAP7_75t_L g350 ( 
.A1(n_276),
.A2(n_179),
.A3(n_157),
.B1(n_172),
.B2(n_165),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_306),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_238),
.B(n_212),
.C(n_169),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_353),
.B(n_289),
.C(n_245),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_360),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_292),
.A2(n_146),
.B1(n_194),
.B2(n_218),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_361),
.A2(n_365),
.B1(n_342),
.B2(n_327),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_262),
.A2(n_158),
.B1(n_143),
.B2(n_162),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_236),
.Y(n_363)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_363),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_279),
.A2(n_143),
.B1(n_162),
.B2(n_295),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_312),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_239),
.B(n_162),
.Y(n_371)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_379),
.Y(n_428)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_381),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_321),
.Y(n_382)
);

NAND2xp33_ASAP7_75t_SL g467 ( 
.A(n_382),
.B(n_396),
.Y(n_467)
);

OAI22xp33_ASAP7_75t_SL g450 ( 
.A1(n_383),
.A2(n_424),
.B1(n_425),
.B2(n_251),
.Y(n_450)
);

INVx13_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_384),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_385),
.B(n_411),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_323),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_386),
.B(n_399),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_327),
.A2(n_312),
.B1(n_293),
.B2(n_302),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_387),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_319),
.B(n_288),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_388),
.B(n_407),
.Y(n_439)
);

INVx13_ASAP7_75t_L g389 ( 
.A(n_337),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_389),
.Y(n_452)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_363),
.Y(n_390)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_390),
.Y(n_438)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_391),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_351),
.A2(n_314),
.B1(n_311),
.B2(n_233),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_392),
.A2(n_414),
.B1(n_333),
.B2(n_368),
.Y(n_432)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

INVx13_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g461 ( 
.A(n_395),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_319),
.B(n_253),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_397),
.B(n_413),
.Y(n_449)
);

INVx13_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_398),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_340),
.B(n_294),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_400),
.B(n_401),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_267),
.Y(n_401)
);

INVx13_ASAP7_75t_L g402 ( 
.A(n_338),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_402),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_358),
.B(n_267),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_403),
.B(n_404),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_357),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_405),
.A2(n_415),
.B1(n_427),
.B2(n_344),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_289),
.Y(n_407)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_409),
.Y(n_453)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_412),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_351),
.A2(n_310),
.B1(n_252),
.B2(n_247),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_376),
.A2(n_303),
.B(n_282),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_416),
.A2(n_396),
.B(n_422),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_282),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_417),
.A2(n_396),
.B(n_369),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_354),
.B(n_290),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_419),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_339),
.B(n_232),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_232),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_421),
.Y(n_448)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_375),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_357),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_426),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_322),
.B(n_353),
.C(n_371),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_397),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_374),
.A2(n_258),
.B1(n_290),
.B2(n_304),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_374),
.A2(n_304),
.B1(n_235),
.B2(n_286),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_320),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_410),
.A2(n_317),
.B1(n_370),
.B2(n_326),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_430),
.A2(n_434),
.B(n_444),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_432),
.A2(n_435),
.B1(n_440),
.B2(n_446),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_433),
.B(n_394),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_416),
.A2(n_365),
.B(n_349),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_405),
.A2(n_359),
.B1(n_343),
.B2(n_368),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_417),
.A2(n_368),
.B1(n_375),
.B2(n_348),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_417),
.A2(n_345),
.B1(n_367),
.B2(n_352),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_443),
.A2(n_469),
.B1(n_392),
.B2(n_399),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_410),
.A2(n_286),
.B(n_235),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_406),
.A2(n_348),
.B1(n_334),
.B2(n_335),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_450),
.A2(n_394),
.B1(n_408),
.B2(n_409),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_406),
.A2(n_385),
.B1(n_380),
.B2(n_414),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_455),
.A2(n_456),
.B1(n_457),
.B2(n_468),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_380),
.A2(n_334),
.B1(n_335),
.B2(n_244),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_420),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_423),
.B(n_345),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_413),
.Y(n_474)
);

OAI32xp33_ASAP7_75t_L g464 ( 
.A1(n_385),
.A2(n_345),
.A3(n_356),
.B1(n_331),
.B2(n_329),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_378),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_466),
.A2(n_426),
.B(n_419),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_411),
.A2(n_328),
.B1(n_346),
.B2(n_344),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_388),
.A2(n_287),
.B1(n_268),
.B2(n_246),
.Y(n_469)
);

BUFx12f_ASAP7_75t_L g470 ( 
.A(n_441),
.Y(n_470)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_470),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_471),
.B(n_489),
.C(n_440),
.Y(n_533)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_428),
.Y(n_472)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_472),
.Y(n_510)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_465),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_473),
.B(n_490),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_474),
.B(n_449),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_404),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_498),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_477),
.A2(n_486),
.B(n_487),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_478),
.B(n_437),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_455),
.A2(n_386),
.B1(n_378),
.B2(n_390),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_479),
.A2(n_456),
.B1(n_469),
.B2(n_460),
.Y(n_534)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_480),
.Y(n_511)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_481),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_412),
.Y(n_482)
);

INVxp33_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_483),
.Y(n_541)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_429),
.Y(n_484)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_484),
.Y(n_537)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_438),
.Y(n_485)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_485),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_466),
.A2(n_381),
.B(n_379),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_433),
.A2(n_382),
.B(n_391),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_488),
.A2(n_504),
.B(n_444),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_427),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_454),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_452),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_491),
.B(n_492),
.Y(n_517)
);

BUFx12f_ASAP7_75t_L g492 ( 
.A(n_441),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_SL g493 ( 
.A(n_443),
.B(n_395),
.C(n_398),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_493),
.B(n_501),
.Y(n_528)
);

BUFx12_ASAP7_75t_L g494 ( 
.A(n_461),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_494),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_453),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_495),
.Y(n_526)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_431),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_496),
.Y(n_535)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_438),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_448),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_507),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_451),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_500),
.B(n_502),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_442),
.B(n_373),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_451),
.Y(n_502)
);

OAI21xp33_ASAP7_75t_L g544 ( 
.A1(n_503),
.A2(n_436),
.B(n_463),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_434),
.A2(n_235),
.B(n_389),
.Y(n_504)
);

INVx11_ASAP7_75t_L g506 ( 
.A(n_460),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_506),
.Y(n_543)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_442),
.B(n_439),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_508),
.B(n_421),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_486),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_509),
.B(n_545),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_449),
.Y(n_518)
);

MAJx2_ASAP7_75t_L g562 ( 
.A(n_518),
.B(n_527),
.C(n_533),
.Y(n_562)
);

INVxp33_ASAP7_75t_L g572 ( 
.A(n_520),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_499),
.A2(n_435),
.B1(n_437),
.B2(n_468),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_521),
.A2(n_532),
.B1(n_540),
.B2(n_447),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_522),
.A2(n_534),
.B1(n_488),
.B2(n_493),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_439),
.Y(n_523)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_523),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_475),
.A2(n_503),
.B(n_504),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_524),
.A2(n_544),
.B(n_487),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_479),
.B(n_437),
.Y(n_529)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_529),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_483),
.B(n_464),
.Y(n_530)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_530),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_475),
.A2(n_467),
.B(n_445),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_531),
.A2(n_524),
.B(n_520),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_478),
.A2(n_430),
.B1(n_432),
.B2(n_459),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_483),
.A2(n_446),
.B1(n_445),
.B2(n_436),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_489),
.B(n_463),
.C(n_453),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_471),
.C(n_485),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_498),
.B(n_431),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_546),
.B(n_496),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_547),
.A2(n_564),
.B(n_526),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_549),
.B(n_553),
.Y(n_586)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_551),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_527),
.B(n_477),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_552),
.B(n_556),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_533),
.B(n_476),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_518),
.B(n_542),
.C(n_519),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_554),
.B(n_567),
.C(n_569),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_538),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_555),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_519),
.B(n_497),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_557),
.A2(n_543),
.B1(n_526),
.B2(n_537),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_523),
.B(n_505),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_558),
.B(n_563),
.Y(n_587)
);

FAx1_ASAP7_75t_SL g559 ( 
.A(n_516),
.B(n_484),
.CI(n_481),
.CON(n_559),
.SN(n_559)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_559),
.A2(n_566),
.B1(n_534),
.B2(n_543),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_515),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_560),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_561),
.A2(n_540),
.B(n_512),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_516),
.B(n_472),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_541),
.A2(n_447),
.B(n_506),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_515),
.B(n_529),
.C(n_532),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_525),
.B(n_393),
.Y(n_568)
);

OA21x2_ASAP7_75t_SL g593 ( 
.A1(n_568),
.A2(n_571),
.B(n_511),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_522),
.B(n_541),
.C(n_521),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_522),
.B(n_366),
.C(n_373),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_570),
.B(n_510),
.C(n_514),
.Y(n_592)
);

NOR3xp33_ASAP7_75t_SL g571 ( 
.A(n_528),
.B(n_494),
.C(n_402),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_530),
.B(n_366),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_578),
.Y(n_588)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_536),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_574),
.Y(n_600)
);

CKINVDCx16_ASAP7_75t_R g575 ( 
.A(n_517),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_575),
.A2(n_579),
.B1(n_512),
.B2(n_511),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_SL g576 ( 
.A(n_531),
.B(n_494),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_SL g584 ( 
.A(n_576),
.B(n_545),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_528),
.B(n_324),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_513),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_580),
.B(n_581),
.Y(n_623)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_582),
.Y(n_620)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_583),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_584),
.B(n_597),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_589),
.A2(n_596),
.B1(n_603),
.B2(n_566),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_554),
.B(n_537),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_591),
.B(n_592),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_593),
.B(n_571),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_549),
.B(n_535),
.C(n_539),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_594),
.B(n_601),
.C(n_602),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_558),
.A2(n_514),
.B1(n_510),
.B2(n_539),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_SL g597 ( 
.A(n_552),
.B(n_562),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_SL g599 ( 
.A(n_562),
.B(n_536),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_606),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_553),
.B(n_535),
.C(n_408),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_556),
.B(n_324),
.C(n_320),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_548),
.A2(n_415),
.B1(n_364),
.B2(n_492),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_578),
.B(n_569),
.C(n_567),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_415),
.C(n_332),
.Y(n_626)
);

XNOR2xp5_ASAP7_75t_SL g606 ( 
.A(n_576),
.B(n_384),
.Y(n_606)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_608),
.Y(n_629)
);

AOI21xp33_ASAP7_75t_L g609 ( 
.A1(n_604),
.A2(n_565),
.B(n_547),
.Y(n_609)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_609),
.Y(n_640)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_611),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_589),
.A2(n_572),
.B(n_550),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_613),
.B(n_616),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_595),
.B(n_563),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_615),
.B(n_619),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_587),
.A2(n_572),
.B(n_577),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_594),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_617),
.Y(n_644)
);

CKINVDCx16_ASAP7_75t_R g619 ( 
.A(n_592),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_600),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_621),
.B(n_620),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_598),
.A2(n_564),
.B1(n_559),
.B2(n_570),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_622),
.B(n_626),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_591),
.B(n_573),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_624),
.B(n_627),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_587),
.B(n_559),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_625),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_584),
.A2(n_492),
.B(n_470),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_601),
.B(n_492),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_588),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_618),
.B(n_590),
.C(n_605),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_631),
.B(n_632),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_607),
.C(n_617),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_623),
.A2(n_608),
.B(n_613),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_635),
.A2(n_623),
.B(n_625),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_612),
.A2(n_602),
.B1(n_606),
.B2(n_585),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_636),
.A2(n_470),
.B1(n_261),
.B2(n_277),
.Y(n_656)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_637),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g657 ( 
.A(n_639),
.B(n_642),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_607),
.B(n_586),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_641),
.B(n_646),
.Y(n_663)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_628),
.B(n_585),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_628),
.B(n_599),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_643),
.B(n_277),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_626),
.B(n_590),
.C(n_586),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_632),
.B(n_612),
.C(n_624),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_648),
.B(n_651),
.Y(n_667)
);

AOI21x1_ASAP7_75t_L g671 ( 
.A1(n_649),
.A2(n_650),
.B(n_647),
.Y(n_671)
);

NOR2xp67_ASAP7_75t_L g650 ( 
.A(n_640),
.B(n_597),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_631),
.B(n_616),
.C(n_588),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_SL g652 ( 
.A1(n_629),
.A2(n_627),
.B1(n_614),
.B2(n_610),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_652),
.B(n_653),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_646),
.B(n_610),
.C(n_614),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_644),
.B(n_470),
.C(n_332),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_655),
.B(n_658),
.C(n_662),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_656),
.B(n_643),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_633),
.B(n_236),
.C(n_261),
.Y(n_658)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_659),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_634),
.A2(n_245),
.B(n_251),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_661),
.A2(n_645),
.B(n_639),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_630),
.B(n_274),
.C(n_642),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_SL g665 ( 
.A1(n_660),
.A2(n_638),
.B(n_634),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_665),
.A2(n_671),
.B(n_657),
.Y(n_682)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_655),
.Y(n_668)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_668),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_669),
.B(n_670),
.Y(n_676)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_658),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g673 ( 
.A(n_651),
.B(n_645),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_673),
.B(n_662),
.Y(n_678)
);

INVx6_ASAP7_75t_L g674 ( 
.A(n_663),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_674),
.B(n_675),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_678),
.B(n_679),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_667),
.B(n_654),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_674),
.B(n_648),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_680),
.B(n_681),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_672),
.B(n_653),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_682),
.A2(n_665),
.B(n_673),
.Y(n_684)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_684),
.Y(n_690)
);

XOR2xp5_ASAP7_75t_L g685 ( 
.A(n_677),
.B(n_657),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_685),
.B(n_686),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_SL g686 ( 
.A1(n_683),
.A2(n_664),
.B(n_669),
.C(n_636),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_690),
.A2(n_687),
.B(n_688),
.C(n_682),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_691),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_692),
.A2(n_689),
.B1(n_676),
.B2(n_656),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_693),
.B(n_666),
.Y(n_694)
);

XNOR2xp5_ASAP7_75t_L g695 ( 
.A(n_694),
.B(n_661),
.Y(n_695)
);


endmodule