module real_jpeg_13240_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_3),
.A2(n_62),
.B1(n_65),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_78),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_4),
.A2(n_62),
.B1(n_65),
.B2(n_80),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_4),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_26),
.B1(n_30),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_5),
.A2(n_51),
.B1(n_62),
.B2(n_65),
.Y(n_161)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_7),
.A2(n_26),
.B1(n_30),
.B2(n_56),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_7),
.A2(n_56),
.B1(n_62),
.B2(n_65),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_26),
.B1(n_30),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_9),
.A2(n_53),
.B1(n_62),
.B2(n_65),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_11),
.A2(n_32),
.B(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_11),
.B(n_91),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_37),
.B1(n_48),
.B2(n_49),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_11),
.A2(n_49),
.B(n_59),
.C(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_11),
.B(n_89),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_11),
.B(n_76),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_11),
.B(n_68),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_11),
.A2(n_30),
.B(n_43),
.C(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_12),
.A2(n_48),
.B1(n_49),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_12),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_12),
.A2(n_62),
.B1(n_65),
.B2(n_67),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_13),
.A2(n_26),
.B1(n_30),
.B2(n_39),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_13),
.A2(n_39),
.B1(n_48),
.B2(n_49),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_13),
.A2(n_39),
.B1(n_62),
.B2(n_65),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_14),
.A2(n_62),
.B1(n_65),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_14),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_119),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_94),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_20),
.B(n_94),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_84),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_21),
.A2(n_22),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_23),
.B(n_41),
.C(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_34),
.B2(n_38),
.Y(n_23)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_24),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_26),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g82 ( 
.A1(n_26),
.A2(n_29),
.A3(n_32),
.B1(n_36),
.B2(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_26),
.B(n_37),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_28),
.B(n_30),
.Y(n_83)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_30),
.A2(n_45),
.A3(n_48),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_37),
.A2(n_60),
.B(n_65),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_37),
.A2(n_74),
.B1(n_76),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_40)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_43),
.A2(n_89),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_46),
.B(n_49),
.Y(n_133)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_47),
.A2(n_87),
.B(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_66),
.B2(n_68),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_55),
.A2(n_57),
.B1(n_68),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_57),
.A2(n_68),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_57),
.A2(n_68),
.B1(n_147),
.B2(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_61)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_61),
.A2(n_100),
.B1(n_127),
.B2(n_185),
.Y(n_184)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_62),
.B(n_170),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_66),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_71),
.B(n_84),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_81),
.B2(n_82),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_74),
.A2(n_76),
.B1(n_93),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_74),
.A2(n_76),
.B1(n_135),
.B2(n_156),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_74),
.A2(n_76),
.B1(n_161),
.B2(n_168),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_75),
.A2(n_103),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.C(n_92),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_85),
.B(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_92),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_107),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_118),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_139),
.B(n_195),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_136),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_122),
.B(n_136),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.C(n_128),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_123),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_130),
.A2(n_131),
.B1(n_134),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_189),
.B(n_194),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_177),
.B(n_188),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_157),
.B(n_176),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_150),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_153),
.C(n_155),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_165),
.B(n_175),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_163),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_171),
.B(n_174),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_179),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_184),
.C(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_190),
.B(n_191),
.Y(n_194)
);


endmodule