module fake_ariane_1985_n_721 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_721);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_721;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_443;
wire n_586;
wire n_286;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_202;
wire n_500;
wire n_665;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_672;
wire n_487;
wire n_422;
wire n_648;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_381;
wire n_344;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_365;
wire n_455;
wire n_429;
wire n_238;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_711;
wire n_453;
wire n_491;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_362;
wire n_543;
wire n_260;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_444;
wire n_355;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_292;
wire n_275;
wire n_704;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_434;
wire n_263;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g195 ( 
.A(n_91),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_100),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_148),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_84),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_99),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_104),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_115),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_179),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_81),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_153),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_42),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_66),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_54),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_150),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_94),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_53),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_129),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_76),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_40),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_114),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_156),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_88),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_126),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_102),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_79),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_33),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_151),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_50),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_138),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_103),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_131),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_139),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_31),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_137),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_49),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_97),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_35),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_72),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_14),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_22),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_165),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_38),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_172),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_162),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_159),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_73),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_178),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_59),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_55),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_8),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_167),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_3),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_69),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_98),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_85),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_17),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_16),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_86),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_71),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_117),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_152),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_82),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_89),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_161),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_189),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_80),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_4),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_185),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_170),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_155),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_105),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_63),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_93),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_101),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_21),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_9),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_30),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_45),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_27),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_144),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_74),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_34),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_119),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_140),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_128),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_70),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_15),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_191),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_90),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_19),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_26),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_136),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_186),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_64),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_183),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_48),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_18),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_29),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_175),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_10),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_65),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_132),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_187),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_21),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_57),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_135),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_7),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_0),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_147),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_116),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_96),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_10),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_11),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_24),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_180),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_23),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_123),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_61),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_13),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_58),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_92),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_171),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_145),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_12),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_169),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_15),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_87),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_111),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_56),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_313),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_249),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_217),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_249),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_227),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_237),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_273),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_285),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_257),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_228),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_318),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_236),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_314),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_251),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_292),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_255),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_239),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_202),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_267),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_269),
.B(n_0),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_274),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_275),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_287),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_207),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_290),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_291),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_304),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_246),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_240),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_275),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_240),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_248),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_248),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_252),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_308),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_256),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_312),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_316),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_219),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_319),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_324),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_326),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_196),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_284),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_219),
.B(n_1),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_284),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_276),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_242),
.B(n_2),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_195),
.B(n_2),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_197),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_199),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_198),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_200),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_201),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_203),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_213),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_204),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_214),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_224),
.B(n_4),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_205),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_206),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_225),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_233),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_208),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_244),
.B(n_5),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_209),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_210),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_247),
.B(n_6),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_298),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_253),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_258),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_259),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_261),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_262),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_298),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_266),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_211),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_212),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_270),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_280),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_245),
.B(n_6),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_283),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_215),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_289),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_295),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_216),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_301),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_302),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_303),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_305),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_218),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_306),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_309),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_220),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_221),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_317),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_381),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_373),
.B(n_321),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_352),
.B(n_320),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_334),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_357),
.B(n_245),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

AND2x6_ASAP7_75t_L g439 ( 
.A(n_358),
.B(n_250),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_330),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_327),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_333),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_342),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_331),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_345),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_428),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_386),
.A2(n_329),
.B(n_328),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_391),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_393),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_397),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_366),
.B(n_250),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_406),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_408),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g458 ( 
.A(n_336),
.B(n_328),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_343),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_363),
.B(n_222),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_346),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_226),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_365),
.B(n_272),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_424),
.B(n_229),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_425),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_367),
.B(n_230),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_377),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_410),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_348),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_351),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_368),
.B(n_231),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_403),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_SL g479 ( 
.A(n_336),
.B(n_272),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_340),
.B(n_232),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_379),
.A2(n_349),
.B(n_383),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_422),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_400),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_400),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_414),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_427),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_353),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_416),
.B(n_234),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_372),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_431),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_354),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_472),
.B(n_385),
.Y(n_494)
);

AND3x2_ASAP7_75t_L g495 ( 
.A(n_459),
.B(n_378),
.C(n_370),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_472),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_387),
.Y(n_497)
);

NAND2x1p5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_380),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_447),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_440),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_388),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_445),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_435),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_446),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_489),
.B(n_389),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_433),
.B(n_390),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_483),
.B(n_392),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_432),
.B(n_362),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_489),
.B(n_395),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_483),
.B(n_396),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_338),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_399),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_401),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_489),
.B(n_402),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_484),
.B(n_382),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_412),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_441),
.B(n_356),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_449),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_489),
.B(n_413),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_449),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_443),
.B(n_359),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_442),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_443),
.B(n_360),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_485),
.B(n_418),
.Y(n_525)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_449),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_467),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_444),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_467),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_467),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_463),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_434),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_454),
.B(n_272),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_463),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_486),
.B(n_436),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_450),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_453),
.Y(n_537)
);

AND2x6_ASAP7_75t_L g538 ( 
.A(n_478),
.B(n_350),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_464),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_455),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_456),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_491),
.B(n_361),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_457),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_468),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_470),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_539),
.B(n_474),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_471),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_518),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_546),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_532),
.B(n_486),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_532),
.A2(n_486),
.B1(n_458),
.B2(n_478),
.Y(n_552)
);

NAND3x1_ASAP7_75t_L g553 ( 
.A(n_508),
.B(n_477),
.C(n_480),
.Y(n_553)
);

AO22x2_ASAP7_75t_L g554 ( 
.A1(n_512),
.A2(n_524),
.B1(n_543),
.B2(n_522),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_501),
.B(n_488),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_516),
.B(n_335),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_523),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_537),
.Y(n_558)
);

OA22x2_ASAP7_75t_L g559 ( 
.A1(n_495),
.A2(n_341),
.B1(n_493),
.B2(n_481),
.Y(n_559)
);

AO22x2_ASAP7_75t_L g560 ( 
.A1(n_505),
.A2(n_337),
.B1(n_437),
.B2(n_344),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_541),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_528),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_496),
.A2(n_462),
.B1(n_479),
.B2(n_421),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_505),
.A2(n_437),
.B1(n_468),
.B2(n_355),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_507),
.B(n_492),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_542),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_544),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_511),
.B(n_371),
.Y(n_568)
);

AO22x2_ASAP7_75t_L g569 ( 
.A1(n_504),
.A2(n_355),
.B1(n_364),
.B2(n_490),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_531),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_494),
.B(n_451),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_534),
.Y(n_572)
);

AO22x2_ASAP7_75t_L g573 ( 
.A1(n_545),
.A2(n_502),
.B1(n_500),
.B2(n_510),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_509),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_513),
.B(n_466),
.Y(n_575)
);

AO22x2_ASAP7_75t_L g576 ( 
.A1(n_515),
.A2(n_364),
.B1(n_490),
.B2(n_374),
.Y(n_576)
);

AND2x6_ASAP7_75t_L g577 ( 
.A(n_513),
.B(n_452),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_514),
.B(n_517),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_497),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_540),
.Y(n_580)
);

AO22x2_ASAP7_75t_L g581 ( 
.A1(n_520),
.A2(n_369),
.B1(n_375),
.B2(n_374),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_521),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_521),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_498),
.B(n_460),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_525),
.A2(n_426),
.B1(n_430),
.B2(n_429),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_SL g586 ( 
.A(n_506),
.B(n_375),
.C(n_376),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_579),
.B(n_536),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_SL g589 ( 
.A(n_578),
.B(n_506),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_575),
.B(n_469),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_547),
.B(n_535),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_555),
.B(n_498),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_565),
.B(n_533),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_568),
.B(n_585),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_552),
.B(n_526),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_549),
.B(n_526),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_563),
.B(n_499),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_551),
.B(n_499),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_554),
.B(n_556),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_548),
.B(n_530),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_557),
.B(n_461),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_577),
.B(n_533),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_562),
.B(n_465),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_577),
.B(n_533),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_587),
.B(n_519),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_580),
.B(n_529),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_550),
.B(n_527),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_571),
.B(n_475),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_582),
.B(n_235),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_583),
.B(n_238),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_559),
.B(n_241),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_570),
.B(n_243),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_572),
.B(n_254),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_558),
.B(n_260),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_571),
.B(n_448),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_561),
.B(n_263),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_601),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_589),
.A2(n_584),
.B(n_573),
.Y(n_618)
);

AO31x2_ASAP7_75t_L g619 ( 
.A1(n_593),
.A2(n_574),
.A3(n_567),
.B(n_566),
.Y(n_619)
);

A2O1A1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_590),
.A2(n_586),
.B(n_573),
.C(n_553),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_608),
.B(n_439),
.Y(n_621)
);

NAND3x1_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_581),
.C(n_576),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_591),
.B(n_564),
.Y(n_623)
);

O2A1O1Ixp5_ASAP7_75t_L g624 ( 
.A1(n_594),
.A2(n_576),
.B(n_581),
.C(n_569),
.Y(n_624)
);

OA21x2_ASAP7_75t_L g625 ( 
.A1(n_592),
.A2(n_265),
.B(n_264),
.Y(n_625)
);

OA21x2_ASAP7_75t_L g626 ( 
.A1(n_597),
.A2(n_271),
.B(n_268),
.Y(n_626)
);

AO31x2_ASAP7_75t_L g627 ( 
.A1(n_602),
.A2(n_569),
.A3(n_560),
.B(n_439),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g628 ( 
.A1(n_598),
.A2(n_439),
.B(n_223),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_603),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_595),
.A2(n_606),
.B(n_605),
.Y(n_630)
);

OAI21x1_ASAP7_75t_L g631 ( 
.A1(n_604),
.A2(n_223),
.B(n_28),
.Y(n_631)
);

OAI22x1_ASAP7_75t_L g632 ( 
.A1(n_611),
.A2(n_278),
.B1(n_279),
.B2(n_277),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_607),
.A2(n_223),
.B(n_32),
.Y(n_633)
);

AO31x2_ASAP7_75t_L g634 ( 
.A1(n_615),
.A2(n_223),
.A3(n_36),
.B(n_37),
.Y(n_634)
);

OAI21xp33_ASAP7_75t_L g635 ( 
.A1(n_588),
.A2(n_596),
.B(n_609),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_610),
.A2(n_282),
.B(n_281),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_612),
.A2(n_288),
.B(n_286),
.Y(n_637)
);

AO21x2_ASAP7_75t_L g638 ( 
.A1(n_613),
.A2(n_41),
.B(n_39),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_600),
.A2(n_44),
.B(n_43),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_618),
.A2(n_616),
.B(n_614),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_628),
.A2(n_47),
.B(n_46),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_629),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_631),
.A2(n_52),
.B(n_51),
.Y(n_643)
);

AO21x2_ASAP7_75t_L g644 ( 
.A1(n_620),
.A2(n_294),
.B(n_293),
.Y(n_644)
);

AO21x2_ASAP7_75t_L g645 ( 
.A1(n_630),
.A2(n_299),
.B(n_296),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_617),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_633),
.A2(n_62),
.B(n_60),
.Y(n_647)
);

OAI21x1_ASAP7_75t_L g648 ( 
.A1(n_639),
.A2(n_68),
.B(n_67),
.Y(n_648)
);

AO31x2_ASAP7_75t_L g649 ( 
.A1(n_623),
.A2(n_141),
.A3(n_194),
.B(n_193),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_624),
.A2(n_325),
.B(n_323),
.C(n_322),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_621),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_626),
.A2(n_130),
.B(n_192),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_625),
.A2(n_127),
.B(n_190),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_619),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_635),
.B(n_20),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_636),
.A2(n_619),
.B(n_637),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_619),
.Y(n_657)
);

AO21x2_ASAP7_75t_L g658 ( 
.A1(n_638),
.A2(n_311),
.B(n_310),
.Y(n_658)
);

AO21x2_ASAP7_75t_L g659 ( 
.A1(n_634),
.A2(n_627),
.B(n_632),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_657),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_642),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_654),
.Y(n_662)
);

AO31x2_ASAP7_75t_L g663 ( 
.A1(n_640),
.A2(n_634),
.A3(n_627),
.B(n_622),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_646),
.Y(n_664)
);

OA21x2_ASAP7_75t_L g665 ( 
.A1(n_656),
.A2(n_118),
.B(n_188),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_643),
.A2(n_641),
.B(n_647),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_659),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_655),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_649),
.Y(n_669)
);

AO21x2_ASAP7_75t_L g670 ( 
.A1(n_645),
.A2(n_121),
.B(n_75),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_652),
.A2(n_122),
.B(n_77),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_644),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_648),
.A2(n_124),
.B(n_78),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_653),
.A2(n_125),
.B(n_83),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_651),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_661),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_R g677 ( 
.A(n_675),
.B(n_95),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_664),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_668),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_662),
.B(n_658),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_672),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_670),
.B(n_650),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_660),
.Y(n_683)
);

AND2x2_ASAP7_75t_SL g684 ( 
.A(n_665),
.B(n_669),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_663),
.B(n_106),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_660),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_683),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_676),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_686),
.Y(n_689)
);

INVx2_ASAP7_75t_R g690 ( 
.A(n_681),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_679),
.B(n_667),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_678),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_684),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_680),
.B(n_666),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_685),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_682),
.B(n_673),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_696),
.B(n_694),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_693),
.B(n_677),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_688),
.Y(n_699)
);

AO21x2_ASAP7_75t_L g700 ( 
.A1(n_695),
.A2(n_671),
.B(n_674),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_697),
.B(n_690),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_699),
.Y(n_702)
);

NAND2x1_ASAP7_75t_L g703 ( 
.A(n_701),
.B(n_697),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_702),
.B(n_698),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_704),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_705),
.B(n_703),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_706),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_707),
.Y(n_708)
);

NOR4xp25_ASAP7_75t_L g709 ( 
.A(n_708),
.B(n_692),
.C(n_687),
.D(n_689),
.Y(n_709)
);

AOI21x1_ASAP7_75t_L g710 ( 
.A1(n_709),
.A2(n_691),
.B(n_689),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_710),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_711),
.B(n_700),
.Y(n_712)
);

OAI32xp33_ASAP7_75t_L g713 ( 
.A1(n_712),
.A2(n_107),
.A3(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_713),
.A2(n_112),
.B(n_113),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_SL g715 ( 
.A1(n_714),
.A2(n_120),
.B1(n_133),
.B2(n_134),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_715),
.A2(n_142),
.B1(n_143),
.B2(n_146),
.Y(n_716)
);

XNOR2xp5_ASAP7_75t_L g717 ( 
.A(n_716),
.B(n_157),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_717),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_718),
.Y(n_719)
);

AOI221xp5_ASAP7_75t_L g720 ( 
.A1(n_719),
.A2(n_166),
.B1(n_173),
.B2(n_176),
.C(n_177),
.Y(n_720)
);

AOI211xp5_ASAP7_75t_L g721 ( 
.A1(n_720),
.A2(n_181),
.B(n_182),
.C(n_184),
.Y(n_721)
);


endmodule