module fake_ariane_457_n_1625 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1625);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1625;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_18),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_69),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_21),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_61),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_0),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_58),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_18),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_8),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_26),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_91),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_16),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_94),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_13),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_17),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_17),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_1),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_28),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_53),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_36),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_93),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_86),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_9),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_44),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_76),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_0),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_15),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_26),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_64),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_99),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_131),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_30),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_127),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_15),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_5),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_134),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_124),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_67),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_70),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_120),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_143),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_83),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_51),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_73),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_54),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_147),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_28),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_78),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_4),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_104),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_14),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_2),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_115),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_4),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_151),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_50),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_7),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_52),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_11),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_6),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_123),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_36),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_44),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_90),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_34),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_56),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_22),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_121),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_24),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_72),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_89),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_32),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_12),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_125),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_71),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_37),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_11),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_110),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_6),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_63),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_60),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_47),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_13),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_109),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_57),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_5),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_32),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_38),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_29),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_116),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_20),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_85),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_37),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_113),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_30),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_136),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_10),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_119),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_66),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_7),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_49),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_148),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_135),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_128),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_138),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_8),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_114),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_21),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_10),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_117),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_101),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_31),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_24),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_9),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_48),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_59),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_88),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_16),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_62),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_75),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_102),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_46),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_40),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_141),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_3),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_65),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_55),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_178),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_168),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_173),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_178),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_180),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_178),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_181),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_162),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_162),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_163),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_294),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_296),
.Y(n_317)
);

BUFx6f_ASAP7_75t_SL g318 ( 
.A(n_165),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_200),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_211),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_218),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_255),
.B(n_1),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_255),
.B(n_3),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_205),
.B(n_12),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_173),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_211),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_287),
.Y(n_330)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_205),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_221),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_223),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_223),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_291),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_154),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_165),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_154),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_165),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_183),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_221),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_206),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_209),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_183),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_160),
.B(n_14),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_187),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_187),
.B(n_19),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_220),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_189),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_221),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_189),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_190),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_221),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_190),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_294),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_225),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_201),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_201),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_216),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_216),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_165),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_233),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_232),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_233),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_157),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_238),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_256),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_274),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_238),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_248),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_167),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_294),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_177),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_179),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_301),
.B(n_169),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_317),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_302),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_305),
.B(n_169),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_316),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_307),
.B(n_280),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_373),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_373),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_337),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_339),
.Y(n_388)
);

AND2x6_ASAP7_75t_L g389 ( 
.A(n_325),
.B(n_176),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_331),
.B(n_249),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_374),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_345),
.B(n_280),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_346),
.A2(n_161),
.B(n_160),
.Y(n_396)
);

CKINVDCx11_ASAP7_75t_R g397 ( 
.A(n_303),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_309),
.B(n_161),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_331),
.B(n_166),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

BUFx8_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_333),
.B(n_166),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_310),
.B(n_248),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_371),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_334),
.B(n_175),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_311),
.B(n_251),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_312),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_313),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_315),
.B(n_294),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_320),
.B(n_175),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g420 ( 
.A(n_335),
.B(n_176),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_338),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_366),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_323),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_361),
.B(n_192),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_324),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

AND2x2_ASAP7_75t_SL g431 ( 
.A(n_328),
.B(n_195),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_336),
.B(n_251),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_326),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_304),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_340),
.B(n_174),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_318),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_327),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_329),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_362),
.B(n_192),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_321),
.B(n_254),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_372),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_403),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_403),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_377),
.B(n_321),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_427),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_403),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_389),
.A2(n_332),
.B1(n_354),
.B2(n_351),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_389),
.A2(n_332),
.B1(n_354),
.B2(n_351),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_254),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_431),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_421),
.B(n_314),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_422),
.B(n_273),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_417),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_389),
.A2(n_342),
.B1(n_298),
.B2(n_285),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_403),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_378),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_421),
.B(n_343),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_421),
.B(n_344),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_431),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_403),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_404),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_405),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_392),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_404),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_423),
.B(n_194),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_404),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_SL g479 ( 
.A(n_421),
.B(n_375),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_377),
.B(n_194),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_423),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_410),
.B(n_303),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_199),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_385),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_385),
.Y(n_486)
);

BUFx6f_ASAP7_75t_SL g487 ( 
.A(n_431),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_439),
.B(n_349),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_381),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_389),
.A2(n_342),
.B1(n_298),
.B2(n_285),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_427),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_389),
.A2(n_273),
.B1(n_294),
.B2(n_197),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_440),
.B(n_199),
.Y(n_494)
);

AND3x2_ASAP7_75t_L g495 ( 
.A(n_391),
.B(n_282),
.C(n_208),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_394),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_439),
.B(n_357),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_L g498 ( 
.A(n_421),
.B(n_212),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_415),
.B(n_186),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_389),
.A2(n_174),
.B1(n_207),
.B2(n_235),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_423),
.B(n_212),
.Y(n_502)
);

NOR3xp33_ASAP7_75t_L g503 ( 
.A(n_399),
.B(n_222),
.C(n_191),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_404),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_381),
.Y(n_506)
);

BUFx10_ASAP7_75t_L g507 ( 
.A(n_421),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_415),
.B(n_224),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_408),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_421),
.B(n_226),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_415),
.B(n_228),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_408),
.Y(n_512)
);

AND3x2_ASAP7_75t_L g513 ( 
.A(n_391),
.B(n_410),
.C(n_434),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_389),
.A2(n_207),
.B1(n_235),
.B2(n_203),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_381),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_381),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_400),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_439),
.A2(n_258),
.B1(n_231),
.B2(n_234),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_405),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_440),
.B(n_214),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_425),
.B(n_430),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_442),
.B(n_443),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_442),
.B(n_214),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_408),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_436),
.B(n_219),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_408),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_436),
.B(n_219),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_436),
.B(n_237),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_442),
.B(n_237),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_408),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_443),
.B(n_239),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_441),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_441),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_381),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_381),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_383),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_383),
.Y(n_537)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_425),
.B(n_243),
.C(n_240),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_389),
.A2(n_195),
.B1(n_203),
.B2(n_210),
.Y(n_539)
);

BUFx4f_ASAP7_75t_L g540 ( 
.A(n_396),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_415),
.B(n_239),
.Y(n_541)
);

OAI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_428),
.A2(n_236),
.B1(n_230),
.B2(n_267),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_389),
.A2(n_210),
.B1(n_261),
.B2(n_244),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_396),
.A2(n_278),
.B1(n_265),
.B2(n_281),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_408),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_383),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_415),
.B(n_252),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_416),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_383),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_416),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_415),
.B(n_259),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_383),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_405),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_425),
.B(n_252),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_395),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_441),
.A2(n_269),
.B1(n_260),
.B2(n_263),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_415),
.B(n_155),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_395),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_416),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_397),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_396),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_383),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_435),
.B(n_253),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_416),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_424),
.B(n_253),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_383),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_379),
.B(n_306),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_416),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_400),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_379),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_425),
.B(n_264),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_424),
.B(n_264),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_401),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_425),
.A2(n_286),
.B1(n_279),
.B2(n_270),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_426),
.B(n_270),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_386),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_SL g578 ( 
.A(n_425),
.B(n_279),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_426),
.B(n_364),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_386),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_401),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_402),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_416),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_430),
.B(n_153),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_434),
.B(n_306),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_430),
.B(n_156),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_556),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_556),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_507),
.B(n_430),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_471),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_522),
.B(n_430),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_456),
.B(n_430),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_492),
.B(n_429),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_446),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_492),
.B(n_429),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_559),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_463),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_507),
.B(n_428),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_463),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_454),
.B(n_409),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_469),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_531),
.A2(n_413),
.B1(n_406),
.B2(n_420),
.Y(n_602)
);

BUFx6f_ASAP7_75t_SL g603 ( 
.A(n_454),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_466),
.B(n_433),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_532),
.B(n_433),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_469),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_561),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_507),
.B(n_416),
.Y(n_608)
);

NOR2x1p5_ASAP7_75t_L g609 ( 
.A(n_561),
.B(n_554),
.Y(n_609)
);

AND2x2_ASAP7_75t_SL g610 ( 
.A(n_461),
.B(n_396),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_523),
.B(n_420),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_571),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_447),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_491),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_532),
.B(n_438),
.Y(n_615)
);

AO22x2_ASAP7_75t_L g616 ( 
.A1(n_466),
.A2(n_437),
.B1(n_432),
.B2(n_438),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_529),
.B(n_449),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_554),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_449),
.B(n_420),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_496),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_568),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_449),
.B(n_420),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_579),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_564),
.A2(n_420),
.B1(n_411),
.B2(n_402),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_488),
.B(n_437),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_448),
.B(n_437),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_497),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_420),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_533),
.B(n_411),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_573),
.B(n_420),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_533),
.B(n_412),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_549),
.B(n_540),
.Y(n_632)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_503),
.B(n_412),
.C(n_432),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_513),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_517),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_575),
.A2(n_420),
.B1(n_396),
.B2(n_388),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_518),
.B(n_432),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_494),
.B(n_420),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_490),
.A2(n_407),
.B1(n_390),
.B2(n_387),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_557),
.B(n_387),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_455),
.B(n_382),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_520),
.B(n_499),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_570),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_499),
.B(n_387),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_476),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_508),
.B(n_388),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_511),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_511),
.B(n_390),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_552),
.B(n_390),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_495),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_485),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_574),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_458),
.B(n_398),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_552),
.B(n_407),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_549),
.B(n_540),
.Y(n_655)
);

NOR2x1p5_ASAP7_75t_L g656 ( 
.A(n_470),
.B(n_398),
.Y(n_656)
);

NOR3xp33_ASAP7_75t_L g657 ( 
.A(n_542),
.B(n_407),
.C(n_419),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_464),
.B(n_419),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_465),
.B(n_409),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_549),
.B(n_409),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_581),
.B(n_418),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_585),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_455),
.B(n_382),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_418),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_457),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_460),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_585),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_486),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_479),
.B(n_393),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_540),
.A2(n_418),
.B(n_414),
.C(n_393),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_445),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_558),
.B(n_418),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_483),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_539),
.A2(n_544),
.B1(n_514),
.B2(n_543),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_558),
.B(n_418),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_479),
.B(n_393),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_558),
.B(n_382),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_459),
.B(n_414),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_482),
.B(n_393),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_576),
.B(n_376),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_459),
.B(n_451),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_482),
.B(n_414),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_541),
.B(n_376),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_547),
.B(n_376),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_480),
.B(n_376),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_525),
.B(n_376),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_444),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_445),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_444),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_452),
.B(n_364),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_521),
.A2(n_386),
.B(n_384),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_447),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_SL g693 ( 
.A1(n_568),
.A2(n_330),
.B1(n_319),
.B2(n_322),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_445),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_525),
.B(n_384),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_453),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_525),
.B(n_384),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_447),
.B(n_158),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_453),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_447),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_447),
.B(n_159),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_470),
.B(n_384),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_578),
.A2(n_384),
.B1(n_185),
.B2(n_242),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_525),
.B(n_164),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_487),
.B(n_19),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_578),
.A2(n_188),
.B1(n_193),
.B2(n_184),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_450),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_525),
.B(n_170),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_450),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_462),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_462),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_477),
.B(n_368),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_487),
.B(n_20),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_467),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_525),
.B(n_171),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_527),
.B(n_172),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_487),
.B(n_22),
.Y(n_717)
);

AND2x6_ASAP7_75t_SL g718 ( 
.A(n_483),
.B(n_308),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_467),
.Y(n_719)
);

OAI21xp5_ASAP7_75t_L g720 ( 
.A1(n_572),
.A2(n_202),
.B(n_300),
.Y(n_720)
);

AO221x1_ASAP7_75t_L g721 ( 
.A1(n_481),
.A2(n_369),
.B1(n_368),
.B2(n_330),
.C(n_322),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_468),
.Y(n_722)
);

INVx8_ASAP7_75t_L g723 ( 
.A(n_527),
.Y(n_723)
);

INVx8_ASAP7_75t_L g724 ( 
.A(n_527),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_527),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_562),
.B(n_23),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_562),
.B(n_510),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_481),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_527),
.B(n_182),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_481),
.B(n_23),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_527),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_468),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_504),
.B(n_25),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_528),
.B(n_196),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_478),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_477),
.B(n_308),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_L g737 ( 
.A(n_493),
.B(n_257),
.C(n_299),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_478),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_472),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_519),
.B(n_198),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_500),
.A2(n_155),
.B1(n_386),
.B2(n_319),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_519),
.B(n_262),
.Y(n_742)
);

OAI21xp5_ASAP7_75t_L g743 ( 
.A1(n_632),
.A2(n_526),
.B(n_545),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_627),
.B(n_528),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_591),
.A2(n_584),
.B(n_586),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_613),
.Y(n_746)
);

AOI21xp33_ASAP7_75t_L g747 ( 
.A1(n_623),
.A2(n_498),
.B(n_538),
.Y(n_747)
);

AOI21x1_ASAP7_75t_L g748 ( 
.A1(n_632),
.A2(n_512),
.B(n_526),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_587),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_613),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_612),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_627),
.B(n_604),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_623),
.B(n_528),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_591),
.A2(n_655),
.B(n_589),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_602),
.A2(n_504),
.B1(n_530),
.B2(n_509),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_660),
.A2(n_498),
.B(n_501),
.C(n_545),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_604),
.B(n_528),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_594),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_588),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_634),
.B(n_528),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_655),
.A2(n_512),
.B(n_505),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_626),
.B(n_528),
.Y(n_762)
);

AO21x1_ASAP7_75t_L g763 ( 
.A1(n_726),
.A2(n_501),
.B(n_505),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_589),
.A2(n_509),
.B(n_524),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_598),
.A2(n_524),
.B(n_530),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_626),
.B(n_474),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_629),
.B(n_474),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_590),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_629),
.B(n_474),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_670),
.A2(n_524),
.B(n_530),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_723),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_647),
.A2(n_555),
.B1(n_474),
.B2(n_484),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_598),
.A2(n_608),
.B(n_592),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_647),
.A2(n_555),
.B1(n_474),
.B2(n_484),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_631),
.B(n_474),
.Y(n_775)
);

OAI21xp5_ASAP7_75t_L g776 ( 
.A1(n_726),
.A2(n_555),
.B(n_551),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_R g777 ( 
.A(n_618),
.B(n_607),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_660),
.A2(n_560),
.B(n_551),
.C(n_548),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_631),
.B(n_484),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_678),
.B(n_484),
.Y(n_780)
);

CKINVDCx10_ASAP7_75t_R g781 ( 
.A(n_712),
.Y(n_781)
);

OAI21xp33_ASAP7_75t_L g782 ( 
.A1(n_605),
.A2(n_548),
.B(n_551),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_608),
.A2(n_548),
.B(n_560),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_702),
.B(n_641),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_642),
.B(n_484),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_592),
.A2(n_560),
.B(n_580),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_621),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_633),
.B(n_653),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_663),
.B(n_484),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_615),
.B(n_502),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_682),
.A2(n_537),
.B(n_580),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_653),
.A2(n_565),
.B(n_569),
.C(n_577),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_613),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_658),
.B(n_502),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_679),
.A2(n_536),
.B(n_577),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_699),
.A2(n_536),
.B(n_489),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_600),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_650),
.B(n_565),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_638),
.A2(n_555),
.B(n_489),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_658),
.B(n_502),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_596),
.A2(n_535),
.B(n_506),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_617),
.B(n_502),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_636),
.A2(n_555),
.B(n_506),
.Y(n_803)
);

OR2x2_ASAP7_75t_SL g804 ( 
.A(n_693),
.B(n_515),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_633),
.B(n_472),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_705),
.B(n_472),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_705),
.B(n_472),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_673),
.B(n_516),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_687),
.A2(n_546),
.B(n_534),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_628),
.A2(n_555),
.B(n_534),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_659),
.B(n_680),
.Y(n_811)
);

OAI321xp33_ASAP7_75t_L g812 ( 
.A1(n_674),
.A2(n_386),
.A3(n_567),
.B1(n_563),
.B2(n_553),
.C(n_546),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_689),
.A2(n_567),
.B(n_563),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_736),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_713),
.B(n_475),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_630),
.A2(n_553),
.B(n_535),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_707),
.A2(n_516),
.B(n_475),
.Y(n_817)
);

NAND2x1_ASAP7_75t_L g818 ( 
.A(n_671),
.B(n_475),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_713),
.B(n_475),
.Y(n_819)
);

BUFx4f_ASAP7_75t_L g820 ( 
.A(n_600),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_662),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_614),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_659),
.B(n_502),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_681),
.B(n_502),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_593),
.B(n_475),
.Y(n_825)
);

AO21x1_ASAP7_75t_L g826 ( 
.A1(n_727),
.A2(n_611),
.B(n_644),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_709),
.A2(n_583),
.B(n_550),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_662),
.B(n_583),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_595),
.B(n_583),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_610),
.B(n_583),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_710),
.A2(n_583),
.B(n_550),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_620),
.B(n_550),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_635),
.B(n_550),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_643),
.B(n_550),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_613),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_610),
.A2(n_473),
.B1(n_266),
.B2(n_297),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_652),
.B(n_473),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_665),
.B(n_473),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_666),
.B(n_473),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_616),
.B(n_473),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_677),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_674),
.A2(n_247),
.B1(n_293),
.B2(n_292),
.Y(n_842)
);

CKINVDCx10_ASAP7_75t_R g843 ( 
.A(n_712),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_711),
.A2(n_246),
.B(n_289),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_616),
.B(n_245),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_714),
.A2(n_722),
.B(n_719),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_717),
.A2(n_241),
.B1(n_288),
.B2(n_283),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_616),
.B(n_229),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_732),
.A2(n_227),
.B(n_277),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_691),
.A2(n_386),
.B(n_276),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_692),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_637),
.B(n_217),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_735),
.A2(n_215),
.B(n_275),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_738),
.A2(n_213),
.B(n_271),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_685),
.B(n_625),
.Y(n_855)
);

O2A1O1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_661),
.A2(n_25),
.B(n_27),
.C(n_31),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_597),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_717),
.B(n_204),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_664),
.A2(n_27),
.B(n_35),
.C(n_38),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_692),
.B(n_268),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_712),
.B(n_667),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_692),
.B(n_250),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_646),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_692),
.Y(n_864)
);

NAND3xp33_ASAP7_75t_L g865 ( 
.A(n_657),
.B(n_39),
.C(n_41),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_700),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_648),
.B(n_649),
.Y(n_867)
);

AOI33xp33_ASAP7_75t_L g868 ( 
.A1(n_624),
.A2(n_41),
.A3(n_42),
.B1(n_43),
.B2(n_45),
.B3(n_46),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_654),
.B(n_42),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_599),
.Y(n_870)
);

OAI21x1_ASAP7_75t_L g871 ( 
.A1(n_694),
.A2(n_96),
.B(n_140),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_657),
.B(n_43),
.Y(n_872)
);

AND2x6_ASAP7_75t_L g873 ( 
.A(n_727),
.B(n_95),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_730),
.A2(n_45),
.B(n_47),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_600),
.A2(n_48),
.B1(n_49),
.B2(n_77),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_694),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_730),
.A2(n_84),
.B(n_92),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_601),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_728),
.A2(n_97),
.B(n_103),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_667),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_683),
.B(n_105),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_728),
.A2(n_107),
.B(n_111),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_698),
.A2(n_126),
.B(n_132),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_609),
.B(n_150),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_700),
.B(n_133),
.Y(n_885)
);

NOR2x1_ASAP7_75t_L g886 ( 
.A(n_656),
.B(n_139),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_684),
.B(n_600),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_733),
.A2(n_720),
.B(n_640),
.C(n_606),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_700),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_645),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_698),
.A2(n_701),
.B(n_739),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_603),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_700),
.B(n_739),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_672),
.B(n_675),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_651),
.Y(n_895)
);

NOR2x1p5_ASAP7_75t_SL g896 ( 
.A(n_668),
.B(n_739),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_701),
.A2(n_739),
.B(n_622),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_723),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_686),
.B(n_697),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_619),
.A2(n_715),
.B(n_729),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_600),
.B(n_725),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_639),
.A2(n_695),
.B(n_737),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_706),
.B(n_703),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_741),
.B(n_669),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_704),
.A2(n_708),
.B(n_716),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_676),
.A2(n_742),
.B(n_740),
.C(n_734),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_721),
.B(n_741),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_SL g908 ( 
.A(n_723),
.B(n_724),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_603),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_731),
.A2(n_724),
.B(n_718),
.Y(n_910)
);

AO21x1_ASAP7_75t_L g911 ( 
.A1(n_591),
.A2(n_726),
.B(n_727),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_627),
.B(n_604),
.Y(n_912)
);

OAI21xp33_ASAP7_75t_L g913 ( 
.A1(n_627),
.A2(n_399),
.B(n_391),
.Y(n_913)
);

NOR2x1p5_ASAP7_75t_SL g914 ( 
.A(n_688),
.B(n_696),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_913),
.A2(n_788),
.B(n_752),
.C(n_912),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_SL g916 ( 
.A(n_797),
.B(n_820),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_822),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_797),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_771),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_SL g920 ( 
.A(n_820),
.B(n_908),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_771),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_811),
.A2(n_874),
.B1(n_872),
.B2(n_767),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_867),
.B(n_841),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_751),
.B(n_784),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_771),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_746),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_857),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_769),
.A2(n_779),
.B(n_775),
.Y(n_928)
);

AOI21x1_ASAP7_75t_L g929 ( 
.A1(n_850),
.A2(n_754),
.B(n_748),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_894),
.B(n_855),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_784),
.B(n_768),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_766),
.A2(n_745),
.B(n_794),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_814),
.B(n_861),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_777),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_771),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_880),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_787),
.B(n_808),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_800),
.A2(n_773),
.B(n_881),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_903),
.A2(n_823),
.B(n_877),
.C(n_757),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_888),
.A2(n_776),
.B(n_762),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_749),
.B(n_759),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_877),
.A2(n_785),
.B(n_906),
.C(n_865),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_870),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_780),
.A2(n_789),
.B1(n_875),
.B2(n_790),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_828),
.B(n_821),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_907),
.A2(n_842),
.B1(n_760),
.B2(n_904),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_899),
.B(n_824),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_755),
.A2(n_792),
.B(n_770),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_887),
.B(n_753),
.Y(n_949)
);

BUFx8_ASAP7_75t_SL g950 ( 
.A(n_884),
.Y(n_950)
);

CKINVDCx16_ASAP7_75t_R g951 ( 
.A(n_909),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_892),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_746),
.Y(n_953)
);

XOR2xp5_ASAP7_75t_L g954 ( 
.A(n_910),
.B(n_847),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_R g955 ( 
.A(n_781),
.B(n_843),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_816),
.A2(n_900),
.B(n_803),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_763),
.A2(n_911),
.B(n_905),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_878),
.B(n_890),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_858),
.B(n_798),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_895),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_869),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_804),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_801),
.A2(n_829),
.B(n_825),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_817),
.A2(n_809),
.B(n_813),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_901),
.B(n_744),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_746),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_805),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_868),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_901),
.B(n_772),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_774),
.B(n_908),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_842),
.B(n_873),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_786),
.A2(n_846),
.B(n_765),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_802),
.A2(n_747),
.B(n_902),
.C(n_778),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_840),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_836),
.A2(n_782),
.B1(n_756),
.B2(n_852),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_896),
.B(n_898),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_836),
.A2(n_845),
.B1(n_848),
.B2(n_873),
.Y(n_977)
);

AOI22xp5_ASAP7_75t_L g978 ( 
.A1(n_830),
.A2(n_873),
.B1(n_806),
.B2(n_807),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_793),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_830),
.B(n_873),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_891),
.A2(n_764),
.B(n_795),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_863),
.A2(n_770),
.B1(n_755),
.B2(n_838),
.Y(n_982)
);

BUFx4f_ASAP7_75t_L g983 ( 
.A(n_793),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_SL g984 ( 
.A(n_856),
.B(n_859),
.C(n_862),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_815),
.A2(n_819),
.B1(n_886),
.B2(n_826),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_832),
.A2(n_837),
.B1(n_834),
.B2(n_833),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_750),
.B(n_851),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_816),
.A2(n_803),
.B(n_897),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_839),
.Y(n_989)
);

BUFx5_ASAP7_75t_L g990 ( 
.A(n_793),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_866),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_866),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_750),
.B(n_835),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_835),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_851),
.B(n_864),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_898),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_864),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_791),
.A2(n_827),
.B(n_831),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_914),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_889),
.B(n_860),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_876),
.B(n_853),
.C(n_854),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_844),
.Y(n_1002)
);

O2A1O1Ixp5_ASAP7_75t_L g1003 ( 
.A1(n_893),
.A2(n_818),
.B(n_761),
.C(n_743),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_849),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_885),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_743),
.B(n_761),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_783),
.B(n_810),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_810),
.A2(n_799),
.B1(n_883),
.B2(n_796),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_SL g1009 ( 
.A1(n_799),
.A2(n_812),
.B1(n_871),
.B2(n_879),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_812),
.A2(n_591),
.B(n_767),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_882),
.B(n_784),
.Y(n_1011)
);

OR2x6_ASAP7_75t_L g1012 ( 
.A(n_797),
.B(n_712),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_752),
.B(n_912),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_746),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_SL g1015 ( 
.A1(n_752),
.A2(n_912),
.B(n_655),
.C(n_632),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_822),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_746),
.Y(n_1017)
);

AO21x2_ASAP7_75t_L g1018 ( 
.A1(n_763),
.A2(n_911),
.B(n_812),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_752),
.B(n_912),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_913),
.A2(n_627),
.B(n_623),
.C(n_788),
.Y(n_1020)
);

CKINVDCx8_ASAP7_75t_R g1021 ( 
.A(n_781),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_752),
.A2(n_912),
.B1(n_627),
.B2(n_602),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_752),
.B(n_912),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_913),
.A2(n_627),
.B(n_788),
.C(n_752),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_752),
.B(n_627),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_797),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_752),
.B(n_912),
.Y(n_1027)
);

INVx3_ASAP7_75t_SL g1028 ( 
.A(n_821),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_SL g1029 ( 
.A(n_797),
.B(n_820),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_752),
.B(n_912),
.Y(n_1030)
);

OAI21xp33_ASAP7_75t_SL g1031 ( 
.A1(n_788),
.A2(n_877),
.B(n_752),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_777),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_797),
.Y(n_1033)
);

BUFx2_ASAP7_75t_SL g1034 ( 
.A(n_751),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_752),
.B(n_912),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_752),
.B(n_912),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_752),
.A2(n_912),
.B1(n_627),
.B2(n_602),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_752),
.B(n_912),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_913),
.A2(n_627),
.B(n_623),
.C(n_788),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_913),
.A2(n_627),
.B(n_623),
.C(n_788),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_752),
.B(n_912),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_752),
.B(n_912),
.Y(n_1042)
);

OR2x6_ASAP7_75t_SL g1043 ( 
.A(n_842),
.B(n_561),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_758),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_1025),
.B(n_1019),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1022),
.A2(n_1037),
.B1(n_1030),
.B2(n_1019),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_972),
.A2(n_981),
.B(n_998),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_1010),
.A2(n_922),
.B(n_940),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_917),
.Y(n_1049)
);

AOI221xp5_ASAP7_75t_L g1050 ( 
.A1(n_922),
.A2(n_1022),
.B1(n_1037),
.B2(n_915),
.C(n_1030),
.Y(n_1050)
);

NAND2x1_ASAP7_75t_L g1051 ( 
.A(n_918),
.B(n_1026),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1038),
.B(n_1042),
.Y(n_1052)
);

CKINVDCx11_ASAP7_75t_R g1053 ( 
.A(n_1021),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_936),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_1020),
.A2(n_1040),
.B(n_1039),
.C(n_1024),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_1013),
.B(n_1023),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_933),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_1032),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1016),
.Y(n_1059)
);

INVx3_ASAP7_75t_SL g1060 ( 
.A(n_1028),
.Y(n_1060)
);

AND2x2_ASAP7_75t_SL g1061 ( 
.A(n_971),
.B(n_946),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_923),
.A2(n_968),
.B1(n_1041),
.B2(n_1036),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_1034),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_942),
.A2(n_961),
.B(n_977),
.C(n_984),
.Y(n_1064)
);

BUFx8_ASAP7_75t_SL g1065 ( 
.A(n_934),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_973),
.A2(n_928),
.B(n_982),
.Y(n_1066)
);

AOI221xp5_ASAP7_75t_SL g1067 ( 
.A1(n_982),
.A2(n_1027),
.B1(n_1035),
.B2(n_948),
.C(n_975),
.Y(n_1067)
);

NOR2xp67_ASAP7_75t_SL g1068 ( 
.A(n_951),
.B(n_918),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_937),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_919),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_952),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_986),
.A2(n_1009),
.B(n_1007),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_1008),
.A2(n_975),
.A3(n_986),
.B(n_999),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_964),
.A2(n_929),
.B(n_963),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_948),
.A2(n_932),
.B(n_957),
.C(n_1008),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_919),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_931),
.Y(n_1077)
);

NAND3xp33_ASAP7_75t_SL g1078 ( 
.A(n_1004),
.B(n_955),
.C(n_945),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_930),
.A2(n_1002),
.B(n_1001),
.C(n_959),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_980),
.A2(n_944),
.A3(n_989),
.B(n_949),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_988),
.A2(n_956),
.B(n_1003),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1015),
.A2(n_970),
.B(n_1011),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_924),
.B(n_941),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_SL g1084 ( 
.A1(n_987),
.A2(n_993),
.B(n_969),
.C(n_941),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_943),
.Y(n_1085)
);

AOI31xp67_ASAP7_75t_L g1086 ( 
.A1(n_985),
.A2(n_978),
.A3(n_1006),
.B(n_965),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_947),
.B(n_962),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1043),
.B(n_1012),
.Y(n_1088)
);

AO32x2_ASAP7_75t_L g1089 ( 
.A1(n_1005),
.A2(n_1018),
.A3(n_974),
.B1(n_921),
.B2(n_935),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_920),
.A2(n_916),
.B(n_1029),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_920),
.A2(n_916),
.B(n_1029),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_966),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_926),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_925),
.A2(n_1033),
.B(n_1026),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1018),
.A2(n_1005),
.B(n_1033),
.Y(n_1095)
);

AO21x1_ASAP7_75t_L g1096 ( 
.A1(n_1000),
.A2(n_954),
.B(n_995),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_967),
.B(n_1012),
.Y(n_1097)
);

CKINVDCx12_ASAP7_75t_R g1098 ( 
.A(n_976),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_925),
.A2(n_996),
.B(n_994),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_950),
.B(n_997),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_927),
.B(n_1044),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_996),
.A2(n_976),
.B(n_958),
.C(n_979),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_960),
.A2(n_921),
.A3(n_935),
.B(n_976),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_990),
.A2(n_926),
.B(n_953),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_926),
.A2(n_953),
.B(n_991),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_953),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_990),
.A2(n_991),
.A3(n_992),
.B(n_1014),
.Y(n_1107)
);

AOI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1017),
.A2(n_913),
.B1(n_391),
.B2(n_1025),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_990),
.A2(n_1014),
.B(n_1017),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_990),
.A2(n_972),
.B(n_981),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1017),
.A2(n_591),
.B(n_939),
.Y(n_1111)
);

BUFx4f_ASAP7_75t_SL g1112 ( 
.A(n_1032),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1031),
.A2(n_627),
.B(n_623),
.C(n_913),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_983),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1025),
.B(n_933),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1031),
.A2(n_913),
.B(n_627),
.C(n_915),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_939),
.A2(n_591),
.B(n_938),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_939),
.A2(n_591),
.B(n_938),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_939),
.A2(n_591),
.B(n_938),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1032),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1025),
.B(n_933),
.Y(n_1121)
);

INVx3_ASAP7_75t_SL g1122 ( 
.A(n_1028),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_939),
.A2(n_591),
.B(n_938),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1019),
.B(n_1030),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_983),
.Y(n_1125)
);

BUFx2_ASAP7_75t_R g1126 ( 
.A(n_1021),
.Y(n_1126)
);

BUFx12f_ASAP7_75t_L g1127 ( 
.A(n_934),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1008),
.A2(n_763),
.A3(n_911),
.B(n_826),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1032),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1025),
.B(n_1038),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_1008),
.A2(n_763),
.A3(n_911),
.B(n_826),
.Y(n_1131)
);

OR2x6_ASAP7_75t_L g1132 ( 
.A(n_1012),
.B(n_797),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_1034),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_917),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_972),
.A2(n_981),
.B(n_998),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1025),
.B(n_933),
.Y(n_1136)
);

OR2x6_ASAP7_75t_L g1137 ( 
.A(n_1012),
.B(n_797),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_936),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_972),
.A2(n_981),
.B(n_998),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_939),
.A2(n_591),
.B(n_938),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1025),
.A2(n_913),
.B1(n_391),
.B2(n_627),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_1008),
.A2(n_763),
.A3(n_911),
.B(n_826),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_972),
.A2(n_981),
.B(n_998),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1031),
.A2(n_913),
.B(n_627),
.C(n_915),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1019),
.B(n_1030),
.Y(n_1145)
);

CKINVDCx6p67_ASAP7_75t_R g1146 ( 
.A(n_1028),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_1019),
.B(n_1030),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_1008),
.A2(n_763),
.A3(n_911),
.B(n_826),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_936),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_939),
.A2(n_591),
.B(n_938),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_983),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1031),
.A2(n_939),
.B(n_922),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1019),
.B(n_1030),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1025),
.B(n_933),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_939),
.A2(n_591),
.B(n_938),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_917),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1025),
.B(n_627),
.Y(n_1157)
);

CKINVDCx11_ASAP7_75t_R g1158 ( 
.A(n_1021),
.Y(n_1158)
);

NOR2xp67_ASAP7_75t_L g1159 ( 
.A(n_925),
.B(n_919),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1025),
.B(n_933),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_917),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_983),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1031),
.A2(n_939),
.B(n_922),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_939),
.A2(n_591),
.B(n_938),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1008),
.A2(n_763),
.A3(n_911),
.B(n_826),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_936),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1045),
.A2(n_1157),
.B1(n_1141),
.B2(n_1130),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1049),
.Y(n_1168)
);

INVx1_ASAP7_75t_SL g1169 ( 
.A(n_1063),
.Y(n_1169)
);

BUFx10_ASAP7_75t_L g1170 ( 
.A(n_1100),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1062),
.A2(n_1108),
.B1(n_1046),
.B2(n_1145),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1065),
.Y(n_1172)
);

CKINVDCx6p67_ASAP7_75t_R g1173 ( 
.A(n_1053),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_1158),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1061),
.A2(n_1062),
.B1(n_1096),
.B2(n_1046),
.Y(n_1175)
);

BUFx4f_ASAP7_75t_SL g1176 ( 
.A(n_1127),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1126),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1152),
.A2(n_1163),
.B1(n_1088),
.B2(n_1087),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1112),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_SL g1180 ( 
.A1(n_1152),
.A2(n_1163),
.B1(n_1066),
.B2(n_1124),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1050),
.A2(n_1147),
.B1(n_1124),
.B2(n_1108),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1066),
.A2(n_1154),
.B1(n_1136),
.B2(n_1115),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1059),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1058),
.Y(n_1184)
);

INVx6_ASAP7_75t_L g1185 ( 
.A(n_1125),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_SL g1186 ( 
.A1(n_1121),
.A2(n_1160),
.B1(n_1083),
.B2(n_1052),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_1151),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_1146),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_1060),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1120),
.Y(n_1190)
);

INVx6_ASAP7_75t_L g1191 ( 
.A(n_1151),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1057),
.A2(n_1056),
.B1(n_1069),
.B2(n_1072),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1153),
.A2(n_1078),
.B1(n_1085),
.B2(n_1134),
.Y(n_1193)
);

OAI22x1_ASAP7_75t_SL g1194 ( 
.A1(n_1063),
.A2(n_1133),
.B1(n_1092),
.B2(n_1122),
.Y(n_1194)
);

CKINVDCx11_ASAP7_75t_R g1195 ( 
.A(n_1071),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1077),
.A2(n_1101),
.B1(n_1161),
.B2(n_1156),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1068),
.A2(n_1067),
.B1(n_1064),
.B2(n_1133),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1138),
.B(n_1149),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1097),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1129),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1048),
.A2(n_1137),
.B1(n_1132),
.B2(n_1166),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1106),
.Y(n_1202)
);

CKINVDCx14_ASAP7_75t_R g1203 ( 
.A(n_1054),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1162),
.Y(n_1204)
);

OAI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1090),
.A2(n_1091),
.B1(n_1082),
.B2(n_1140),
.Y(n_1205)
);

INVxp67_ASAP7_75t_SL g1206 ( 
.A(n_1081),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1116),
.A2(n_1144),
.B1(n_1055),
.B2(n_1113),
.Y(n_1207)
);

BUFx8_ASAP7_75t_SL g1208 ( 
.A(n_1070),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1117),
.A2(n_1164),
.B1(n_1155),
.B2(n_1118),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1095),
.A2(n_1111),
.B1(n_1093),
.B2(n_1119),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1079),
.A2(n_1123),
.B1(n_1150),
.B2(n_1051),
.Y(n_1211)
);

BUFx10_ASAP7_75t_L g1212 ( 
.A(n_1093),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1109),
.A2(n_1081),
.B1(n_1099),
.B2(n_1070),
.Y(n_1213)
);

INVx6_ASAP7_75t_L g1214 ( 
.A(n_1098),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_SL g1215 ( 
.A1(n_1086),
.A2(n_1073),
.B1(n_1080),
.B2(n_1084),
.Y(n_1215)
);

NAND2x1p5_ASAP7_75t_L g1216 ( 
.A(n_1076),
.B(n_1159),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1109),
.A2(n_1073),
.B1(n_1159),
.B2(n_1105),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_SL g1218 ( 
.A(n_1073),
.B(n_1075),
.Y(n_1218)
);

INVx4_ASAP7_75t_L g1219 ( 
.A(n_1107),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1107),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_1047),
.Y(n_1221)
);

BUFx12f_ASAP7_75t_L g1222 ( 
.A(n_1107),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1102),
.A2(n_1128),
.B(n_1148),
.Y(n_1223)
);

BUFx8_ASAP7_75t_L g1224 ( 
.A(n_1089),
.Y(n_1224)
);

CKINVDCx11_ASAP7_75t_R g1225 ( 
.A(n_1089),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1094),
.A2(n_1104),
.B1(n_1074),
.B2(n_1110),
.Y(n_1226)
);

CKINVDCx6p67_ASAP7_75t_R g1227 ( 
.A(n_1103),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1089),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1135),
.A2(n_1139),
.B1(n_1143),
.B2(n_1128),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1128),
.A2(n_1131),
.B1(n_1142),
.B2(n_1148),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1142),
.B(n_1148),
.Y(n_1231)
);

CKINVDCx14_ASAP7_75t_R g1232 ( 
.A(n_1165),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1061),
.A2(n_690),
.B1(n_451),
.B2(n_452),
.Y(n_1233)
);

INVx6_ASAP7_75t_L g1234 ( 
.A(n_1114),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1053),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1157),
.A2(n_804),
.B1(n_1045),
.B2(n_693),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1114),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1057),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1114),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1053),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1100),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1063),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1112),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1141),
.A2(n_391),
.B1(n_1043),
.B2(n_1062),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1157),
.A2(n_627),
.B(n_623),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1061),
.A2(n_690),
.B1(n_451),
.B2(n_452),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1141),
.A2(n_391),
.B1(n_1043),
.B2(n_1062),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1045),
.A2(n_391),
.B1(n_1157),
.B2(n_913),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1061),
.A2(n_690),
.B1(n_693),
.B2(n_585),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1065),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1141),
.A2(n_391),
.B1(n_1043),
.B2(n_1062),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1114),
.Y(n_1252)
);

CKINVDCx11_ASAP7_75t_R g1253 ( 
.A(n_1053),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1053),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1053),
.Y(n_1255)
);

CKINVDCx11_ASAP7_75t_R g1256 ( 
.A(n_1053),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1141),
.A2(n_391),
.B1(n_1043),
.B2(n_1062),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1053),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1112),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1061),
.A2(n_690),
.B1(n_391),
.B2(n_368),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1219),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1198),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1232),
.B(n_1180),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1231),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1180),
.B(n_1168),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1206),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1248),
.A2(n_1207),
.B(n_1167),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1205),
.A2(n_1211),
.B(n_1171),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1228),
.A2(n_1224),
.B1(n_1236),
.B2(n_1247),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1183),
.Y(n_1270)
);

AND2x2_ASAP7_75t_SL g1271 ( 
.A(n_1175),
.B(n_1225),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1223),
.A2(n_1209),
.B(n_1229),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1254),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1209),
.A2(n_1210),
.B(n_1226),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1194),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1220),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1230),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1230),
.Y(n_1278)
);

BUFx4f_ASAP7_75t_L g1279 ( 
.A(n_1214),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1238),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1206),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1222),
.Y(n_1282)
);

NAND2x1_ASAP7_75t_L g1283 ( 
.A(n_1213),
.B(n_1217),
.Y(n_1283)
);

CKINVDCx11_ASAP7_75t_R g1284 ( 
.A(n_1235),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1224),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1227),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1214),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1215),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1215),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1202),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1218),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1221),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1182),
.B(n_1178),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1221),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1199),
.B(n_1171),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1205),
.Y(n_1296)
);

BUFx12f_ASAP7_75t_L g1297 ( 
.A(n_1253),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1169),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1212),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1182),
.B(n_1178),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1199),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1175),
.B(n_1186),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1181),
.B(n_1186),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1181),
.B(n_1192),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1217),
.A2(n_1201),
.B(n_1216),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1242),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1192),
.B(n_1201),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1196),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1197),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1212),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1244),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1244),
.A2(n_1257),
.B(n_1251),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1237),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1252),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1208),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1247),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1251),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1257),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1193),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1245),
.B(n_1184),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1203),
.B(n_1190),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1233),
.A2(n_1246),
.B(n_1260),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1267),
.A2(n_1249),
.B(n_1243),
.C(n_1179),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1282),
.B(n_1250),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_SL g1325 ( 
.A1(n_1315),
.A2(n_1188),
.B(n_1189),
.C(n_1256),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1306),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1301),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1273),
.B(n_1259),
.Y(n_1328)
);

AO21x1_ASAP7_75t_L g1329 ( 
.A1(n_1304),
.A2(n_1187),
.B(n_1259),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1268),
.A2(n_1260),
.B(n_1187),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1274),
.A2(n_1239),
.B(n_1234),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1301),
.B(n_1173),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1280),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1269),
.A2(n_1177),
.B(n_1204),
.C(n_1200),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1304),
.A2(n_1172),
.B(n_1255),
.C(n_1240),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1279),
.B(n_1176),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1262),
.B(n_1170),
.Y(n_1337)
);

AO32x2_ASAP7_75t_L g1338 ( 
.A1(n_1287),
.A2(n_1170),
.A3(n_1241),
.B1(n_1195),
.B2(n_1176),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1312),
.A2(n_1239),
.B1(n_1191),
.B2(n_1185),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1263),
.B(n_1241),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1263),
.B(n_1265),
.Y(n_1341)
);

OR2x6_ASAP7_75t_L g1342 ( 
.A(n_1305),
.B(n_1174),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1265),
.B(n_1258),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1270),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1297),
.Y(n_1345)
);

NAND4xp25_ASAP7_75t_L g1346 ( 
.A(n_1302),
.B(n_1300),
.C(n_1293),
.D(n_1303),
.Y(n_1346)
);

AO32x2_ASAP7_75t_L g1347 ( 
.A1(n_1287),
.A2(n_1310),
.A3(n_1299),
.B1(n_1295),
.B2(n_1308),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1295),
.A2(n_1293),
.B(n_1300),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1282),
.B(n_1285),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1291),
.A2(n_1274),
.B(n_1305),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1321),
.B(n_1285),
.Y(n_1351)
);

AO32x2_ASAP7_75t_L g1352 ( 
.A1(n_1299),
.A2(n_1310),
.A3(n_1308),
.B1(n_1312),
.B2(n_1319),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1320),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1286),
.B(n_1313),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1319),
.A2(n_1302),
.B(n_1309),
.C(n_1312),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1296),
.A2(n_1272),
.B(n_1283),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1303),
.A2(n_1271),
.B1(n_1322),
.B2(n_1307),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1264),
.B(n_1296),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1321),
.B(n_1298),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1313),
.B(n_1314),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1290),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_1320),
.Y(n_1362)
);

CKINVDCx6p67_ASAP7_75t_R g1363 ( 
.A(n_1297),
.Y(n_1363)
);

AO32x2_ASAP7_75t_L g1364 ( 
.A1(n_1266),
.A2(n_1277),
.A3(n_1278),
.B1(n_1288),
.B2(n_1289),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1314),
.B(n_1276),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1315),
.B(n_1284),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1341),
.B(n_1272),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1361),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1333),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1353),
.B(n_1266),
.Y(n_1370)
);

BUFx2_ASAP7_75t_SL g1371 ( 
.A(n_1329),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1347),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1344),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1340),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1339),
.B(n_1271),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1347),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1346),
.A2(n_1318),
.B1(n_1311),
.B2(n_1317),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1347),
.B(n_1272),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1350),
.B(n_1272),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1350),
.B(n_1281),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1365),
.B(n_1261),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1362),
.B(n_1281),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1346),
.A2(n_1322),
.B1(n_1307),
.B2(n_1317),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1327),
.B(n_1358),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1354),
.B(n_1261),
.Y(n_1385)
);

CKINVDCx16_ASAP7_75t_R g1386 ( 
.A(n_1345),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1360),
.B(n_1292),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1326),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1349),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1364),
.B(n_1294),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1364),
.Y(n_1391)
);

OAI31xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1377),
.A2(n_1348),
.A3(n_1343),
.B(n_1351),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1389),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1379),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1379),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_L g1396 ( 
.A(n_1372),
.B(n_1356),
.C(n_1348),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1372),
.B(n_1376),
.Y(n_1397)
);

INVxp67_ASAP7_75t_SL g1398 ( 
.A(n_1380),
.Y(n_1398)
);

AO22x1_ASAP7_75t_L g1399 ( 
.A1(n_1378),
.A2(n_1318),
.B1(n_1316),
.B2(n_1311),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1372),
.B(n_1357),
.C(n_1355),
.Y(n_1400)
);

INVx5_ASAP7_75t_L g1401 ( 
.A(n_1379),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1367),
.B(n_1352),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1380),
.Y(n_1403)
);

OAI31xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1377),
.A2(n_1316),
.A3(n_1275),
.B(n_1359),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1367),
.B(n_1352),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1382),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1367),
.B(n_1352),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1389),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1369),
.Y(n_1409)
);

NOR2x1_ASAP7_75t_SL g1410 ( 
.A(n_1371),
.B(n_1375),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1369),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1376),
.B(n_1364),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1376),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1378),
.A2(n_1331),
.B(n_1357),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1389),
.B(n_1339),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1370),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1382),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1373),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1390),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1390),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1373),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1390),
.Y(n_1422)
);

AOI211x1_ASAP7_75t_SL g1423 ( 
.A1(n_1375),
.A2(n_1335),
.B(n_1334),
.C(n_1330),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1383),
.A2(n_1288),
.B1(n_1289),
.B2(n_1332),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1381),
.B(n_1385),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1418),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1418),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1421),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1419),
.B(n_1374),
.Y(n_1429)
);

OR2x6_ASAP7_75t_L g1430 ( 
.A(n_1399),
.B(n_1342),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1394),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1394),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1419),
.B(n_1374),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1419),
.B(n_1387),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1421),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1406),
.Y(n_1436)
);

INVx5_ASAP7_75t_L g1437 ( 
.A(n_1401),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1409),
.B(n_1368),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1406),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1409),
.B(n_1368),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1411),
.B(n_1391),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1419),
.B(n_1387),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1401),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1394),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1411),
.B(n_1384),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1394),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1401),
.B(n_1403),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1401),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1417),
.B(n_1384),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1397),
.B(n_1370),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1397),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1397),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1438),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1451),
.B(n_1412),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1437),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1431),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1429),
.B(n_1413),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1429),
.B(n_1413),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1429),
.B(n_1413),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1431),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1438),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1431),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1437),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1426),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1440),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1426),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1433),
.B(n_1425),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1433),
.B(n_1425),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1452),
.B(n_1412),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1437),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1450),
.B(n_1416),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1430),
.A2(n_1400),
.B1(n_1396),
.B2(n_1424),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1427),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1427),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1428),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1428),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1450),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1445),
.B(n_1412),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1435),
.Y(n_1480)
);

NAND2x1_ASAP7_75t_L g1481 ( 
.A(n_1448),
.B(n_1403),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1435),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1432),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1445),
.B(n_1420),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1449),
.B(n_1416),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1436),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1433),
.B(n_1425),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1436),
.Y(n_1488)
);

NOR2x1_ASAP7_75t_L g1489 ( 
.A(n_1448),
.B(n_1366),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1432),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1439),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1434),
.B(n_1393),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1440),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1439),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1494),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1493),
.B(n_1423),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1457),
.Y(n_1497)
);

AOI33xp33_ASAP7_75t_L g1498 ( 
.A1(n_1473),
.A2(n_1493),
.A3(n_1460),
.B1(n_1459),
.B2(n_1458),
.B3(n_1491),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1489),
.B(n_1437),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1465),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1478),
.B(n_1423),
.Y(n_1501)
);

INVx3_ASAP7_75t_SL g1502 ( 
.A(n_1456),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_SL g1503 ( 
.A(n_1489),
.B(n_1363),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1453),
.B(n_1392),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1472),
.B(n_1449),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1465),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1481),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1462),
.B(n_1386),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1467),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1467),
.Y(n_1510)
);

NOR2x1_ASAP7_75t_L g1511 ( 
.A(n_1456),
.B(n_1315),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1466),
.B(n_1386),
.Y(n_1512)
);

INVxp67_ASAP7_75t_SL g1513 ( 
.A(n_1456),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1458),
.B(n_1392),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1492),
.B(n_1434),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1485),
.B(n_1325),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1457),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1485),
.B(n_1328),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1459),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1460),
.B(n_1402),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1492),
.B(n_1434),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1468),
.B(n_1442),
.Y(n_1522)
);

INVx1_ASAP7_75t_SL g1523 ( 
.A(n_1472),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1479),
.A2(n_1396),
.B1(n_1400),
.B2(n_1398),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1455),
.B(n_1441),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1456),
.B(n_1437),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1464),
.B(n_1437),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1474),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1455),
.B(n_1441),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1500),
.Y(n_1530)
);

OA211x2_ASAP7_75t_L g1531 ( 
.A1(n_1503),
.A2(n_1481),
.B(n_1470),
.C(n_1454),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1496),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1501),
.A2(n_1410),
.B(n_1404),
.Y(n_1533)
);

AOI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1524),
.A2(n_1504),
.B1(n_1514),
.B2(n_1523),
.C(n_1512),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1498),
.A2(n_1404),
.B(n_1407),
.C(n_1405),
.Y(n_1535)
);

XOR2x1_ASAP7_75t_L g1536 ( 
.A(n_1499),
.B(n_1324),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_1519),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1506),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1498),
.B(n_1454),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1515),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1518),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1518),
.B(n_1479),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1509),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1510),
.Y(n_1544)
);

AOI321xp33_ASAP7_75t_L g1545 ( 
.A1(n_1520),
.A2(n_1424),
.A3(n_1383),
.B1(n_1470),
.B2(n_1402),
.C(n_1405),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1528),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1495),
.A2(n_1398),
.B(n_1422),
.C(n_1420),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1515),
.Y(n_1548)
);

OAI32xp33_ASAP7_75t_L g1549 ( 
.A1(n_1499),
.A2(n_1484),
.A3(n_1448),
.B1(n_1447),
.B2(n_1422),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1497),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1505),
.B(n_1484),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1497),
.Y(n_1552)
);

AOI32xp33_ASAP7_75t_L g1553 ( 
.A1(n_1516),
.A2(n_1402),
.A3(n_1405),
.B1(n_1407),
.B2(n_1447),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1508),
.B(n_1486),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1541),
.B(n_1508),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1532),
.B(n_1512),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1532),
.B(n_1521),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1550),
.Y(n_1558)
);

NOR2xp67_ASAP7_75t_L g1559 ( 
.A(n_1540),
.B(n_1507),
.Y(n_1559)
);

AOI32xp33_ASAP7_75t_L g1560 ( 
.A1(n_1534),
.A2(n_1516),
.A3(n_1525),
.B1(n_1529),
.B2(n_1511),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1548),
.Y(n_1561)
);

OAI31xp33_ASAP7_75t_L g1562 ( 
.A1(n_1535),
.A2(n_1407),
.A3(n_1517),
.B(n_1526),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1537),
.B(n_1522),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1539),
.B(n_1542),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1533),
.A2(n_1513),
.B(n_1527),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1534),
.A2(n_1517),
.B1(n_1322),
.B2(n_1461),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1551),
.B(n_1468),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1552),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1536),
.B(n_1469),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1554),
.B(n_1469),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1533),
.A2(n_1430),
.B1(n_1399),
.B2(n_1414),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1530),
.Y(n_1572)
);

AOI32xp33_ASAP7_75t_L g1573 ( 
.A1(n_1545),
.A2(n_1447),
.A3(n_1395),
.B1(n_1507),
.B2(n_1448),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1573),
.A2(n_1531),
.B1(n_1553),
.B2(n_1526),
.Y(n_1574)
);

NOR2x1_ASAP7_75t_L g1575 ( 
.A(n_1556),
.B(n_1507),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1563),
.B(n_1538),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1565),
.A2(n_1527),
.B(n_1549),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1569),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1557),
.Y(n_1579)
);

OAI32xp33_ASAP7_75t_L g1580 ( 
.A1(n_1564),
.A2(n_1546),
.A3(n_1544),
.B1(n_1543),
.B2(n_1443),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1555),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_SL g1582 ( 
.A1(n_1564),
.A2(n_1547),
.B1(n_1476),
.B2(n_1475),
.C(n_1480),
.Y(n_1582)
);

NAND4xp75_ASAP7_75t_L g1583 ( 
.A(n_1562),
.B(n_1471),
.C(n_1464),
.D(n_1415),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1561),
.Y(n_1584)
);

NOR3xp33_ASAP7_75t_L g1585 ( 
.A(n_1581),
.B(n_1561),
.C(n_1560),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1584),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_SL g1587 ( 
.A(n_1577),
.B(n_1566),
.C(n_1571),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1583),
.A2(n_1569),
.B(n_1559),
.Y(n_1588)
);

NOR2x1_ASAP7_75t_L g1589 ( 
.A(n_1575),
.B(n_1558),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1574),
.B(n_1570),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1582),
.A2(n_1566),
.B1(n_1568),
.B2(n_1572),
.C(n_1547),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1578),
.Y(n_1592)
);

NOR3x1_ASAP7_75t_SL g1593 ( 
.A(n_1579),
.B(n_1388),
.C(n_1570),
.Y(n_1593)
);

OAI21xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1589),
.A2(n_1567),
.B(n_1576),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1593),
.A2(n_1582),
.B(n_1487),
.Y(n_1595)
);

AOI21xp33_ASAP7_75t_L g1596 ( 
.A1(n_1592),
.A2(n_1580),
.B(n_1461),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_SL g1597 ( 
.A(n_1585),
.B(n_1336),
.C(n_1323),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1586),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1595),
.A2(n_1587),
.B(n_1590),
.C(n_1591),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1598),
.A2(n_1502),
.B1(n_1596),
.B2(n_1486),
.Y(n_1600)
);

NAND4xp75_ASAP7_75t_SL g1601 ( 
.A(n_1594),
.B(n_1588),
.C(n_1597),
.D(n_1502),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1595),
.A2(n_1471),
.B(n_1490),
.C(n_1457),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1598),
.Y(n_1603)
);

OAI21xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1595),
.A2(n_1487),
.B(n_1491),
.Y(n_1604)
);

XOR2xp5_ASAP7_75t_L g1605 ( 
.A(n_1601),
.B(n_1324),
.Y(n_1605)
);

XNOR2xp5_ASAP7_75t_L g1606 ( 
.A(n_1600),
.B(n_1430),
.Y(n_1606)
);

NAND4xp25_ASAP7_75t_L g1607 ( 
.A(n_1599),
.B(n_1443),
.C(n_1408),
.D(n_1393),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1604),
.A2(n_1490),
.B1(n_1483),
.B2(n_1461),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1603),
.Y(n_1609)
);

NOR3xp33_ASAP7_75t_L g1610 ( 
.A(n_1609),
.B(n_1602),
.C(n_1483),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1607),
.A2(n_1483),
.B(n_1463),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1606),
.A2(n_1490),
.B1(n_1463),
.B2(n_1488),
.C(n_1480),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1610),
.A2(n_1605),
.B1(n_1608),
.B2(n_1463),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1613),
.A2(n_1611),
.B1(n_1612),
.B2(n_1488),
.Y(n_1614)
);

XOR2x2_ASAP7_75t_L g1615 ( 
.A(n_1614),
.B(n_1410),
.Y(n_1615)
);

AOI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1614),
.A2(n_1475),
.B(n_1474),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1616),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1615),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1617),
.B(n_1476),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1618),
.A2(n_1482),
.B(n_1477),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1619),
.A2(n_1482),
.B(n_1477),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1621),
.B(n_1620),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1622),
.Y(n_1623)
);

AOI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1623),
.A2(n_1432),
.B1(n_1446),
.B2(n_1444),
.C(n_1443),
.Y(n_1624)
);

AOI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1624),
.A2(n_1338),
.B(n_1337),
.C(n_1443),
.Y(n_1625)
);


endmodule