module real_aes_6883_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_L g436 ( .A1(n_0), .A2(n_7), .B1(n_437), .B2(n_708), .C1(n_713), .C2(n_714), .Y(n_436) );
NAND3xp33_ASAP7_75t_SL g102 ( .A(n_1), .B(n_103), .C(n_104), .Y(n_102) );
INVx1_ASAP7_75t_L g431 ( .A(n_1), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_2), .A2(n_138), .B(n_143), .C(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_3), .A2(n_133), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g449 ( .A(n_4), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_5), .B(n_157), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_6), .B(n_433), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_7), .Y(n_713) );
AOI21xp33_ASAP7_75t_L g466 ( .A1(n_8), .A2(n_133), .B(n_467), .Y(n_466) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g167 ( .A(n_10), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_11), .B(n_43), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_12), .A2(n_245), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_13), .B(n_148), .Y(n_184) );
INVx1_ASAP7_75t_L g471 ( .A(n_14), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_15), .B(n_147), .Y(n_519) );
INVx1_ASAP7_75t_L g131 ( .A(n_16), .Y(n_131) );
INVx1_ASAP7_75t_L g531 ( .A(n_17), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_18), .A2(n_168), .B(n_193), .C(n_195), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_19), .B(n_157), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_20), .B(n_460), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_21), .B(n_133), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_22), .B(n_253), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_23), .A2(n_147), .B(n_149), .C(n_153), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_24), .B(n_157), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_25), .B(n_148), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_26), .A2(n_151), .B(n_195), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_27), .B(n_148), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_28), .Y(n_213) );
INVx1_ASAP7_75t_L g227 ( .A(n_29), .Y(n_227) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_30), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_31), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_32), .B(n_148), .Y(n_450) );
INVx1_ASAP7_75t_L g250 ( .A(n_33), .Y(n_250) );
INVx1_ASAP7_75t_L g484 ( .A(n_34), .Y(n_484) );
INVx2_ASAP7_75t_L g136 ( .A(n_35), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_36), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_37), .A2(n_147), .B(n_206), .C(n_208), .Y(n_205) );
INVxp67_ASAP7_75t_L g251 ( .A(n_38), .Y(n_251) );
CKINVDCx14_ASAP7_75t_R g204 ( .A(n_39), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_40), .A2(n_143), .B(n_226), .C(n_232), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_41), .A2(n_138), .B(n_143), .C(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_42), .A2(n_116), .B1(n_117), .B2(n_424), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_42), .Y(n_424) );
INVx1_ASAP7_75t_L g483 ( .A(n_44), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_45), .A2(n_165), .B(n_166), .C(n_169), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_46), .B(n_148), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_47), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_48), .Y(n_247) );
INVx1_ASAP7_75t_L g141 ( .A(n_49), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g485 ( .A(n_50), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_51), .B(n_133), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_52), .A2(n_143), .B1(n_153), .B2(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_53), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_54), .Y(n_446) );
CKINVDCx14_ASAP7_75t_R g163 ( .A(n_55), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_56), .A2(n_165), .B(n_208), .C(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_57), .Y(n_512) );
INVx1_ASAP7_75t_L g468 ( .A(n_58), .Y(n_468) );
INVx1_ASAP7_75t_L g139 ( .A(n_59), .Y(n_139) );
INVx1_ASAP7_75t_L g130 ( .A(n_60), .Y(n_130) );
INVx1_ASAP7_75t_SL g207 ( .A(n_61), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_62), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_63), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g216 ( .A(n_64), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_SL g459 ( .A1(n_65), .A2(n_208), .B(n_460), .C(n_461), .Y(n_459) );
INVxp67_ASAP7_75t_L g462 ( .A(n_66), .Y(n_462) );
INVx1_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_68), .A2(n_133), .B(n_162), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_69), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_70), .A2(n_133), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_71), .Y(n_487) );
INVx1_ASAP7_75t_L g506 ( .A(n_72), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_73), .A2(n_245), .B(n_246), .Y(n_244) );
INVx1_ASAP7_75t_L g191 ( .A(n_74), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g224 ( .A(n_75), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_76), .A2(n_138), .B(n_143), .C(n_508), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_77), .A2(n_133), .B(n_140), .Y(n_132) );
INVx1_ASAP7_75t_L g194 ( .A(n_78), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_79), .B(n_228), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_80), .A2(n_100), .B1(n_109), .B2(n_719), .Y(n_99) );
INVx2_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
INVx1_ASAP7_75t_L g181 ( .A(n_82), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_83), .B(n_460), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_84), .A2(n_138), .B(n_143), .C(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g103 ( .A(n_85), .Y(n_103) );
OR2x2_ASAP7_75t_L g428 ( .A(n_85), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g707 ( .A(n_85), .B(n_430), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_86), .A2(n_143), .B(n_215), .C(n_218), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_87), .B(n_160), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_88), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_89), .A2(n_138), .B(n_143), .C(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_90), .Y(n_523) );
INVx1_ASAP7_75t_L g458 ( .A(n_91), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_92), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_93), .B(n_228), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_94), .B(n_126), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_95), .B(n_126), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_96), .B(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_98), .A2(n_133), .B(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_101), .Y(n_721) );
OR2x2_ASAP7_75t_SL g101 ( .A(n_102), .B(n_107), .Y(n_101) );
OR2x2_ASAP7_75t_L g706 ( .A(n_103), .B(n_430), .Y(n_706) );
NOR2x2_ASAP7_75t_L g716 ( .A(n_103), .B(n_429), .Y(n_716) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g430 ( .A(n_108), .B(n_431), .Y(n_430) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_114), .B(n_435), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g718 ( .A(n_113), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_425), .B(n_432), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g437 ( .A1(n_118), .A2(n_438), .B1(n_706), .B2(n_707), .Y(n_437) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g712 ( .A(n_119), .Y(n_712) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_350), .Y(n_119) );
NOR4xp25_ASAP7_75t_L g120 ( .A(n_121), .B(n_292), .C(n_322), .D(n_332), .Y(n_120) );
OAI211xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_197), .B(n_255), .C(n_282), .Y(n_121) );
OAI222xp33_ASAP7_75t_L g377 ( .A1(n_122), .A2(n_297), .B1(n_378), .B2(n_379), .C1(n_380), .C2(n_381), .Y(n_377) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_172), .Y(n_122) );
AOI33xp33_ASAP7_75t_L g303 ( .A1(n_123), .A2(n_290), .A3(n_291), .B1(n_304), .B2(n_309), .B3(n_311), .Y(n_303) );
OAI211xp5_ASAP7_75t_SL g360 ( .A1(n_123), .A2(n_361), .B(n_363), .C(n_365), .Y(n_360) );
OR2x2_ASAP7_75t_L g376 ( .A(n_123), .B(n_362), .Y(n_376) );
INVx1_ASAP7_75t_L g409 ( .A(n_123), .Y(n_409) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_159), .Y(n_123) );
INVx2_ASAP7_75t_L g286 ( .A(n_124), .Y(n_286) );
AND2x2_ASAP7_75t_L g302 ( .A(n_124), .B(n_188), .Y(n_302) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_124), .Y(n_337) );
AND2x2_ASAP7_75t_L g366 ( .A(n_124), .B(n_159), .Y(n_366) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_132), .B(n_156), .Y(n_124) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_125), .A2(n_189), .B(n_196), .Y(n_188) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_125), .A2(n_202), .B(n_210), .Y(n_201) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx4_ASAP7_75t_L g158 ( .A(n_126), .Y(n_158) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_126), .A2(n_456), .B(n_463), .Y(n_455) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g243 ( .A(n_127), .Y(n_243) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_128), .B(n_129), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
BUFx2_ASAP7_75t_L g245 ( .A(n_133), .Y(n_245) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_134), .B(n_138), .Y(n_178) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g231 ( .A(n_135), .Y(n_231) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx1_ASAP7_75t_L g154 ( .A(n_136), .Y(n_154) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_137), .Y(n_152) );
INVx3_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
INVx1_ASAP7_75t_L g460 ( .A(n_137), .Y(n_460) );
INVx4_ASAP7_75t_SL g155 ( .A(n_138), .Y(n_155) );
BUFx3_ASAP7_75t_L g232 ( .A(n_138), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_142), .B(n_146), .C(n_155), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_SL g162 ( .A1(n_142), .A2(n_155), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_142), .A2(n_155), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_142), .A2(n_155), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_SL g246 ( .A1(n_142), .A2(n_155), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_142), .A2(n_155), .B(n_458), .C(n_459), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_142), .A2(n_155), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_142), .A2(n_155), .B(n_528), .C(n_529), .Y(n_527) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_144), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_147), .B(n_207), .Y(n_206) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g165 ( .A(n_148), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_151), .B(n_194), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g249 ( .A1(n_151), .A2(n_228), .B1(n_250), .B2(n_251), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_151), .B(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
OAI22xp5_ASAP7_75t_SL g482 ( .A1(n_152), .A2(n_183), .B1(n_483), .B2(n_484), .Y(n_482) );
INVx2_ASAP7_75t_L g451 ( .A(n_153), .Y(n_451) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g218 ( .A(n_155), .Y(n_218) );
OAI22xp33_ASAP7_75t_L g480 ( .A1(n_155), .A2(n_178), .B1(n_481), .B2(n_485), .Y(n_480) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_157), .A2(n_466), .B(n_472), .Y(n_465) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_158), .B(n_187), .Y(n_186) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_158), .A2(n_212), .B(n_219), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_158), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_SL g502 ( .A(n_158), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g266 ( .A(n_159), .Y(n_266) );
BUFx3_ASAP7_75t_L g274 ( .A(n_159), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_159), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g285 ( .A(n_159), .B(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_159), .B(n_173), .Y(n_314) );
AND2x2_ASAP7_75t_L g383 ( .A(n_159), .B(n_317), .Y(n_383) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_171), .Y(n_159) );
INVx1_ASAP7_75t_L g175 ( .A(n_160), .Y(n_175) );
INVx2_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_160), .A2(n_178), .B(n_224), .C(n_225), .Y(n_223) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_160), .A2(n_526), .B(n_532), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx5_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_168), .B(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_168), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g195 ( .A(n_170), .Y(n_195) );
INVx2_ASAP7_75t_SL g277 ( .A(n_172), .Y(n_277) );
OR2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_188), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_173), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g319 ( .A(n_173), .Y(n_319) );
AND2x2_ASAP7_75t_L g330 ( .A(n_173), .B(n_286), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_173), .B(n_315), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_173), .B(n_317), .Y(n_362) );
AND2x2_ASAP7_75t_L g421 ( .A(n_173), .B(n_366), .Y(n_421) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g291 ( .A(n_174), .B(n_188), .Y(n_291) );
AND2x2_ASAP7_75t_L g301 ( .A(n_174), .B(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g323 ( .A(n_174), .Y(n_323) );
AND3x2_ASAP7_75t_L g382 ( .A(n_174), .B(n_383), .C(n_384), .Y(n_382) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_186), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_175), .B(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_175), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_175), .B(n_523), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_178), .A2(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_178), .A2(n_446), .B(n_447), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_178), .A2(n_506), .B(n_507), .Y(n_505) );
O2A1O1Ixp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_184), .C(n_185), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_182), .A2(n_185), .B(n_216), .C(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_185), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_185), .A2(n_509), .B(n_510), .Y(n_508) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_188), .Y(n_273) );
INVx1_ASAP7_75t_SL g317 ( .A(n_188), .Y(n_317) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_188), .B(n_266), .C(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_235), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_198), .A2(n_301), .B(n_353), .C(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_200), .B(n_222), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_200), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_SL g369 ( .A(n_200), .Y(n_369) );
AND2x2_ASAP7_75t_L g390 ( .A(n_200), .B(n_237), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_200), .B(n_299), .Y(n_418) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
AND2x2_ASAP7_75t_L g263 ( .A(n_201), .B(n_254), .Y(n_263) );
INVx2_ASAP7_75t_L g270 ( .A(n_201), .Y(n_270) );
AND2x2_ASAP7_75t_L g290 ( .A(n_201), .B(n_237), .Y(n_290) );
AND2x2_ASAP7_75t_L g340 ( .A(n_201), .B(n_222), .Y(n_340) );
INVx1_ASAP7_75t_L g344 ( .A(n_201), .Y(n_344) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_209), .Y(n_520) );
INVx2_ASAP7_75t_SL g254 ( .A(n_211), .Y(n_254) );
BUFx2_ASAP7_75t_L g280 ( .A(n_211), .Y(n_280) );
AND2x2_ASAP7_75t_L g407 ( .A(n_211), .B(n_222), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
INVx1_ASAP7_75t_L g253 ( .A(n_221), .Y(n_253) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_221), .A2(n_515), .B(n_522), .Y(n_514) );
INVx3_ASAP7_75t_SL g237 ( .A(n_222), .Y(n_237) );
AND2x2_ASAP7_75t_L g262 ( .A(n_222), .B(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g269 ( .A(n_222), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g299 ( .A(n_222), .B(n_259), .Y(n_299) );
OR2x2_ASAP7_75t_L g308 ( .A(n_222), .B(n_254), .Y(n_308) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_222), .Y(n_326) );
AND2x2_ASAP7_75t_L g331 ( .A(n_222), .B(n_284), .Y(n_331) );
AND2x2_ASAP7_75t_L g359 ( .A(n_222), .B(n_239), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_222), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g397 ( .A(n_222), .B(n_238), .Y(n_397) );
OR2x6_ASAP7_75t_L g222 ( .A(n_223), .B(n_233), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_229), .C(n_230), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_228), .A2(n_449), .B(n_450), .C(n_451), .Y(n_448) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_231), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_L g321 ( .A(n_237), .B(n_270), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_237), .B(n_263), .Y(n_349) );
AND2x2_ASAP7_75t_L g367 ( .A(n_237), .B(n_284), .Y(n_367) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_254), .Y(n_238) );
AND2x2_ASAP7_75t_L g268 ( .A(n_239), .B(n_254), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_239), .B(n_297), .Y(n_296) );
BUFx3_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
OR2x2_ASAP7_75t_L g354 ( .A(n_239), .B(n_274), .Y(n_354) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_244), .B(n_252), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_241), .A2(n_260), .B(n_261), .Y(n_259) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_241), .A2(n_505), .B(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_SL g496 ( .A1(n_242), .A2(n_497), .B(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_243), .A2(n_445), .B(n_452), .Y(n_444) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_243), .A2(n_480), .B(n_486), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_243), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g260 ( .A(n_244), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_252), .Y(n_261) );
AND2x2_ASAP7_75t_L g289 ( .A(n_254), .B(n_259), .Y(n_289) );
INVx1_ASAP7_75t_L g297 ( .A(n_254), .Y(n_297) );
AND2x2_ASAP7_75t_L g392 ( .A(n_254), .B(n_270), .Y(n_392) );
AOI222xp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_264), .B1(n_267), .B2(n_271), .C1(n_275), .C2(n_278), .Y(n_255) );
INVx1_ASAP7_75t_L g387 ( .A(n_256), .Y(n_387) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_262), .Y(n_256) );
AND2x2_ASAP7_75t_L g283 ( .A(n_257), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g294 ( .A(n_257), .B(n_263), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_257), .B(n_285), .Y(n_310) );
OAI222xp33_ASAP7_75t_L g332 ( .A1(n_257), .A2(n_333), .B1(n_338), .B2(n_339), .C1(n_347), .C2(n_349), .Y(n_332) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g320 ( .A(n_259), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_259), .B(n_340), .Y(n_380) );
AND2x2_ASAP7_75t_L g391 ( .A(n_259), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g399 ( .A(n_262), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_264), .B(n_315), .Y(n_378) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_266), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g336 ( .A(n_266), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx3_ASAP7_75t_L g281 ( .A(n_269), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g371 ( .A1(n_269), .A2(n_372), .B(n_375), .C(n_377), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_269), .B(n_306), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_269), .B(n_289), .Y(n_411) );
AND2x2_ASAP7_75t_L g284 ( .A(n_270), .B(n_280), .Y(n_284) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g311 ( .A(n_273), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_274), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g363 ( .A(n_274), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g402 ( .A(n_274), .B(n_302), .Y(n_402) );
INVx1_ASAP7_75t_L g414 ( .A(n_274), .Y(n_414) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_277), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g395 ( .A(n_280), .Y(n_395) );
A2O1A1Ixp33_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_285), .B(n_287), .C(n_291), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_283), .A2(n_313), .B1(n_328), .B2(n_331), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_284), .B(n_298), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_284), .B(n_306), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_285), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g348 ( .A(n_285), .Y(n_348) );
AND2x2_ASAP7_75t_L g355 ( .A(n_285), .B(n_335), .Y(n_355) );
INVx2_ASAP7_75t_L g316 ( .A(n_286), .Y(n_316) );
INVxp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NOR4xp25_ASAP7_75t_L g293 ( .A(n_290), .B(n_294), .C(n_295), .D(n_298), .Y(n_293) );
INVx1_ASAP7_75t_SL g364 ( .A(n_291), .Y(n_364) );
AND2x2_ASAP7_75t_L g408 ( .A(n_291), .B(n_409), .Y(n_408) );
OAI211xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_300), .B(n_303), .C(n_312), .Y(n_292) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_299), .B(n_369), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_301), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_419) );
INVx1_ASAP7_75t_SL g374 ( .A(n_302), .Y(n_374) );
AND2x2_ASAP7_75t_L g413 ( .A(n_302), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_306), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_310), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_311), .B(n_336), .Y(n_396) );
OAI21xp5_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_318), .B(n_320), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g388 ( .A(n_315), .Y(n_388) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_L g416 ( .A(n_316), .Y(n_416) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_317), .Y(n_343) );
OAI21xp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B(n_327), .Y(n_322) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_323), .Y(n_335) );
OR2x2_ASAP7_75t_L g373 ( .A(n_323), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI21xp33_ASAP7_75t_SL g368 ( .A1(n_326), .A2(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_330), .A2(n_357), .B1(n_360), .B2(n_367), .C(n_368), .Y(n_356) );
INVx1_ASAP7_75t_SL g400 ( .A(n_331), .Y(n_400) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
OR2x2_ASAP7_75t_L g347 ( .A(n_335), .B(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g384 ( .A(n_337), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_344), .B2(n_345), .Y(n_339) );
INVx1_ASAP7_75t_L g379 ( .A(n_340), .Y(n_379) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_343), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NOR4xp25_ASAP7_75t_L g350 ( .A(n_351), .B(n_385), .C(n_398), .D(n_410), .Y(n_350) );
NAND3xp33_ASAP7_75t_SL g351 ( .A(n_352), .B(n_356), .C(n_371), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_354), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_361), .B(n_366), .Y(n_370) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI221xp5_ASAP7_75t_SL g398 ( .A1(n_373), .A2(n_399), .B1(n_400), .B2(n_401), .C(n_403), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_375), .A2(n_390), .B(n_391), .C(n_393), .Y(n_389) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_376), .A2(n_394), .B1(n_396), .B2(n_397), .Y(n_393) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_388), .C(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g404 ( .A(n_397), .Y(n_404) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_405), .B(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_412), .B1(n_415), .B2(n_417), .C(n_419), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_428), .Y(n_434) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_432), .A2(n_436), .B(n_717), .Y(n_435) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g709 ( .A(n_438), .Y(n_709) );
NAND2x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_622), .Y(n_438) );
NOR5xp2_ASAP7_75t_L g439 ( .A(n_440), .B(n_545), .C(n_577), .D(n_592), .E(n_609), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_473), .B(n_492), .C(n_533), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_454), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_442), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_442), .B(n_597), .Y(n_660) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_443), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_443), .B(n_489), .Y(n_546) );
AND2x2_ASAP7_75t_L g587 ( .A(n_443), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_443), .B(n_556), .Y(n_591) );
OR2x2_ASAP7_75t_L g628 ( .A(n_443), .B(n_479), .Y(n_628) );
INVx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g478 ( .A(n_444), .B(n_479), .Y(n_478) );
INVx3_ASAP7_75t_L g536 ( .A(n_444), .Y(n_536) );
OR2x2_ASAP7_75t_L g699 ( .A(n_444), .B(n_539), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_454), .A2(n_602), .B1(n_603), .B2(n_606), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_454), .B(n_536), .Y(n_685) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_464), .Y(n_454) );
AND2x2_ASAP7_75t_L g491 ( .A(n_455), .B(n_479), .Y(n_491) );
AND2x2_ASAP7_75t_L g538 ( .A(n_455), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g543 ( .A(n_455), .Y(n_543) );
INVx3_ASAP7_75t_L g556 ( .A(n_455), .Y(n_556) );
OR2x2_ASAP7_75t_L g576 ( .A(n_455), .B(n_539), .Y(n_576) );
AND2x2_ASAP7_75t_L g595 ( .A(n_455), .B(n_465), .Y(n_595) );
BUFx2_ASAP7_75t_L g627 ( .A(n_455), .Y(n_627) );
AND2x4_ASAP7_75t_L g542 ( .A(n_464), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g477 ( .A(n_465), .Y(n_477) );
INVx2_ASAP7_75t_L g490 ( .A(n_465), .Y(n_490) );
OR2x2_ASAP7_75t_L g558 ( .A(n_465), .B(n_539), .Y(n_558) );
AND2x2_ASAP7_75t_L g588 ( .A(n_465), .B(n_479), .Y(n_588) );
AND2x2_ASAP7_75t_L g605 ( .A(n_465), .B(n_536), .Y(n_605) );
AND2x2_ASAP7_75t_L g645 ( .A(n_465), .B(n_556), .Y(n_645) );
AND2x2_ASAP7_75t_SL g681 ( .A(n_465), .B(n_491), .Y(n_681) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp33_ASAP7_75t_SL g474 ( .A(n_475), .B(n_488), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_476), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_477), .A2(n_491), .B(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_477), .B(n_479), .Y(n_675) );
AND2x2_ASAP7_75t_L g611 ( .A(n_478), .B(n_612), .Y(n_611) );
INVx3_ASAP7_75t_L g539 ( .A(n_479), .Y(n_539) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_479), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_488), .B(n_536), .Y(n_704) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_489), .A2(n_647), .B1(n_648), .B2(n_653), .Y(n_646) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AND2x2_ASAP7_75t_L g537 ( .A(n_490), .B(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g575 ( .A(n_490), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g612 ( .A(n_490), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_491), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g666 ( .A(n_491), .Y(n_666) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_513), .Y(n_493) );
INVx4_ASAP7_75t_L g552 ( .A(n_494), .Y(n_552) );
AND2x2_ASAP7_75t_L g630 ( .A(n_494), .B(n_597), .Y(n_630) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
INVx3_ASAP7_75t_L g549 ( .A(n_495), .Y(n_549) );
AND2x2_ASAP7_75t_L g563 ( .A(n_495), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g567 ( .A(n_495), .Y(n_567) );
INVx2_ASAP7_75t_L g581 ( .A(n_495), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_495), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g638 ( .A(n_495), .B(n_633), .Y(n_638) );
AND2x2_ASAP7_75t_L g703 ( .A(n_495), .B(n_673), .Y(n_703) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
AND2x2_ASAP7_75t_L g544 ( .A(n_504), .B(n_525), .Y(n_544) );
INVx2_ASAP7_75t_L g564 ( .A(n_504), .Y(n_564) );
INVx1_ASAP7_75t_L g569 ( .A(n_513), .Y(n_569) );
AND2x2_ASAP7_75t_L g615 ( .A(n_513), .B(n_563), .Y(n_615) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_524), .Y(n_513) );
INVx2_ASAP7_75t_L g554 ( .A(n_514), .Y(n_554) );
INVx1_ASAP7_75t_L g562 ( .A(n_514), .Y(n_562) );
AND2x2_ASAP7_75t_L g580 ( .A(n_514), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_514), .B(n_564), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_521), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
AND2x2_ASAP7_75t_L g597 ( .A(n_524), .B(n_554), .Y(n_597) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g550 ( .A(n_525), .Y(n_550) );
AND2x2_ASAP7_75t_L g633 ( .A(n_525), .B(n_564), .Y(n_633) );
OAI21xp5_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_540), .B(n_544), .Y(n_533) );
INVx1_ASAP7_75t_SL g578 ( .A(n_534), .Y(n_578) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_535), .B(n_542), .Y(n_635) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g584 ( .A(n_536), .B(n_539), .Y(n_584) );
AND2x2_ASAP7_75t_L g613 ( .A(n_536), .B(n_557), .Y(n_613) );
OR2x2_ASAP7_75t_L g616 ( .A(n_536), .B(n_576), .Y(n_616) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_537), .A2(n_629), .B1(n_681), .B2(n_682), .C1(n_684), .C2(n_686), .Y(n_680) );
BUFx2_ASAP7_75t_L g594 ( .A(n_539), .Y(n_594) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g583 ( .A(n_542), .B(n_584), .Y(n_583) );
INVx3_ASAP7_75t_SL g600 ( .A(n_542), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_542), .B(n_594), .Y(n_654) );
AND2x2_ASAP7_75t_L g589 ( .A(n_544), .B(n_549), .Y(n_589) );
INVx1_ASAP7_75t_L g608 ( .A(n_544), .Y(n_608) );
OAI221xp5_ASAP7_75t_SL g545 ( .A1(n_546), .A2(n_547), .B1(n_551), .B2(n_555), .C(n_559), .Y(n_545) );
OR2x2_ASAP7_75t_L g617 ( .A(n_547), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
AND2x2_ASAP7_75t_L g602 ( .A(n_549), .B(n_572), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_549), .B(n_562), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_549), .B(n_597), .Y(n_647) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_549), .Y(n_657) );
NAND2x1_ASAP7_75t_SL g668 ( .A(n_549), .B(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g553 ( .A(n_550), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g573 ( .A(n_550), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_550), .B(n_568), .Y(n_599) );
INVx1_ASAP7_75t_L g665 ( .A(n_550), .Y(n_665) );
INVx1_ASAP7_75t_L g640 ( .A(n_551), .Y(n_640) );
OR2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g652 ( .A(n_552), .Y(n_652) );
NOR2xp67_ASAP7_75t_L g664 ( .A(n_552), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g669 ( .A(n_553), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_553), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g572 ( .A(n_554), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_554), .B(n_564), .Y(n_585) );
INVx1_ASAP7_75t_L g651 ( .A(n_554), .Y(n_651) );
INVx1_ASAP7_75t_L g672 ( .A(n_555), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI21xp5_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_565), .B(n_574), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
AND2x2_ASAP7_75t_L g705 ( .A(n_561), .B(n_638), .Y(n_705) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g673 ( .A(n_562), .B(n_633), .Y(n_673) );
AOI32xp33_ASAP7_75t_L g586 ( .A1(n_563), .A2(n_569), .A3(n_587), .B1(n_589), .B2(n_590), .Y(n_586) );
AOI322xp5_ASAP7_75t_L g688 ( .A1(n_563), .A2(n_595), .A3(n_678), .B1(n_689), .B2(n_690), .C1(n_691), .C2(n_693), .Y(n_688) );
INVx2_ASAP7_75t_L g568 ( .A(n_564), .Y(n_568) );
INVx1_ASAP7_75t_L g678 ( .A(n_564), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_566), .B(n_572), .Y(n_621) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_567), .B(n_633), .Y(n_683) );
INVx1_ASAP7_75t_L g570 ( .A(n_568), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_568), .B(n_597), .Y(n_687) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_576), .B(n_671), .Y(n_670) );
OAI221xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_579), .B1(n_582), .B2(n_585), .C(n_586), .Y(n_577) );
OR2x2_ASAP7_75t_L g598 ( .A(n_579), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g607 ( .A(n_579), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g632 ( .A(n_580), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g636 ( .A(n_590), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_596), .B1(n_598), .B2(n_600), .C(n_601), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_594), .A2(n_625), .B1(n_629), .B2(n_630), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_595), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g700 ( .A(n_595), .Y(n_700) );
INVx1_ASAP7_75t_L g694 ( .A(n_597), .Y(n_694) );
INVx1_ASAP7_75t_SL g629 ( .A(n_598), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_600), .B(n_628), .Y(n_690) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_605), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g671 ( .A(n_605), .Y(n_671) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
OAI221xp5_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_614), .B1(n_616), .B2(n_617), .C(n_619), .Y(n_609) );
NOR2xp33_ASAP7_75t_SL g610 ( .A(n_611), .B(n_613), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_611), .A2(n_629), .B1(n_675), .B2(n_676), .Y(n_674) );
CKINVDCx14_ASAP7_75t_R g614 ( .A(n_615), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_616), .A2(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR3xp33_ASAP7_75t_SL g622 ( .A(n_623), .B(n_655), .C(n_679), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_631), .C(n_639), .D(n_646), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g702 ( .A(n_627), .Y(n_702) );
INVx3_ASAP7_75t_SL g696 ( .A(n_628), .Y(n_696) );
OR2x2_ASAP7_75t_L g701 ( .A(n_628), .B(n_702), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B1(n_636), .B2(n_638), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_633), .B(n_651), .Y(n_692) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_641), .B(n_643), .Y(n_639) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI211xp5_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_658), .B(n_661), .C(n_674), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g689 ( .A(n_660), .Y(n_689) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_666), .B1(n_667), .B2(n_670), .C1(n_672), .C2(n_673), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND4xp25_ASAP7_75t_SL g698 ( .A(n_671), .B(n_699), .C(n_700), .D(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND3xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_688), .C(n_697), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_706), .A2(n_709), .B1(n_710), .B2(n_712), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_707), .Y(n_711) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
endmodule