module fake_netlist_5_933_n_139 (n_16, n_0, n_12, n_9, n_25, n_18, n_22, n_1, n_8, n_10, n_24, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_139);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_139;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_124;
wire n_86;
wire n_136;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_101;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_128;
wire n_73;
wire n_92;
wire n_120;
wire n_135;
wire n_30;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_29;
wire n_79;
wire n_131;
wire n_47;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_118;
wire n_28;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_1),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g66 ( 
.A(n_30),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_28),
.B(n_4),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_45),
.B1(n_29),
.B2(n_43),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_47),
.B1(n_28),
.B2(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_55),
.Y(n_73)
);

INVxp67_ASAP7_75t_SL g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_12),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_25),
.B(n_67),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_65),
.B(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_63),
.B1(n_62),
.B2(n_53),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_79),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_78),
.B(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_81),
.Y(n_96)
);

NAND4xp25_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_69),
.C(n_80),
.D(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_82),
.Y(n_98)
);

OA21x2_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_83),
.B(n_88),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_91),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_94),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_97),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_76),
.B1(n_90),
.B2(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

NOR2xp67_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_106),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_108),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_75),
.C(n_49),
.Y(n_117)
);

NAND4xp75_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_105),
.C(n_52),
.D(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_116),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_52),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_54),
.Y(n_126)
);

AO22x2_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_59),
.B1(n_65),
.B2(n_56),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_76),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_50),
.Y(n_129)
);

NOR2x1p5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_59),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_56),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_61),
.B(n_83),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_61),
.B1(n_50),
.B2(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_61),
.B(n_58),
.C(n_89),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_126),
.B(n_127),
.Y(n_136)
);

OAI21x1_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_130),
.B(n_127),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_133),
.C(n_135),
.Y(n_138)
);

OAI221xp5_ASAP7_75t_R g139 ( 
.A1(n_138),
.A2(n_137),
.B1(n_131),
.B2(n_61),
.C(n_58),
.Y(n_139)
);


endmodule