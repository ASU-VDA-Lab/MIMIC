module fake_jpeg_17730_n_333 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_43),
.B(n_68),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_49),
.Y(n_82)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_14),
.B(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_57),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_0),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_0),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_62),
.Y(n_100)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_28),
.Y(n_71)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_65),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_21),
.B(n_5),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_67),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_68),
.B1(n_64),
.B2(n_40),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_70),
.A2(n_87),
.B1(n_91),
.B2(n_99),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_71),
.B(n_107),
.Y(n_139)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_109),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_27),
.B(n_26),
.C(n_28),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_74),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_75),
.B(n_83),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_32),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_46),
.B1(n_45),
.B2(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_47),
.A2(n_37),
.B1(n_20),
.B2(n_35),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_92),
.B(n_94),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_37),
.B1(n_20),
.B2(n_35),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_93),
.A2(n_95),
.B1(n_117),
.B2(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_24),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_18),
.B1(n_15),
.B2(n_38),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_96),
.B(n_105),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_61),
.A2(n_18),
.B1(n_15),
.B2(n_38),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_32),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g106 ( 
.A(n_42),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_32),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_54),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g110 ( 
.A(n_57),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_112),
.Y(n_123)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

CKINVDCx12_ASAP7_75t_R g112 ( 
.A(n_57),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_59),
.A2(n_9),
.B1(n_11),
.B2(n_2),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_54),
.A2(n_32),
.B1(n_24),
.B2(n_3),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_57),
.B(n_0),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_24),
.Y(n_124)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_167),
.Y(n_168)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_1),
.B(n_3),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_126),
.A2(n_153),
.B(n_139),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_154),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_7),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_129),
.B(n_140),
.Y(n_185)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_76),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_131),
.A2(n_145),
.B1(n_146),
.B2(n_149),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_143),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_11),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_142),
.C(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_78),
.B(n_108),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_82),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_104),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_147),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_99),
.B1(n_116),
.B2(n_103),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_150),
.Y(n_181)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_87),
.C(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_119),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_91),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_160),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_79),
.Y(n_160)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_125),
.Y(n_190)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_101),
.B(n_97),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_134),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_89),
.B(n_111),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_166),
.B(n_81),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_80),
.B(n_77),
.C(n_120),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_80),
.B1(n_81),
.B2(n_101),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_186),
.B1(n_195),
.B2(n_157),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_171),
.B(n_178),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_133),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_154),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_176),
.A2(n_201),
.B(n_203),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_127),
.A2(n_142),
.B1(n_152),
.B2(n_156),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_123),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_180),
.B(n_191),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_136),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_168),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_137),
.B1(n_167),
.B2(n_128),
.Y(n_186)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_139),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_137),
.A2(n_151),
.B1(n_163),
.B2(n_145),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_135),
.B(n_176),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_200),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_162),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_198),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_126),
.Y(n_200)
);

NAND2x1_ASAP7_75t_SL g201 ( 
.A(n_130),
.B(n_122),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_175),
.Y(n_233)
);

NAND2x1_ASAP7_75t_SL g203 ( 
.A(n_138),
.B(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_199),
.B1(n_194),
.B2(n_182),
.Y(n_245)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_212),
.Y(n_240)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_132),
.B1(n_135),
.B2(n_189),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_231),
.B1(n_233),
.B2(n_179),
.Y(n_248)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_230),
.B(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_218),
.Y(n_261)
);

CKINVDCx12_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_220),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_188),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_222),
.C(n_201),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_183),
.Y(n_222)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_222),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_202),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_208),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_168),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_203),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_169),
.A2(n_168),
.B1(n_176),
.B2(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_187),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_236),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_242),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_177),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_199),
.B(n_182),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_259),
.B1(n_236),
.B2(n_211),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_194),
.C(n_179),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_255),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_262),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_259),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_224),
.A2(n_216),
.B1(n_231),
.B2(n_214),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_263),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_206),
.A2(n_224),
.B1(n_218),
.B2(n_215),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_223),
.A2(n_209),
.B(n_213),
.Y(n_262)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_228),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_266),
.A2(n_268),
.B1(n_280),
.B2(n_245),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_212),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_207),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_207),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_232),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_282),
.B1(n_284),
.B2(n_276),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_235),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_283),
.C(n_246),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_261),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_265),
.Y(n_298)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_286),
.C(n_287),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_238),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_258),
.C(n_260),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_294),
.C(n_296),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_258),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_260),
.C(n_261),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_266),
.A2(n_251),
.B1(n_270),
.B2(n_267),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_264),
.Y(n_301)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_265),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_291),
.B1(n_293),
.B2(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_304),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_277),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_275),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_308),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_286),
.B(n_275),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_303),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_294),
.B(n_285),
.CI(n_296),
.CON(n_307),
.SN(n_307)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_309),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_297),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_292),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_310),
.Y(n_318)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_303),
.C(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_311),
.B(n_316),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_301),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

INVx13_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_318),
.B1(n_312),
.B2(n_314),
.Y(n_327)
);

OAI21x1_ASAP7_75t_SL g329 ( 
.A1(n_327),
.A2(n_328),
.B(n_321),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_319),
.Y(n_328)
);

A2O1A1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_329),
.A2(n_330),
.B(n_326),
.C(n_328),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_327),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_322),
.B1(n_313),
.B2(n_315),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_313),
.Y(n_333)
);


endmodule