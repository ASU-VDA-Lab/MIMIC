module fake_jpeg_2189_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_6),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_1),
.B(n_2),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_3),
.B(n_4),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_12),
.B1(n_16),
.B2(n_18),
.Y(n_54)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_12),
.B1(n_24),
.B2(n_16),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_56),
.B1(n_33),
.B2(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_38),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_32),
.A2(n_3),
.B1(n_4),
.B2(n_9),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_10),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_60),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_64),
.B1(n_65),
.B2(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_11),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_66),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_29),
.B1(n_26),
.B2(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_11),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_69),
.B(n_54),
.Y(n_76)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_31),
.A3(n_41),
.B1(n_26),
.B2(n_40),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_54),
.C(n_53),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_54),
.B1(n_40),
.B2(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_67),
.C(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_84),
.Y(n_88)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_61),
.B(n_66),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_77),
.B(n_72),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_87),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_89),
.A2(n_90),
.B(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_92),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_90),
.A2(n_84),
.B(n_75),
.C(n_78),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_94),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_98),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_96),
.A3(n_93),
.B1(n_89),
.B2(n_74),
.C1(n_30),
.C2(n_47),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_74),
.B1(n_47),
.B2(n_52),
.Y(n_100)
);

OAI211xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_44),
.B(n_52),
.C(n_95),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_44),
.Y(n_102)
);


endmodule