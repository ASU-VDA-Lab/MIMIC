module fake_jpeg_10572_n_293 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_23),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_21),
.B1(n_34),
.B2(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_48),
.B1(n_53),
.B2(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_34),
.B1(n_18),
.B2(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_50),
.B(n_54),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_34),
.B1(n_18),
.B2(n_19),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_27),
.B(n_33),
.C(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_43),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_19),
.B1(n_24),
.B2(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_20),
.B(n_17),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_17),
.A3(n_29),
.B1(n_30),
.B2(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_65),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_32),
.B1(n_31),
.B2(n_17),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_98),
.B(n_8),
.Y(n_116)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_75),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_32),
.B1(n_17),
.B2(n_24),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_70),
.A2(n_86),
.B(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_88),
.B1(n_100),
.B2(n_49),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_96),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_23),
.B(n_2),
.C(n_3),
.Y(n_113)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_79),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_43),
.C(n_42),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_3),
.C(n_4),
.Y(n_123)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_89),
.Y(n_103)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_0),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_30),
.B1(n_26),
.B2(n_29),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_23),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_26),
.B1(n_43),
.B2(n_41),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_62),
.B1(n_49),
.B2(n_64),
.Y(n_104)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_44),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_64),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_42),
.B1(n_41),
.B2(n_39),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_0),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_108),
.B1(n_74),
.B2(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_49),
.B1(n_64),
.B2(n_23),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_113),
.B1(n_127),
.B2(n_74),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_23),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_97),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_1),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_68),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_86),
.B(n_97),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_68),
.B1(n_73),
.B2(n_88),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_121),
.B1(n_113),
.B2(n_127),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_67),
.A2(n_9),
.B1(n_14),
.B2(n_5),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_125),
.C(n_84),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_87),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_82),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_4),
.C(n_5),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_66),
.A2(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_135),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_152),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_66),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_136),
.C(n_158),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_69),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_125),
.B(n_123),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_104),
.B1(n_108),
.B2(n_109),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_150),
.B1(n_107),
.B2(n_129),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_156),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_93),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_148),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_75),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_147),
.B(n_151),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_102),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_149),
.A2(n_157),
.B1(n_143),
.B2(n_146),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_113),
.A2(n_73),
.B1(n_72),
.B2(n_95),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_83),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_4),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_86),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_155),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_89),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_101),
.B1(n_79),
.B2(n_87),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_107),
.B(n_96),
.C(n_80),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_129),
.A2(n_90),
.B1(n_6),
.B2(n_7),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_121),
.B(n_102),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_180),
.B(n_184),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_164),
.B1(n_168),
.B2(n_158),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_188),
.B1(n_141),
.B2(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_138),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_165),
.B(n_171),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_111),
.B(n_124),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_170),
.B(n_139),
.Y(n_203)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_111),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_120),
.C(n_112),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_187),
.C(n_174),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_137),
.A2(n_90),
.B(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_182),
.Y(n_197)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_115),
.B(n_99),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_112),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_133),
.B(n_144),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_85),
.B1(n_114),
.B2(n_115),
.Y(n_188)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_198),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_204),
.B1(n_207),
.B2(n_179),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_208),
.Y(n_216)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_205),
.C(n_210),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_167),
.A2(n_154),
.B1(n_132),
.B2(n_151),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_162),
.B1(n_173),
.B2(n_175),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_203),
.B(n_172),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_147),
.B1(n_153),
.B2(n_142),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_131),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_181),
.A2(n_142),
.B1(n_8),
.B2(n_10),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_164),
.B(n_169),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_179),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_85),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_114),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_184),
.C(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_7),
.Y(n_213)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_221),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_211),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_176),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_223),
.C(n_233),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_225),
.B(n_209),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_166),
.B(n_171),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_163),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_231),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_183),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_169),
.C(n_170),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_232),
.B(n_196),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_247),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_219),
.A2(n_166),
.B1(n_191),
.B2(n_195),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_241),
.B1(n_168),
.B2(n_220),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_193),
.B1(n_202),
.B2(n_203),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_244),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_177),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_243),
.A2(n_248),
.B(n_249),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_205),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_246),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_204),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_230),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_214),
.C(n_233),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_255),
.C(n_256),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_192),
.B1(n_226),
.B2(n_225),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_254),
.A2(n_180),
.B(n_246),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_216),
.C(n_229),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_209),
.C(n_217),
.Y(n_256)
);

XNOR2x1_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_215),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_258),
.A2(n_262),
.B1(n_249),
.B2(n_241),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_227),
.B(n_224),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_242),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_238),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_231),
.Y(n_262)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_263),
.A2(n_265),
.B1(n_267),
.B2(n_271),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_R g268 ( 
.A(n_258),
.B(n_239),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_270),
.B(n_261),
.Y(n_276)
);

AOI31xp67_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_206),
.A3(n_228),
.B(n_183),
.Y(n_269)
);

OA21x2_ASAP7_75t_SL g280 ( 
.A1(n_269),
.A2(n_10),
.B(n_12),
.Y(n_280)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_259),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_253),
.C(n_265),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_274),
.C(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_257),
.C(n_256),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_268),
.B(n_264),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_259),
.B1(n_254),
.B2(n_161),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_278),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_280),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_283),
.B(n_114),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_267),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_285),
.A2(n_251),
.B(n_13),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_284),
.A2(n_274),
.B(n_278),
.C(n_275),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_287),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_251),
.B(n_13),
.C(n_15),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_288),
.B(n_289),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_281),
.B(n_12),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_290),
.B(n_12),
.Y(n_293)
);


endmodule