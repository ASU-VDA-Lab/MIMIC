module fake_jpeg_27707_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_6),
.B(n_4),
.Y(n_9)
);

HAxp5_ASAP7_75t_SL g10 ( 
.A(n_3),
.B(n_5),
.CON(n_10),
.SN(n_10)
);

INVx4_ASAP7_75t_SL g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_4),
.B(n_1),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_15),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_28)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.C(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_21),
.Y(n_26)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_3),
.B1(n_6),
.B2(n_14),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_12),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_8),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_7),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_11),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_11),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_24)
);

OAI21x1_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_23),
.B(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.C(n_29),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_36),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_26),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.C(n_28),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_28),
.B(n_20),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.B(n_9),
.Y(n_43)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_22),
.A3(n_9),
.B1(n_16),
.B2(n_19),
.C1(n_17),
.C2(n_25),
.Y(n_42)
);


endmodule