module fake_netlist_6_629_n_81 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_81);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_81;

wire n_52;
wire n_46;
wire n_39;
wire n_63;
wire n_73;
wire n_68;
wire n_50;
wire n_49;
wire n_77;
wire n_42;
wire n_54;
wire n_32;
wire n_66;
wire n_78;
wire n_47;
wire n_62;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_38;
wire n_61;
wire n_59;
wire n_76;
wire n_36;
wire n_55;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_40;
wire n_80;
wire n_41;
wire n_71;
wire n_74;
wire n_72;
wire n_60;
wire n_35;
wire n_69;
wire n_79;
wire n_43;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_19),
.Y(n_34)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_3),
.B(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_4),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp67_ASAP7_75t_L g47 ( 
.A(n_11),
.B(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_23),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx11_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

OR2x6_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_7),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_10),
.Y(n_56)
);

O2A1O1Ixp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_14),
.B(n_16),
.C(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_63),
.Y(n_70)
);

NAND2x1p5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_61),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_64),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_73),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_72),
.B1(n_56),
.B2(n_47),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_34),
.B(n_41),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_44),
.A3(n_45),
.B1(n_51),
.B2(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_78),
.B(n_57),
.Y(n_81)
);


endmodule