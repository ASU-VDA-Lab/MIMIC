module fake_jpeg_1164_n_85 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx3_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_36),
.Y(n_39)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_31),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_47),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_52),
.B(n_30),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_0),
.Y(n_63)
);

OAI22x1_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_36),
.B1(n_30),
.B2(n_29),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_65)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NOR3xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_4),
.C(n_5),
.Y(n_68)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_56),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_26),
.B(n_1),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_66),
.B(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_67),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_12),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_3),
.B(n_4),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_70),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_6),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_59),
.B1(n_58),
.B2(n_5),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_78),
.B1(n_73),
.B2(n_8),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_75),
.B(n_72),
.C(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_79),
.B(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_7),
.Y(n_82)
);

AOI322xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.C1(n_17),
.C2(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_19),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_20),
.Y(n_85)
);


endmodule