module fake_jpeg_22024_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx12f_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_7),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_10),
.C(n_11),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_9),
.B1(n_12),
.B2(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_16),
.B(n_15),
.C(n_17),
.Y(n_27)
);

NOR2x1_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_12),
.B1(n_9),
.B2(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_16),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_38),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_20),
.B1(n_16),
.B2(n_1),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_29),
.C(n_28),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_21),
.C(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_39),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_32),
.B1(n_39),
.B2(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

OA21x2_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_39),
.B(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_41),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_47),
.C(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_52),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_47),
.C(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_53),
.Y(n_59)
);

AOI322xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_7),
.A3(n_35),
.B1(n_36),
.B2(n_44),
.C1(n_49),
.C2(n_58),
.Y(n_60)
);


endmodule