module real_jpeg_32876_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_470;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_0),
.A2(n_58),
.B1(n_62),
.B2(n_65),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_0),
.A2(n_65),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_0),
.A2(n_65),
.B1(n_355),
.B2(n_358),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_0),
.A2(n_65),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_89),
.B1(n_94),
.B2(n_95),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_1),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_1),
.A2(n_94),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_1),
.A2(n_94),
.B1(n_395),
.B2(n_399),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_1),
.A2(n_94),
.B1(n_404),
.B2(n_445),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_2),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g279 ( 
.A(n_2),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_2),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_3),
.A2(n_173),
.B1(n_273),
.B2(n_276),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_3),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_6),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_6),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_6),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_7),
.B(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_7),
.A2(n_129),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_7),
.Y(n_326)
);

OAI32xp33_ASAP7_75t_L g361 ( 
.A1(n_7),
.A2(n_112),
.A3(n_362),
.B1(n_365),
.B2(n_366),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_7),
.B(n_25),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_L g459 ( 
.A1(n_7),
.A2(n_136),
.B1(n_444),
.B2(n_460),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_7),
.A2(n_326),
.B1(n_485),
.B2(n_490),
.Y(n_484)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_8),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_8),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_9),
.A2(n_146),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_9),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_11),
.A2(n_79),
.B1(n_83),
.B2(n_86),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_11),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_11),
.A2(n_62),
.B1(n_86),
.B2(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_11),
.A2(n_86),
.B1(n_432),
.B2(n_435),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_11),
.A2(n_86),
.B1(n_449),
.B2(n_452),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_12),
.A2(n_144),
.B1(n_145),
.B2(n_149),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_12),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_12),
.A2(n_144),
.B1(n_211),
.B2(n_215),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_13),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_36)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_13),
.A2(n_41),
.B1(n_238),
.B2(n_241),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_13),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_13),
.A2(n_41),
.B1(n_370),
.B2(n_372),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_15),
.A2(n_178),
.B1(n_179),
.B2(n_184),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_15),
.Y(n_178)
);

AOI22x1_ASAP7_75t_SL g260 ( 
.A1(n_15),
.A2(n_178),
.B1(n_261),
.B2(n_265),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_15),
.A2(n_178),
.B1(n_316),
.B2(n_321),
.Y(n_315)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_16),
.Y(n_194)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_16),
.Y(n_201)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_16),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_17),
.A2(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_17),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_17),
.A2(n_164),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_297),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_244),
.B(n_294),
.Y(n_19)
);

NAND2xp67_ASAP7_75t_SL g296 ( 
.A(n_20),
.B(n_245),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_169),
.C(n_221),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_21),
.B(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_109),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_66),
.B1(n_107),
.B2(n_108),
.Y(n_22)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_36),
.B1(n_48),
.B2(n_57),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_24),
.A2(n_48),
.B1(n_57),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_24),
.A2(n_48),
.B1(n_260),
.B2(n_266),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_24),
.A2(n_48),
.B1(n_224),
.B2(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_24),
.A2(n_48),
.B1(n_306),
.B2(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AO21x2_ASAP7_75t_L g48 ( 
.A1(n_26),
.A2(n_49),
.B(n_53),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_26)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_27),
.Y(n_400)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_29),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_29),
.Y(n_217)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_34),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_34),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_34),
.Y(n_364)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_34),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_40),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_40),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_40),
.Y(n_492)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_46),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_53),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_54),
.Y(n_265)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_60),
.Y(n_227)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_60),
.Y(n_308)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_66),
.B(n_107),
.C(n_109),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_77),
.B1(n_87),
.B2(n_97),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_68),
.A2(n_88),
.B1(n_98),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_68),
.A2(n_78),
.B1(n_98),
.B2(n_252),
.Y(n_251)
);

NOR2x1_ASAP7_75t_L g325 ( 
.A(n_68),
.B(n_326),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_100),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g489 ( 
.A(n_73),
.Y(n_489)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_82),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_82),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_93),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_103),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_133),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_110),
.A2(n_133),
.B1(n_134),
.B2(n_328),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.A3(n_117),
.B1(n_120),
.B2(n_128),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g329 ( 
.A1(n_111),
.A2(n_114),
.A3(n_120),
.B1(n_128),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_143),
.B1(n_154),
.B2(n_158),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_135),
.A2(n_143),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_135),
.A2(n_315),
.B1(n_369),
.B2(n_376),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_135),
.A2(n_470),
.B1(n_471),
.B2(n_472),
.Y(n_469)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_155),
.B1(n_159),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_136),
.A2(n_172),
.B1(n_272),
.B2(n_277),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_136),
.A2(n_418),
.B1(n_420),
.B2(n_421),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_136),
.A2(n_444),
.B1(n_448),
.B2(n_455),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

BUFx2_ASAP7_75t_R g314 ( 
.A(n_137),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_137),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_138),
.Y(n_456)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_138),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_142),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_142),
.Y(n_324)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_148),
.Y(n_320)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_148),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_153),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_153),
.Y(n_466)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_163),
.Y(n_427)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_168),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_170),
.B(n_222),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_171),
.B(n_176),
.Y(n_248)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_173),
.Y(n_422)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_189),
.B1(n_210),
.B2(n_218),
.Y(n_176)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_183),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_184),
.B(n_326),
.Y(n_366)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_188),
.Y(n_288)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_188),
.Y(n_434)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_189),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_189),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_189),
.A2(n_218),
.B1(n_431),
.B2(n_437),
.Y(n_430)
);

AO21x2_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_197),
.B(n_202),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_196),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g415 ( 
.A(n_197),
.Y(n_415)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_208),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_210),
.Y(n_283)
);

BUFx4f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_213),
.Y(n_289)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_217),
.Y(n_388)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.C(n_235),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_223),
.B(n_235),
.Y(n_302)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_228),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI22x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_242),
.B2(n_243),
.Y(n_235)
);

AO22x1_ASAP7_75t_L g353 ( 
.A1(n_236),
.A2(n_237),
.B1(n_290),
.B2(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_243),
.A2(n_385),
.B1(n_393),
.B2(n_394),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2x2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_293),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_268),
.B1(n_269),
.B2(n_292),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_247),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_259),
.B2(n_267),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_280),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_277),
.B(n_326),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_279),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_287),
.Y(n_358)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_290),
.A2(n_354),
.B1(n_393),
.B2(n_482),
.Y(n_481)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_291),
.B(n_326),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_336),
.B(n_507),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_334),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_300),
.B(n_334),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_327),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_301),
.B(n_341),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_327),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_312),
.C(n_325),
.Y(n_304)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_312),
.A2(n_346),
.B(n_347),
.Y(n_351)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_313),
.Y(n_348)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_320),
.Y(n_414)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_320),
.Y(n_447)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_324),
.Y(n_451)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_325),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_350),
.Y(n_349)
);

OAI21xp33_ASAP7_75t_SL g385 ( 
.A1(n_326),
.A2(n_386),
.B(n_389),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_326),
.B(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AOI21x1_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_378),
.B(n_506),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_SL g506 ( 
.A(n_340),
.B(n_342),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_353),
.C(n_359),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_343),
.B(n_501),
.Y(n_500)
);

AOI22x1_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_349),
.B1(n_351),
.B2(n_352),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_345),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_353),
.A2(n_502),
.B(n_503),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_353),
.B(n_360),
.Y(n_503)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_359),
.Y(n_502)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_367),
.Y(n_360)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_361),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_361),
.B(n_368),
.Y(n_497)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_367),
.Y(n_496)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx4f_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_499),
.B(n_505),
.Y(n_378)
);

AOI21x1_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_476),
.B(n_498),
.Y(n_379)
);

OAI21x1_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_440),
.B(n_475),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_416),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_382),
.B(n_416),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_401),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_383),
.A2(n_384),
.B1(n_401),
.B2(n_402),
.Y(n_473)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_389),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_394),
.Y(n_437)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_410),
.B1(n_411),
.B2(n_415),
.Y(n_402)
);

NAND2xp33_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_406),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_428),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_417),
.B(n_430),
.C(n_438),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_421),
.Y(n_471)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_438),
.B2(n_439),
.Y(n_428)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_429),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_430),
.Y(n_439)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_431),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

AOI21x1_ASAP7_75t_SL g440 ( 
.A1(n_441),
.A2(n_468),
.B(n_474),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_458),
.B(n_467),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_457),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_443),
.B(n_457),
.Y(n_467)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx8_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_459),
.B(n_461),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

BUFx2_ASAP7_75t_SL g465 ( 
.A(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_473),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_469),
.B(n_473),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NOR2x1_ASAP7_75t_L g498 ( 
.A(n_477),
.B(n_478),
.Y(n_498)
);

XNOR2x1_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_494),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_480),
.A2(n_481),
.B1(n_483),
.B2(n_493),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_481),
.B(n_493),
.C(n_494),
.Y(n_504)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_483),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_486),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_492),
.Y(n_491)
);

AOI21x1_ASAP7_75t_L g494 ( 
.A1(n_495),
.A2(n_496),
.B(n_497),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_504),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_504),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);


endmodule