module fake_jpeg_29806_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_5),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.Y(n_73)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_1),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_59),
.B1(n_58),
.B2(n_47),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_74),
.B1(n_43),
.B2(n_50),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_76),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_58),
.B1(n_42),
.B2(n_55),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_2),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_78),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_75),
.B(n_69),
.C(n_49),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_95),
.B(n_3),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_46),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_86),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_52),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_88),
.Y(n_101)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_68),
.B1(n_55),
.B2(n_42),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_2),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_80),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_44),
.A3(n_21),
.B1(n_22),
.B2(n_39),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_19),
.B1(n_37),
.B2(n_35),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_105),
.B1(n_14),
.B2(n_17),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_102),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_7),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_7),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_8),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_118),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_12),
.B(n_13),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_125),
.B(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_18),
.C(n_20),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_24),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_108),
.B1(n_26),
.B2(n_29),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_117),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_101),
.B(n_111),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_116),
.C(n_126),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_134),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_138),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_137),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_135),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_139),
.C(n_123),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_115),
.C(n_122),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_136),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_133),
.B1(n_129),
.B2(n_120),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_121),
.C(n_33),
.Y(n_148)
);


endmodule