module fake_jpeg_26517_n_102 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_0),
.C(n_1),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_0),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_59),
.B1(n_62),
.B2(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_54),
.B(n_53),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_29),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_36),
.B1(n_35),
.B2(n_37),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_30),
.B1(n_38),
.B2(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_5),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_30),
.B1(n_19),
.B2(n_22),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_17),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_1),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_73),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_76),
.Y(n_82)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_7),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_8),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_10),
.B(n_11),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_70),
.B(n_73),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_90),
.B(n_91),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_92),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_95),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_82),
.C(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_94),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_83),
.B1(n_79),
.B2(n_85),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_87),
.B(n_23),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_14),
.Y(n_102)
);


endmodule