module fake_jpeg_2124_n_185 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_63),
.Y(n_69)
);

BUFx12f_ASAP7_75t_SL g62 ( 
.A(n_55),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_60),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_50),
.B1(n_46),
.B2(n_57),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_74),
.B1(n_66),
.B2(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_44),
.Y(n_82)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_44),
.B1(n_56),
.B2(n_58),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_52),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_62),
.B(n_52),
.C(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_88),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_90),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_65),
.B1(n_64),
.B2(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_6),
.Y(n_111)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_72),
.B(n_47),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_0),
.C(n_1),
.Y(n_101)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_66),
.B1(n_64),
.B2(n_59),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_75),
.B1(n_47),
.B2(n_2),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_13),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_76),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_100),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_20),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_112),
.C(n_109),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_75),
.B1(n_47),
.B2(n_21),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_101),
.Y(n_117)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_10),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_35),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_85),
.C(n_79),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_122),
.C(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_11),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_119),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_12),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_87),
.C(n_28),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_27),
.C(n_42),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_14),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_14),
.Y(n_126)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_15),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_131),
.B(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_15),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_16),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_99),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_134),
.C(n_146),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_95),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_104),
.B(n_17),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_138),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_17),
.B(n_18),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_19),
.A3(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_143),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_150),
.B1(n_38),
.B2(n_43),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_33),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_123),
.B1(n_39),
.B2(n_40),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_156),
.B1(n_157),
.B2(n_159),
.Y(n_162)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_149),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_147),
.C(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_133),
.C(n_146),
.Y(n_164)
);

XOR2x2_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_153),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_169),
.A2(n_162),
.B1(n_144),
.B2(n_155),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_161),
.B(n_140),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_161),
.C(n_168),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_173),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_172),
.C(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_143),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_169),
.B(n_175),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_160),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_136),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_160),
.Y(n_185)
);


endmodule