module real_jpeg_14325_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_273, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_273;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_3),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_3),
.A2(n_64),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_3),
.B(n_141),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_149),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_3),
.A2(n_43),
.B(n_48),
.C(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_3),
.B(n_109),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_3),
.B(n_32),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_3),
.B(n_53),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_3),
.A2(n_62),
.B(n_73),
.C(n_247),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_4),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_4),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_68),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_29),
.B1(n_35),
.B2(n_68),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_52),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_6),
.A2(n_52),
.B1(n_59),
.B2(n_62),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_7),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_7),
.A2(n_59),
.B1(n_62),
.B2(n_102),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_102),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_7),
.A2(n_29),
.B1(n_35),
.B2(n_102),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_8),
.A2(n_59),
.B1(n_62),
.B2(n_70),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_70),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_8),
.A2(n_29),
.B1(n_35),
.B2(n_70),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_12),
.A2(n_59),
.B1(n_62),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_79),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_79),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_13),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_13),
.A2(n_59),
.B1(n_62),
.B2(n_138),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_138),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_138),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_14),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_15),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_15),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_111)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_17),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_17),
.A2(n_45),
.B1(n_59),
.B2(n_62),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_17),
.A2(n_29),
.B1(n_35),
.B2(n_45),
.Y(n_145)
);

HAxp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_125),
.CON(n_18),
.SN(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_103),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_103),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_81),
.C(n_87),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_23),
.B(n_81),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_24),
.B(n_56),
.C(n_71),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_26),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_162)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_28),
.A2(n_32),
.B(n_37),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_28),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_28),
.A2(n_32),
.B1(n_93),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_28),
.A2(n_32),
.B1(n_145),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_28),
.A2(n_32),
.B1(n_181),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_28),
.A2(n_32),
.B1(n_192),
.B2(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_28),
.A2(n_32),
.B1(n_149),
.B2(n_232),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_28),
.A2(n_32),
.B1(n_225),
.B2(n_232),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_29),
.B(n_234),
.Y(n_233)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_31),
.A2(n_34),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_31),
.A2(n_91),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_35),
.A2(n_49),
.B(n_149),
.Y(n_213)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_42),
.A2(n_50),
.B1(n_95),
.B2(n_97),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_44),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_43),
.B(n_76),
.Y(n_190)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_44),
.A2(n_62),
.A3(n_75),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_46),
.A2(n_53),
.B1(n_85),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_46),
.A2(n_53),
.B1(n_96),
.B2(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_46),
.A2(n_53),
.B1(n_154),
.B2(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_46),
.A2(n_53),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_46),
.A2(n_53),
.B1(n_211),
.B2(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_50),
.A2(n_97),
.B1(n_184),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_57),
.A2(n_58),
.B1(n_137),
.B2(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_62),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_59),
.A2(n_61),
.A3(n_64),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_59),
.B(n_149),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_60),
.B(n_62),
.Y(n_147)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_65),
.B(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_77),
.B1(n_78),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_72),
.A2(n_77),
.B1(n_133),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_109),
.B1(n_132),
.B2(n_134),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_73),
.A2(n_109),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_77),
.A2(n_176),
.B(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_83),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_87),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.C(n_100),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_88),
.A2(n_89),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_90),
.B(n_94),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_100),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_123),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_113),
.B1(n_114),
.B2(n_122),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_110),
.B(n_112),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_110),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_121),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_266),
.B(n_270),
.Y(n_125)
);

OAI221xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_169),
.B1(n_264),
.B2(n_265),
.C(n_273),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_160),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_128),
.B(n_160),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_150),
.C(n_151),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_129),
.B(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_142),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_135),
.C(n_142),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_150),
.B(n_151),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_157),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_162),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_162),
.B(n_167),
.C(n_168),
.Y(n_267)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_260),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_203),
.B(n_259),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_193),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_172),
.B(n_193),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_182),
.C(n_185),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_173),
.B(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_179),
.C(n_180),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_182),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_189),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_191),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_198),
.B2(n_202),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_194),
.B(n_199),
.C(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_253),
.B(n_258),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_241),
.B(n_252),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_221),
.B(n_240),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_217),
.C(n_219),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_220),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_229),
.B(n_239),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_223),
.B(n_227),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_235),
.B(n_238),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_243),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_248),
.C(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_262),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);


endmodule