module fake_jpeg_1468_n_535 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_535);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_535;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_58),
.Y(n_202)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_60),
.Y(n_187)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_64),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_69),
.B(n_77),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_72),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_76),
.Y(n_208)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_18),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_95),
.Y(n_152)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_85),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_24),
.B(n_16),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_100),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_24),
.Y(n_95)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_96),
.Y(n_195)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_98),
.B(n_105),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_99),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_54),
.B(n_15),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_102),
.Y(n_207)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_56),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_109),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_23),
.B(n_15),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_2),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_56),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_164)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_25),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_114),
.Y(n_170)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_25),
.Y(n_114)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_121),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_56),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_117),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_57),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_28),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_118),
.B(n_120),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx5_ASAP7_75t_SL g134 ( 
.A(n_119),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_122),
.B(n_123),
.Y(n_201)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_29),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_37),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_29),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_7),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_85),
.A2(n_50),
.B1(n_22),
.B2(n_47),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_126),
.A2(n_133),
.B1(n_143),
.B2(n_145),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_68),
.A2(n_31),
.B(n_53),
.C(n_44),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_127),
.A2(n_162),
.B(n_129),
.C(n_152),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_108),
.B1(n_70),
.B2(n_73),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_128),
.A2(n_131),
.B1(n_144),
.B2(n_147),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_50),
.B1(n_22),
.B2(n_47),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_85),
.A2(n_50),
.B1(n_22),
.B2(n_46),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_27),
.B1(n_53),
.B2(n_44),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_106),
.A2(n_55),
.B1(n_31),
.B2(n_36),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_60),
.A2(n_33),
.B1(n_48),
.B2(n_46),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_55),
.B1(n_36),
.B2(n_42),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_60),
.A2(n_48),
.B1(n_37),
.B2(n_33),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_150),
.A2(n_160),
.B1(n_161),
.B2(n_174),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_156),
.B(n_193),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_89),
.A2(n_41),
.B1(n_39),
.B2(n_42),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_41),
.B1(n_39),
.B2(n_5),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_124),
.B(n_15),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_163),
.B(n_196),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_164),
.A2(n_199),
.B1(n_204),
.B2(n_209),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_186),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_183),
.B(n_142),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_80),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_86),
.A2(n_99),
.B1(n_102),
.B2(n_104),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_175),
.A2(n_177),
.B1(n_190),
.B2(n_198),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_92),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_90),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_189),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_123),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_62),
.B(n_76),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_200),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_82),
.B(n_8),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_121),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_122),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_113),
.B(n_14),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_65),
.A2(n_14),
.B1(n_72),
.B2(n_87),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_203),
.A2(n_154),
.B1(n_185),
.B2(n_209),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_114),
.A2(n_115),
.B1(n_97),
.B2(n_58),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_58),
.A2(n_51),
.B1(n_30),
.B2(n_43),
.Y(n_209)
);

INVx4_ASAP7_75t_SL g210 ( 
.A(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_210),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_127),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_211),
.B(n_216),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_212),
.Y(n_315)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_213),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_214),
.B(n_225),
.Y(n_307)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

INVx4_ASAP7_75t_SL g290 ( 
.A(n_215),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_141),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_201),
.A2(n_199),
.B1(n_128),
.B2(n_137),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_219),
.A2(n_239),
.B1(n_233),
.B2(n_229),
.Y(n_306)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_220),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_221),
.B(n_230),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_224),
.B(n_237),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_170),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_181),
.A2(n_176),
.B(n_177),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_226),
.A2(n_271),
.B(n_272),
.Y(n_332)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_146),
.Y(n_227)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

BUFx8_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_184),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_229),
.B(n_245),
.Y(n_318)
);

NOR2x1_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_170),
.Y(n_230)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_139),
.B(n_155),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_234),
.B(n_260),
.Y(n_328)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_202),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_202),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_238),
.B(n_242),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_140),
.A2(n_149),
.B1(n_166),
.B2(n_148),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g241 ( 
.A(n_153),
.Y(n_241)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_132),
.B(n_197),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_130),
.Y(n_243)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_243),
.Y(n_319)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_187),
.Y(n_244)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_159),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_151),
.B(n_157),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_246),
.A2(n_249),
.B(n_224),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_247),
.Y(n_281)
);

NAND2x1_ASAP7_75t_SL g249 ( 
.A(n_154),
.B(n_151),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_250),
.A2(n_276),
.B1(n_272),
.B2(n_271),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_132),
.B(n_197),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_253),
.Y(n_301)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_159),
.B(n_208),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_167),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_254),
.B(n_259),
.Y(n_302)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_168),
.Y(n_255)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_256),
.Y(n_291)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_257),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_208),
.B(n_157),
.C(n_136),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_271),
.C(n_272),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_136),
.B(n_153),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_149),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_188),
.Y(n_261)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_204),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_262),
.B(n_263),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_145),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_150),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_265),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_193),
.B(n_207),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_266),
.B(n_270),
.Y(n_323)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_206),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_267),
.B(n_268),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_140),
.B(n_205),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_167),
.B(n_205),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_269),
.B(n_273),
.Y(n_331)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_135),
.B(n_182),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_135),
.B(n_182),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_180),
.B(n_126),
.Y(n_273)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_180),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_275),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_179),
.A2(n_195),
.B1(n_133),
.B2(n_134),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_195),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_279),
.Y(n_325)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_146),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_278),
.A2(n_241),
.B1(n_215),
.B2(n_246),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_179),
.B(n_146),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_264),
.B(n_226),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_284),
.A2(n_297),
.B(n_326),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_286),
.Y(n_352)
);

AOI32xp33_ASAP7_75t_L g288 ( 
.A1(n_211),
.A2(n_235),
.A3(n_225),
.B1(n_230),
.B2(n_273),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_288),
.B(n_330),
.Y(n_355)
);

O2A1O1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_236),
.A2(n_223),
.B(n_262),
.C(n_231),
.Y(n_297)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_227),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_298),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_217),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_305),
.B(n_321),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_306),
.A2(n_308),
.B1(n_311),
.B2(n_267),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_219),
.A2(n_274),
.B1(n_214),
.B2(n_265),
.Y(n_308)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_210),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_274),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_248),
.A2(n_260),
.B1(n_240),
.B2(n_234),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_316),
.A2(n_245),
.B1(n_244),
.B2(n_213),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_317),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_246),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_322),
.A2(n_325),
.B1(n_303),
.B2(n_300),
.Y(n_366)
);

O2A1O1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_246),
.A2(n_249),
.B(n_258),
.C(n_261),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_216),
.B(n_222),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_278),
.Y(n_345)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_270),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_343),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_311),
.A2(n_275),
.B1(n_232),
.B2(n_252),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_335),
.A2(n_336),
.B1(n_340),
.B2(n_360),
.Y(n_381)
);

NOR2x1_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_257),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_337),
.B(n_338),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_324),
.B(n_256),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_255),
.C(n_220),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_346),
.C(n_299),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_308),
.A2(n_243),
.B1(n_218),
.B2(n_239),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_341),
.Y(n_402)
);

AO21x1_ASAP7_75t_L g398 ( 
.A1(n_342),
.A2(n_345),
.B(n_361),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_277),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_228),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_329),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_350),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_316),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_301),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_362),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_314),
.A2(n_286),
.B(n_312),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_353),
.A2(n_296),
.B(n_299),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_305),
.B(n_302),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_354),
.B(n_367),
.Y(n_373)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_356),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_293),
.Y(n_358)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_358),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_318),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_SL g374 ( 
.A(n_359),
.B(n_291),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_306),
.A2(n_297),
.B1(n_284),
.B2(n_280),
.Y(n_360)
);

AO21x2_ASAP7_75t_L g361 ( 
.A1(n_322),
.A2(n_280),
.B(n_326),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_288),
.B(n_304),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_332),
.A2(n_295),
.B1(n_304),
.B2(n_318),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_363),
.A2(n_320),
.B1(n_327),
.B2(n_296),
.Y(n_386)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_290),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_366),
.A2(n_282),
.B1(n_291),
.B2(n_290),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_285),
.B(n_281),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_285),
.B(n_315),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_320),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_318),
.A2(n_303),
.B1(n_293),
.B2(n_282),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_369),
.A2(n_352),
.B1(n_357),
.B2(n_359),
.Y(n_392)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_283),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_289),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_371),
.B(n_372),
.Y(n_401)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_289),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_374),
.A2(n_383),
.B(n_392),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_375),
.A2(n_347),
.B1(n_345),
.B2(n_359),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_348),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_382),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_330),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_388),
.C(n_399),
.Y(n_413)
);

XOR2x2_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_296),
.Y(n_378)
);

XOR2x1_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_345),
.Y(n_416)
);

NAND3xp33_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_389),
.C(n_400),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_364),
.A2(n_290),
.B(n_296),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_386),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_313),
.C(n_327),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_313),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_350),
.A2(n_319),
.B1(n_294),
.B2(n_298),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_394),
.A2(n_395),
.B1(n_396),
.B2(n_344),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_361),
.A2(n_319),
.B1(n_294),
.B2(n_287),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_361),
.A2(n_294),
.B1(n_287),
.B2(n_292),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_292),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_310),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_340),
.A2(n_361),
.B1(n_364),
.B2(n_335),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_403),
.A2(n_356),
.B1(n_370),
.B2(n_341),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_406),
.A2(n_415),
.B1(n_419),
.B2(n_423),
.Y(n_457)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_405),
.Y(n_410)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_410),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_373),
.B(n_338),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_411),
.B(n_426),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_346),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_417),
.C(n_421),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_343),
.Y(n_414)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_403),
.A2(n_361),
.B1(n_352),
.B2(n_357),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_416),
.A2(n_425),
.B(n_430),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_339),
.C(n_353),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_420),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_337),
.C(n_369),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_333),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_432),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_381),
.A2(n_342),
.B1(n_372),
.B2(n_371),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_424),
.A2(n_429),
.B1(n_395),
.B2(n_396),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_375),
.A2(n_358),
.B1(n_365),
.B2(n_348),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_390),
.B(n_358),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_401),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_427),
.B(n_433),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_378),
.C(n_379),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_382),
.C(n_393),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_381),
.A2(n_392),
.B1(n_379),
.B2(n_398),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_383),
.A2(n_382),
.B(n_374),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_387),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_431),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_404),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_376),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_434),
.A2(n_415),
.B1(n_423),
.B2(n_406),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_378),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_443),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_422),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_437),
.B(n_450),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_427),
.B(n_393),
.Y(n_440)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_425),
.Y(n_442)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_386),
.Y(n_443)
);

XNOR2x2_ASAP7_75t_SL g444 ( 
.A(n_414),
.B(n_432),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_444),
.B(n_448),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_408),
.B(n_391),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_445),
.B(n_455),
.Y(n_464)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_429),
.Y(n_446)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_446),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_387),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_424),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_398),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_407),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_421),
.B(n_391),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_458),
.C(n_413),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_409),
.B(n_402),
.C(n_397),
.Y(n_458)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_460),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_440),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_465),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_439),
.B(n_437),
.Y(n_463)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_463),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_407),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_452),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_468),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_439),
.B(n_419),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_454),
.A2(n_430),
.B(n_418),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_469),
.A2(n_436),
.B(n_441),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_435),
.B(n_410),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_478),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_472),
.A2(n_447),
.B1(n_449),
.B2(n_441),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_474),
.B(n_451),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_454),
.A2(n_418),
.B(n_398),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_475),
.A2(n_457),
.B(n_453),
.Y(n_481)
);

AOI322xp5_ASAP7_75t_SL g477 ( 
.A1(n_435),
.A2(n_416),
.A3(n_428),
.B1(n_409),
.B2(n_431),
.C1(n_394),
.C2(n_402),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_477),
.A2(n_456),
.B1(n_453),
.B2(n_443),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_438),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_476),
.A2(n_446),
.B1(n_434),
.B2(n_449),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_479),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_480),
.B(n_462),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_481),
.A2(n_489),
.B(n_475),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_474),
.B(n_458),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_480),
.Y(n_494)
);

NOR2x1_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_462),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_485),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_448),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_487),
.B(n_493),
.C(n_469),
.Y(n_502)
);

A2O1A1Ixp33_ASAP7_75t_L g492 ( 
.A1(n_476),
.A2(n_444),
.B(n_451),
.C(n_438),
.Y(n_492)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_492),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_397),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_496),
.Y(n_510)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_486),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_498),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_490),
.B(n_466),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_499),
.A2(n_505),
.B(n_491),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_485),
.A2(n_463),
.B1(n_459),
.B2(n_468),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_501),
.B(n_503),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_502),
.B(n_487),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_464),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_504),
.A2(n_482),
.B(n_464),
.Y(n_507)
);

BUFx24_ASAP7_75t_SL g506 ( 
.A(n_499),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_509),
.Y(n_519)
);

NOR3xp33_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_470),
.C(n_505),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_483),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_514),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_489),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_495),
.B(n_500),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_495),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_501),
.Y(n_518)
);

AOI322xp5_ASAP7_75t_L g526 ( 
.A1(n_516),
.A2(n_465),
.A3(n_486),
.B1(n_488),
.B2(n_477),
.C1(n_467),
.C2(n_498),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_492),
.C(n_481),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_518),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_496),
.C(n_497),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_522),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_479),
.C(n_493),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_523),
.A2(n_467),
.B(n_472),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_526),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_518),
.Y(n_531)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_520),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_519),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_530),
.B(n_531),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_524),
.C(n_525),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_478),
.B(n_471),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_532),
.Y(n_535)
);


endmodule