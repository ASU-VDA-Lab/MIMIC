module fake_jpeg_9465_n_107 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_24),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_39),
.B1(n_12),
.B2(n_1),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_22),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_16),
.C(n_13),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_18),
.B1(n_14),
.B2(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_50),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_32),
.B1(n_21),
.B2(n_18),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_55),
.B1(n_58),
.B2(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_43),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_59),
.B(n_61),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_31),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_10),
.C(n_11),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_25),
.B1(n_20),
.B2(n_13),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_20),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_15),
.B(n_23),
.C(n_2),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_41),
.B1(n_29),
.B2(n_26),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_44),
.B(n_29),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_55),
.C(n_50),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_29),
.B(n_26),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_51),
.B(n_54),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_60),
.B(n_61),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_57),
.Y(n_78)
);

AOI221xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_81),
.B1(n_71),
.B2(n_70),
.C(n_59),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_49),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_82),
.C(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_90),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_80),
.C(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_42),
.B1(n_5),
.B2(n_7),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_93),
.B(n_85),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_73),
.B1(n_66),
.B2(n_68),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_42),
.B1(n_5),
.B2(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_89),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_92),
.B(n_93),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_99),
.A3(n_8),
.B1(n_9),
.B2(n_0),
.C1(n_4),
.C2(n_26),
.Y(n_102)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_88),
.C(n_44),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_9),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_4),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.C(n_101),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_68),
.B(n_53),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_4),
.Y(n_107)
);


endmodule