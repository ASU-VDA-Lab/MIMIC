module real_jpeg_8178_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_1),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_2),
.A2(n_34),
.B1(n_38),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_2),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_34),
.B1(n_38),
.B2(n_56),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_10),
.A2(n_34),
.B1(n_38),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_43),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_43),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_11),
.A2(n_34),
.B1(n_38),
.B2(n_48),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_23),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_12),
.A2(n_22),
.B(n_23),
.C(n_59),
.D(n_61),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_12),
.B(n_73),
.Y(n_72)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_12),
.A2(n_26),
.B(n_50),
.C(n_84),
.D(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_12),
.B(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_12),
.B(n_60),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_12),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_12),
.A2(n_109),
.B(n_110),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_89),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_88),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_64),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_17),
.B(n_64),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_45),
.C(n_58),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_18),
.A2(n_19),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_31),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_24),
.A2(n_28),
.B(n_30),
.C(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_60)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_51),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_39),
.B(n_41),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_33),
.A2(n_40),
.B1(n_44),
.B2(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_38),
.B1(n_51),
.B2(n_52),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_34),
.A2(n_53),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_38),
.B(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_38),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_39),
.A2(n_41),
.B(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_39),
.B(n_122),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_40),
.B(n_42),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_40),
.A2(n_44),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_45),
.A2(n_46),
.B1(n_58),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_47),
.A2(n_57),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_55),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_50),
.B(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_57),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_68),
.B(n_69),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_80),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_79),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_85),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_131),
.B(n_137),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_111),
.B(n_130),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_92),
.B(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_95),
.B1(n_96),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_107),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_104),
.C(n_107),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B(n_110),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_119),
.B(n_129),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_113),
.B(n_117),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_124),
.B(n_128),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);


endmodule