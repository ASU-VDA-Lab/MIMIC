module real_jpeg_4079_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_1),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_1),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_1),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_1),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_1),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_1),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_1),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_1),
.B(n_371),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_2),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_2),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_2),
.B(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_2),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_2),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_2),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_2),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_2),
.B(n_392),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_3),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_96),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_4),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_4),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_4),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_4),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_4),
.B(n_408),
.Y(n_407)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_6),
.Y(n_191)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_6),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_6),
.Y(n_392)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_7),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g224 ( 
.A(n_7),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_8),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_8),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_8),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_8),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_8),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_8),
.B(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_10),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_10),
.Y(n_219)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_10),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_11),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_11),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_12),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_12),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_12),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_12),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_12),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_13),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_14),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_14),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_14),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_14),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_14),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_15),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_15),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_15),
.B(n_96),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_15),
.B(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_15),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_15),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_15),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_15),
.B(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_172),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_170),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_145),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_19),
.B(n_145),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_101),
.C(n_112),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g468 ( 
.A(n_20),
.B(n_101),
.CI(n_112),
.CON(n_468),
.SN(n_468)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_58),
.B1(n_99),
.B2(n_100),
.Y(n_20)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_22),
.B(n_40),
.C(n_100),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.C(n_35),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_23),
.B(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.C(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_47),
.C(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_24),
.A2(n_29),
.B1(n_69),
.B2(n_126),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_24),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_24),
.A2(n_121),
.B1(n_126),
.B2(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_24),
.A2(n_126),
.B1(n_377),
.B2(n_378),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_67),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g133 ( 
.A(n_25),
.B(n_134),
.Y(n_133)
);

OR2x2_ASAP7_75t_SL g163 ( 
.A(n_25),
.B(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_27),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_27),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_29),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_29),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_29),
.B(n_60),
.C(n_66),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_29),
.B(n_315),
.C(n_319),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_29),
.A2(n_69),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g426 ( 
.A(n_32),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_33),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_35),
.A2(n_36),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_35),
.A2(n_36),
.B1(n_139),
.B2(n_140),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_36),
.B(n_129),
.C(n_139),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_38),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_38),
.Y(n_275)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_39),
.Y(n_195)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_39),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_57),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_41),
.B(n_47),
.C(n_52),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_52),
.B2(n_56),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_46),
.A2(n_47),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_50),
.Y(n_241)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_70),
.C(n_84),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_59),
.B(n_350),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_65),
.A2(n_66),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_65),
.B(n_104),
.C(n_106),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_65),
.A2(n_66),
.B1(n_121),
.B2(n_290),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_66),
.B(n_121),
.C(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_70),
.B(n_84),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.C(n_79),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_71),
.A2(n_117),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_71),
.B(n_106),
.C(n_239),
.Y(n_265)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_75),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_79),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_78),
.Y(n_380)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_82),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_82),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_82),
.Y(n_394)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_83),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_95),
.B2(n_98),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_86)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_94),
.C(n_95),
.Y(n_111)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_88),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_89),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_89),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_89),
.B(n_268),
.C(n_272),
.Y(n_282)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_97),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_108),
.B2(n_109),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_110),
.C(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_106),
.A2(n_107),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_106),
.A2(n_107),
.B1(n_238),
.B2(n_243),
.Y(n_237)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_128),
.C(n_142),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_113),
.A2(n_114),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_123),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_120),
.Y(n_335)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_121),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_122),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_123),
.B(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_126),
.B(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_128),
.B(n_142),
.Y(n_352)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_130),
.B(n_342),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_136),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_132),
.B(n_137),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_133),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_133),
.Y(n_284)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g470 ( 
.A(n_145),
.Y(n_470)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_147),
.CI(n_148),
.CON(n_145),
.SN(n_145)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_158),
.B2(n_169),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_157),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_156),
.Y(n_235)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_163),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_163),
.B(n_213),
.C(n_218),
.Y(n_296)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_164),
.Y(n_321)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_466),
.B(n_469),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AO21x2_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_345),
.B(n_354),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_329),
.B(n_344),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_305),
.B(n_328),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_177),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_277),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_178),
.B(n_277),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_236),
.C(n_263),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_179),
.B(n_327),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_179),
.Y(n_472)
);

FAx1_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_210),
.CI(n_221),
.CON(n_179),
.SN(n_179)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_180),
.B(n_210),
.C(n_221),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_196),
.C(n_202),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_181),
.B(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_192),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_183),
.B(n_188),
.C(n_192),
.Y(n_276)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_186),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_187),
.Y(n_401)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_196),
.A2(n_202),
.B1(n_203),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_196),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_197),
.B(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_322)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_207),
.Y(n_418)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_212)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_213),
.A2(n_220),
.B1(n_249),
.B2(n_250),
.Y(n_386)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_223),
.B(n_225),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_222),
.B(n_229),
.C(n_232),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_227),
.B(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_233),
.B(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_233),
.B(n_383),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_233),
.B(n_416),
.Y(n_415)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_236),
.B(n_263),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_244),
.C(n_246),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_237),
.A2(n_244),
.B1(n_245),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_246),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.C(n_258),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_247),
.A2(n_248),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_259),
.Y(n_454)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_276),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_266),
.C(n_276),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_280),
.C(n_304),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_291),
.B1(n_303),
.B2(n_304),
.Y(n_279)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_287),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_282),
.B(n_283),
.C(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_301),
.C(n_340),
.Y(n_339)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_326),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_306),
.B(n_326),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_311),
.C(n_323),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_307),
.A2(n_308),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_311),
.B(n_323),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.C(n_322),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_312),
.B(n_446),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_314),
.B(n_322),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_315),
.A2(n_316),
.B1(n_319),
.B2(n_320),
.Y(n_374)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_330),
.B(n_345),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_332),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_346),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_332),
.B(n_346),
.Y(n_465)
);

FAx1_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_336),
.CI(n_343),
.CON(n_332),
.SN(n_332)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_339),
.C(n_341),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_347),
.B(n_349),
.C(n_351),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

OAI31xp33_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_462),
.A3(n_463),
.B(n_465),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_456),
.B(n_461),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_441),
.B(n_455),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_396),
.B(n_440),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_387),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_359),
.B(n_387),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_375),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_372),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_361),
.B(n_372),
.C(n_375),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.C(n_369),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_362),
.A2(n_363),
.B1(n_365),
.B2(n_366),
.Y(n_389)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_369),
.B(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_381),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_376),
.B(n_450),
.C(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_386),
.Y(n_381)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_386),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.C(n_395),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_388),
.B(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_390),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_390),
.A2(n_395),
.B1(n_432),
.B2(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_391),
.Y(n_430)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_392),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_393),
.Y(n_431)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_395),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_434),
.B(n_439),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_420),
.B(n_433),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_405),
.B(n_419),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_415),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_415),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_410),
.B(n_414),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_410),
.Y(n_414)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_414),
.A2(n_422),
.B1(n_427),
.B2(n_428),
.Y(n_421)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_414),
.Y(n_427)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx8_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_429),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_429),
.Y(n_433)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_422),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_423),
.A2(n_424),
.B(n_427),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_430),
.A2(n_431),
.B(n_432),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_435),
.B(n_436),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_443),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_447),
.B2(n_448),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_449),
.C(n_452),
.Y(n_457)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_457),
.B(n_458),
.Y(n_461)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_459),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_467),
.B(n_468),
.Y(n_469)
);

BUFx24_ASAP7_75t_SL g471 ( 
.A(n_468),
.Y(n_471)
);


endmodule