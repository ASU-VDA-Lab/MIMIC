module fake_jpeg_2985_n_203 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_203);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_5),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_1),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_73),
.Y(n_89)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_79),
.Y(n_90)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_0),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_57),
.B1(n_61),
.B2(n_66),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_89),
.B1(n_84),
.B2(n_80),
.Y(n_94)
);

BUFx12f_ASAP7_75t_SL g84 ( 
.A(n_73),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_88),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_57),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_55),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_64),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_72),
.B1(n_90),
.B2(n_80),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_3),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_74),
.B(n_66),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_70),
.C(n_49),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_72),
.B1(n_55),
.B2(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_61),
.B1(n_57),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_109),
.B1(n_59),
.B2(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_26),
.Y(n_116)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_110),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_50),
.B(n_54),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

OR2x4_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_50),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_60),
.B1(n_59),
.B2(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_67),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_115),
.B1(n_125),
.B2(n_117),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_70),
.B1(n_49),
.B2(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_3),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_127),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_70),
.B1(n_49),
.B2(n_63),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_5),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_6),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_105),
.B1(n_107),
.B2(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_140),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_27),
.B(n_45),
.C(n_44),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_149),
.B(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_143),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_24),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_122),
.B1(n_120),
.B2(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_146),
.B(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_15),
.B(n_18),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_12),
.B(n_14),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_15),
.B(n_16),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_171),
.B(n_138),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_31),
.C(n_17),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_163),
.Y(n_179)
);

OR2x6_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_145),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_32),
.Y(n_164)
);

OAI322xp33_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_139),
.A3(n_143),
.B1(n_25),
.B2(n_29),
.C1(n_30),
.C2(n_33),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_139),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

NAND2x1p5_ASAP7_75t_R g171 ( 
.A(n_142),
.B(n_21),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_172),
.Y(n_174)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_180),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

INVxp33_ASAP7_75t_SL g182 ( 
.A(n_171),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_182),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_137),
.B(n_23),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_160),
.B(n_165),
.C(n_167),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_183),
.B1(n_163),
.B2(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_164),
.C(n_161),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_191),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_168),
.A3(n_163),
.B1(n_173),
.B2(n_159),
.C1(n_172),
.C2(n_42),
.Y(n_191)
);

AOI211xp5_ASAP7_75t_L g197 ( 
.A1(n_192),
.A2(n_194),
.B(n_185),
.C(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_176),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_189),
.C(n_184),
.Y(n_196)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

AOI211xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_197),
.B(n_198),
.C(n_195),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_193),
.B(n_188),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_22),
.B(n_34),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_37),
.Y(n_203)
);


endmodule