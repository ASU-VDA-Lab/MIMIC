module real_jpeg_29206_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_50;
wire n_29;
wire n_55;
wire n_49;
wire n_52;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_47;
wire n_14;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_53;
wire n_18;
wire n_22;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_48;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_0),
.A2(n_17),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B1(n_25),
.B2(n_26),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

NOR3xp33_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_8),
.C(n_16),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_2),
.A2(n_16),
.B(n_19),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_2),
.A2(n_6),
.B(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_2),
.B(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_2),
.B(n_48),
.Y(n_47)
);

OAI31xp33_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_3),
.A3(n_19),
.B(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_6),
.A2(n_18),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_7),
.B(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_20),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

OAI31xp33_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_30),
.A3(n_33),
.B(n_37),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_27),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_15),
.A2(n_25),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_44),
.C(n_51),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);


endmodule