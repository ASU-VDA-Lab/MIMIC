module real_aes_8713_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g429 ( .A(n_0), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_1), .A2(n_115), .B(n_118), .C(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g181 ( .A(n_2), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_3), .A2(n_110), .B(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_4), .B(n_191), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g192 ( .A1(n_5), .A2(n_110), .B(n_193), .Y(n_192) );
AND2x6_ASAP7_75t_L g115 ( .A(n_6), .B(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_7), .A2(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_8), .B(n_41), .Y(n_430) );
INVx1_ASAP7_75t_L g443 ( .A(n_9), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_10), .B(n_151), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_11), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g198 ( .A(n_12), .Y(n_198) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_13), .A2(n_19), .B1(n_101), .B2(n_701), .C1(n_702), .C2(n_706), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_13), .Y(n_701) );
INVx1_ASAP7_75t_L g136 ( .A(n_14), .Y(n_136) );
INVx1_ASAP7_75t_L g169 ( .A(n_15), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_16), .A2(n_124), .B(n_170), .C(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_17), .B(n_191), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_18), .B(n_126), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_20), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_21), .B(n_544), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_22), .A2(n_150), .B(n_184), .C(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_23), .B(n_191), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_24), .B(n_151), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g165 ( .A1(n_25), .A2(n_166), .B(n_168), .C(n_170), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_26), .B(n_151), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_27), .Y(n_493) );
INVx1_ASAP7_75t_L g482 ( .A(n_28), .Y(n_482) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_29), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_30), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_31), .B(n_151), .Y(n_182) );
INVx1_ASAP7_75t_L g540 ( .A(n_32), .Y(n_540) );
INVx1_ASAP7_75t_L g208 ( .A(n_33), .Y(n_208) );
INVx2_ASAP7_75t_L g113 ( .A(n_34), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_35), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_36), .A2(n_150), .B(n_199), .C(n_506), .Y(n_505) );
INVxp67_ASAP7_75t_L g541 ( .A(n_37), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g117 ( .A1(n_38), .A2(n_115), .B(n_118), .C(n_121), .Y(n_117) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_39), .A2(n_118), .B(n_481), .C(n_486), .Y(n_480) );
CKINVDCx14_ASAP7_75t_R g504 ( .A(n_40), .Y(n_504) );
INVx1_ASAP7_75t_L g206 ( .A(n_42), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g441 ( .A1(n_43), .A2(n_128), .B(n_196), .C(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_44), .B(n_151), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_45), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_46), .Y(n_537) );
INVx1_ASAP7_75t_L g471 ( .A(n_47), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_48), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_49), .B(n_110), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_50), .A2(n_118), .B1(n_184), .B2(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_51), .Y(n_138) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_52), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_53), .A2(n_196), .B(n_197), .C(n_199), .Y(n_195) );
CKINVDCx14_ASAP7_75t_R g440 ( .A(n_54), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_55), .Y(n_246) );
INVx1_ASAP7_75t_L g194 ( .A(n_56), .Y(n_194) );
INVx1_ASAP7_75t_L g116 ( .A(n_57), .Y(n_116) );
INVx1_ASAP7_75t_L g135 ( .A(n_58), .Y(n_135) );
INVx1_ASAP7_75t_SL g507 ( .A(n_59), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_60), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_61), .B(n_191), .Y(n_475) );
INVx1_ASAP7_75t_L g496 ( .A(n_62), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_SL g216 ( .A1(n_63), .A2(n_126), .B(n_199), .C(n_217), .Y(n_216) );
INVxp67_ASAP7_75t_L g218 ( .A(n_64), .Y(n_218) );
INVx1_ASAP7_75t_L g714 ( .A(n_65), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_66), .A2(n_110), .B(n_439), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_67), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_68), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_69), .A2(n_110), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g239 ( .A(n_70), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_71), .A2(n_161), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g450 ( .A(n_72), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_73), .Y(n_479) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_74), .A2(n_99), .B1(n_710), .B2(n_719), .C1(n_729), .C2(n_735), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g721 ( .A1(n_74), .A2(n_431), .B1(n_722), .B2(n_723), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_74), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_75), .A2(n_115), .B(n_118), .C(n_241), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_76), .A2(n_110), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g453 ( .A(n_77), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_78), .B(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
INVx1_ASAP7_75t_L g462 ( .A(n_80), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_81), .B(n_126), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_82), .A2(n_115), .B(n_118), .C(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g427 ( .A(n_83), .Y(n_427) );
OR2x2_ASAP7_75t_L g700 ( .A(n_83), .B(n_428), .Y(n_700) );
OR2x2_ASAP7_75t_L g718 ( .A(n_83), .B(n_705), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_84), .A2(n_118), .B(n_495), .C(n_498), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_85), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_86), .B(n_144), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_87), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_88), .A2(n_115), .B(n_118), .C(n_147), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_89), .Y(n_156) );
INVx1_ASAP7_75t_L g215 ( .A(n_90), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g163 ( .A(n_91), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_92), .B(n_123), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_93), .B(n_140), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_94), .B(n_140), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_95), .A2(n_110), .B(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g474 ( .A(n_96), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_97), .B(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_426), .B1(n_431), .B2(n_700), .Y(n_101) );
INVx2_ASAP7_75t_L g707 ( .A(n_102), .Y(n_707) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_395), .Y(n_102) );
NOR3xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_288), .C(n_361), .Y(n_103) );
OAI211xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_173), .B(n_220), .C(n_272), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_141), .Y(n_106) );
AND2x2_ASAP7_75t_L g236 ( .A(n_107), .B(n_237), .Y(n_236) );
INVx3_ASAP7_75t_L g255 ( .A(n_107), .Y(n_255) );
INVx2_ASAP7_75t_L g270 ( .A(n_107), .Y(n_270) );
INVx1_ASAP7_75t_L g300 ( .A(n_107), .Y(n_300) );
AND2x2_ASAP7_75t_L g350 ( .A(n_107), .B(n_271), .Y(n_350) );
AOI32xp33_ASAP7_75t_L g377 ( .A1(n_107), .A2(n_305), .A3(n_378), .B1(n_380), .B2(n_381), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_107), .B(n_226), .Y(n_383) );
AND2x2_ASAP7_75t_L g410 ( .A(n_107), .B(n_253), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_107), .B(n_419), .Y(n_418) );
OR2x6_ASAP7_75t_L g107 ( .A(n_108), .B(n_137), .Y(n_107) );
AOI21xp5_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_117), .B(n_130), .Y(n_108) );
BUFx2_ASAP7_75t_L g161 ( .A(n_110), .Y(n_161) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_115), .Y(n_110) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_111), .B(n_115), .Y(n_178) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
INVx1_ASAP7_75t_L g485 ( .A(n_112), .Y(n_485) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g119 ( .A(n_113), .Y(n_119) );
INVx1_ASAP7_75t_L g185 ( .A(n_113), .Y(n_185) );
INVx1_ASAP7_75t_L g120 ( .A(n_114), .Y(n_120) );
INVx3_ASAP7_75t_L g124 ( .A(n_114), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_114), .Y(n_126) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_114), .Y(n_167) );
INVx4_ASAP7_75t_SL g171 ( .A(n_115), .Y(n_171) );
BUFx3_ASAP7_75t_L g486 ( .A(n_115), .Y(n_486) );
INVx5_ASAP7_75t_L g164 ( .A(n_118), .Y(n_164) );
AND2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
BUFx3_ASAP7_75t_L g129 ( .A(n_119), .Y(n_129) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B(n_127), .Y(n_121) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_123), .A2(n_181), .B(n_182), .C(n_183), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_123), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_123), .A2(n_166), .B1(n_540), .B2(n_541), .Y(n_539) );
INVx5_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_124), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_124), .B(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_124), .B(n_443), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_127), .A2(n_242), .B(n_243), .Y(n_241) );
O2A1O1Ixp5_ASAP7_75t_L g461 ( .A1(n_127), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_127), .A2(n_463), .B(n_496), .C(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
INVx1_ASAP7_75t_L g244 ( .A(n_130), .Y(n_244) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_131), .A2(n_176), .B(n_186), .Y(n_175) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_131), .A2(n_203), .B(n_210), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_131), .B(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_133), .B(n_134), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
NOR2xp33_ASAP7_75t_SL g137 ( .A(n_138), .B(n_139), .Y(n_137) );
INVx3_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_139), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_139), .B(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_139), .A2(n_492), .B(n_499), .Y(n_491) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_140), .A2(n_213), .B(n_219), .Y(n_212) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_140), .Y(n_447) );
AND2x2_ASAP7_75t_L g299 ( .A(n_141), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g321 ( .A(n_141), .Y(n_321) );
AND2x2_ASAP7_75t_L g406 ( .A(n_141), .B(n_236), .Y(n_406) );
AND2x2_ASAP7_75t_L g409 ( .A(n_141), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_158), .Y(n_141) );
INVx2_ASAP7_75t_L g228 ( .A(n_142), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_142), .B(n_253), .Y(n_259) );
AND2x2_ASAP7_75t_L g269 ( .A(n_142), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g305 ( .A(n_142), .Y(n_305) );
AO21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B(n_155), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_143), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g544 ( .A(n_143), .Y(n_544) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_144), .A2(n_160), .B(n_172), .Y(n_159) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_144), .A2(n_438), .B(n_444), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_144), .A2(n_178), .B(n_479), .C(n_480), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_154), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_152), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_150), .B(n_507), .Y(n_506) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g199 ( .A(n_153), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_157), .B(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_157), .B(n_246), .Y(n_245) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_157), .A2(n_458), .B(n_465), .Y(n_457) );
AND2x2_ASAP7_75t_L g247 ( .A(n_158), .B(n_228), .Y(n_247) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g229 ( .A(n_159), .Y(n_229) );
AND2x2_ASAP7_75t_L g271 ( .A(n_159), .B(n_253), .Y(n_271) );
AND2x2_ASAP7_75t_L g340 ( .A(n_159), .B(n_237), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_165), .C(n_171), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_164), .A2(n_171), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_164), .A2(n_171), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g439 ( .A1(n_164), .A2(n_171), .B(n_440), .C(n_441), .Y(n_439) );
O2A1O1Ixp33_ASAP7_75t_SL g449 ( .A1(n_164), .A2(n_171), .B(n_450), .C(n_451), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_SL g470 ( .A1(n_164), .A2(n_171), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_164), .A2(n_171), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_164), .A2(n_171), .B(n_537), .C(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_166), .B(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_166), .B(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_166), .B(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI22xp5_ASAP7_75t_SL g205 ( .A1(n_167), .A2(n_206), .B1(n_207), .B2(n_208), .Y(n_205) );
INVx2_ASAP7_75t_L g207 ( .A(n_167), .Y(n_207) );
OAI22xp33_ASAP7_75t_L g203 ( .A1(n_171), .A2(n_178), .B1(n_204), .B2(n_209), .Y(n_203) );
INVx1_ASAP7_75t_L g498 ( .A(n_171), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_188), .Y(n_173) );
OR2x2_ASAP7_75t_L g234 ( .A(n_174), .B(n_202), .Y(n_234) );
INVx1_ASAP7_75t_L g313 ( .A(n_174), .Y(n_313) );
AND2x2_ASAP7_75t_L g327 ( .A(n_174), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_174), .B(n_201), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_174), .B(n_325), .Y(n_379) );
AND2x2_ASAP7_75t_L g387 ( .A(n_174), .B(n_388), .Y(n_387) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g224 ( .A(n_175), .Y(n_224) );
AND2x2_ASAP7_75t_L g294 ( .A(n_175), .B(n_202), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_178), .A2(n_239), .B(n_240), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_178), .A2(n_459), .B(n_460), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_178), .A2(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_188), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g421 ( .A(n_188), .Y(n_421) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_201), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_189), .B(n_265), .Y(n_287) );
OR2x2_ASAP7_75t_L g316 ( .A(n_189), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g348 ( .A(n_189), .B(n_328), .Y(n_348) );
INVx1_ASAP7_75t_SL g368 ( .A(n_189), .Y(n_368) );
AND2x2_ASAP7_75t_L g372 ( .A(n_189), .B(n_233), .Y(n_372) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_SL g225 ( .A(n_190), .B(n_201), .Y(n_225) );
AND2x2_ASAP7_75t_L g232 ( .A(n_190), .B(n_212), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_190), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g275 ( .A(n_190), .B(n_257), .Y(n_275) );
INVx1_ASAP7_75t_SL g282 ( .A(n_190), .Y(n_282) );
BUFx2_ASAP7_75t_L g293 ( .A(n_190), .Y(n_293) );
AND2x2_ASAP7_75t_L g309 ( .A(n_190), .B(n_224), .Y(n_309) );
AND2x2_ASAP7_75t_L g324 ( .A(n_190), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g388 ( .A(n_190), .B(n_202), .Y(n_388) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_200), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_201), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g312 ( .A(n_201), .B(n_313), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_201), .A2(n_330), .B1(n_333), .B2(n_336), .C(n_341), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_201), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_212), .Y(n_201) );
INVx3_ASAP7_75t_L g257 ( .A(n_202), .Y(n_257) );
INVx2_ASAP7_75t_L g463 ( .A(n_207), .Y(n_463) );
BUFx2_ASAP7_75t_L g267 ( .A(n_212), .Y(n_267) );
AND2x2_ASAP7_75t_L g281 ( .A(n_212), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g298 ( .A(n_212), .Y(n_298) );
OR2x2_ASAP7_75t_L g317 ( .A(n_212), .B(n_257), .Y(n_317) );
INVx3_ASAP7_75t_L g325 ( .A(n_212), .Y(n_325) );
AND2x2_ASAP7_75t_L g328 ( .A(n_212), .B(n_257), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_226), .B1(n_230), .B2(n_235), .C(n_248), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_223), .B(n_297), .Y(n_422) );
OR2x2_ASAP7_75t_L g425 ( .A(n_223), .B(n_256), .Y(n_425) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
OAI221xp5_ASAP7_75t_SL g248 ( .A1(n_224), .A2(n_249), .B1(n_256), .B2(n_258), .C(n_261), .Y(n_248) );
AND2x2_ASAP7_75t_L g265 ( .A(n_224), .B(n_257), .Y(n_265) );
AND2x2_ASAP7_75t_L g273 ( .A(n_224), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_224), .B(n_281), .Y(n_280) );
NAND2x1_ASAP7_75t_L g323 ( .A(n_224), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g375 ( .A(n_224), .B(n_317), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_226), .A2(n_335), .B1(n_364), .B2(n_366), .Y(n_363) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AOI322xp5_ASAP7_75t_L g272 ( .A1(n_227), .A2(n_236), .A3(n_273), .B1(n_276), .B2(n_279), .C1(n_283), .C2(n_286), .Y(n_272) );
OR2x2_ASAP7_75t_L g284 ( .A(n_227), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_228), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g263 ( .A(n_228), .B(n_237), .Y(n_263) );
INVx1_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
AND2x2_ASAP7_75t_L g344 ( .A(n_228), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g254 ( .A(n_229), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g345 ( .A(n_229), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_229), .B(n_253), .Y(n_419) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_233), .B(n_368), .Y(n_367) );
INVx3_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g319 ( .A(n_234), .B(n_266), .Y(n_319) );
OR2x2_ASAP7_75t_L g416 ( .A(n_234), .B(n_267), .Y(n_416) );
INVx1_ASAP7_75t_L g397 ( .A(n_235), .Y(n_397) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_247), .Y(n_235) );
INVx4_ASAP7_75t_L g285 ( .A(n_236), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_236), .B(n_304), .Y(n_310) );
INVx2_ASAP7_75t_L g253 ( .A(n_237), .Y(n_253) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_244), .B(n_245), .Y(n_237) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_244), .A2(n_534), .B(n_542), .Y(n_533) );
INVx1_ASAP7_75t_L g551 ( .A(n_244), .Y(n_551) );
INVx1_ASAP7_75t_L g335 ( .A(n_247), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_247), .B(n_307), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g322 ( .A1(n_249), .A2(n_323), .B(n_326), .Y(n_322) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_254), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g307 ( .A(n_253), .Y(n_307) );
INVx1_ASAP7_75t_L g334 ( .A(n_253), .Y(n_334) );
INVx1_ASAP7_75t_L g260 ( .A(n_254), .Y(n_260) );
AND2x2_ASAP7_75t_L g262 ( .A(n_254), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g358 ( .A(n_255), .B(n_344), .Y(n_358) );
AND2x2_ASAP7_75t_L g380 ( .A(n_255), .B(n_340), .Y(n_380) );
BUFx2_ASAP7_75t_L g332 ( .A(n_257), .Y(n_332) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AOI32xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_264), .A3(n_265), .B1(n_266), .B2(n_268), .Y(n_261) );
INVx1_ASAP7_75t_L g342 ( .A(n_262), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_262), .A2(n_390), .B1(n_391), .B2(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_265), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_265), .B(n_324), .Y(n_365) );
AND2x2_ASAP7_75t_L g412 ( .A(n_265), .B(n_297), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_266), .B(n_313), .Y(n_360) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g413 ( .A(n_268), .Y(n_413) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g338 ( .A(n_269), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_271), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g385 ( .A(n_271), .B(n_305), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_271), .B(n_300), .Y(n_392) );
INVx1_ASAP7_75t_SL g374 ( .A(n_273), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_274), .B(n_325), .Y(n_352) );
NOR4xp25_ASAP7_75t_L g398 ( .A(n_274), .B(n_297), .C(n_399), .D(n_402), .Y(n_398) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_275), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_L g355 ( .A(n_278), .Y(n_355) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_281), .A2(n_372), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g297 ( .A(n_282), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g346 ( .A(n_285), .Y(n_346) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND4xp25_ASAP7_75t_SL g288 ( .A(n_289), .B(n_314), .C(n_329), .D(n_349), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_295), .B(n_299), .C(n_301), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g381 ( .A(n_294), .B(n_324), .Y(n_381) );
AND2x2_ASAP7_75t_L g390 ( .A(n_294), .B(n_368), .Y(n_390) );
INVx3_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_297), .B(n_332), .Y(n_394) );
AND2x2_ASAP7_75t_L g306 ( .A(n_300), .B(n_307), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_308), .B1(n_310), .B2(n_311), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
AND2x2_ASAP7_75t_L g404 ( .A(n_304), .B(n_350), .Y(n_404) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_306), .B(n_355), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_307), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B(n_320), .C(n_322), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_315), .A2(n_350), .B1(n_351), .B2(n_353), .C(n_356), .Y(n_349) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_323), .A2(n_408), .B1(n_411), .B2(n_413), .C(n_414), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_324), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_332), .B(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g362 ( .A(n_334), .Y(n_362) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_337), .A2(n_357), .B1(n_359), .B2(n_360), .Y(n_356) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI21xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B(n_347), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_346), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_357), .A2(n_383), .B1(n_421), .B2(n_422), .C(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g402 ( .A(n_359), .Y(n_402) );
OAI211xp5_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_363), .B(n_369), .C(n_389), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI211xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_372), .B(n_373), .C(n_382), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
A2O1A1Ixp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B(n_376), .C(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g423 ( .A1(n_380), .A2(n_406), .B(n_424), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_386), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI21xp5_ASAP7_75t_SL g415 ( .A1(n_392), .A2(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_407), .C(n_420), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_403), .C(n_405), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
CKINVDCx14_ASAP7_75t_R g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g709 ( .A(n_426), .Y(n_709) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NOR2x2_ASAP7_75t_L g704 ( .A(n_427), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_428), .Y(n_705) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g722 ( .A(n_431), .Y(n_722) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g706 ( .A1(n_432), .A2(n_700), .B1(n_707), .B2(n_708), .Y(n_706) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_630), .Y(n_432) );
NAND5xp2_ASAP7_75t_L g433 ( .A(n_434), .B(n_545), .C(n_577), .D(n_594), .E(n_617), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_476), .B1(n_509), .B2(n_513), .C(n_517), .Y(n_434) );
INVx1_ASAP7_75t_L g657 ( .A(n_435), .Y(n_657) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_455), .Y(n_435) );
AND3x2_ASAP7_75t_L g632 ( .A(n_436), .B(n_457), .C(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_445), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_437), .B(n_515), .Y(n_514) );
BUFx3_ASAP7_75t_L g524 ( .A(n_437), .Y(n_524) );
AND2x2_ASAP7_75t_L g528 ( .A(n_437), .B(n_467), .Y(n_528) );
INVx2_ASAP7_75t_L g554 ( .A(n_437), .Y(n_554) );
OR2x2_ASAP7_75t_L g565 ( .A(n_437), .B(n_468), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_437), .B(n_456), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_437), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g644 ( .A(n_437), .B(n_468), .Y(n_644) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_445), .Y(n_527) );
AND2x2_ASAP7_75t_L g585 ( .A(n_445), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_445), .B(n_456), .Y(n_604) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g516 ( .A(n_446), .B(n_456), .Y(n_516) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_446), .Y(n_523) );
AND2x2_ASAP7_75t_L g571 ( .A(n_446), .B(n_468), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g596 ( .A(n_446), .B(n_455), .C(n_554), .Y(n_596) );
AND2x2_ASAP7_75t_L g661 ( .A(n_446), .B(n_457), .Y(n_661) );
AND2x2_ASAP7_75t_L g695 ( .A(n_446), .B(n_456), .Y(n_695) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_454), .Y(n_446) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_447), .A2(n_469), .B(n_475), .Y(n_468) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_447), .A2(n_502), .B(n_508), .Y(n_501) );
INVxp67_ASAP7_75t_L g525 ( .A(n_455), .Y(n_525) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_467), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_456), .B(n_554), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_456), .B(n_585), .Y(n_593) );
AND2x2_ASAP7_75t_L g643 ( .A(n_456), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g671 ( .A(n_456), .Y(n_671) );
INVx4_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g578 ( .A(n_457), .B(n_571), .Y(n_578) );
BUFx3_ASAP7_75t_L g610 ( .A(n_457), .Y(n_610) );
INVx2_ASAP7_75t_L g586 ( .A(n_467), .Y(n_586) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_468), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_476), .A2(n_646), .B1(n_648), .B2(n_649), .Y(n_645) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_489), .Y(n_476) );
AND2x2_ASAP7_75t_L g509 ( .A(n_477), .B(n_510), .Y(n_509) );
INVx3_ASAP7_75t_SL g520 ( .A(n_477), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_477), .B(n_549), .Y(n_581) );
OR2x2_ASAP7_75t_L g600 ( .A(n_477), .B(n_490), .Y(n_600) );
AND2x2_ASAP7_75t_L g605 ( .A(n_477), .B(n_557), .Y(n_605) );
AND2x2_ASAP7_75t_L g608 ( .A(n_477), .B(n_550), .Y(n_608) );
AND2x2_ASAP7_75t_L g620 ( .A(n_477), .B(n_501), .Y(n_620) );
AND2x2_ASAP7_75t_L g636 ( .A(n_477), .B(n_491), .Y(n_636) );
AND2x4_ASAP7_75t_L g639 ( .A(n_477), .B(n_511), .Y(n_639) );
OR2x2_ASAP7_75t_L g656 ( .A(n_477), .B(n_592), .Y(n_656) );
OR2x2_ASAP7_75t_L g687 ( .A(n_477), .B(n_533), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_477), .B(n_615), .Y(n_689) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_487), .Y(n_477) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_485), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g563 ( .A(n_489), .B(n_531), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_489), .B(n_550), .Y(n_682) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_501), .Y(n_489) );
AND2x2_ASAP7_75t_L g519 ( .A(n_490), .B(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g549 ( .A(n_490), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g557 ( .A(n_490), .B(n_533), .Y(n_557) );
AND2x2_ASAP7_75t_L g575 ( .A(n_490), .B(n_511), .Y(n_575) );
OR2x2_ASAP7_75t_L g592 ( .A(n_490), .B(n_550), .Y(n_592) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g512 ( .A(n_491), .Y(n_512) );
AND2x2_ASAP7_75t_L g615 ( .A(n_491), .B(n_501), .Y(n_615) );
INVx2_ASAP7_75t_L g511 ( .A(n_501), .Y(n_511) );
INVx1_ASAP7_75t_L g627 ( .A(n_501), .Y(n_627) );
AND2x2_ASAP7_75t_L g677 ( .A(n_501), .B(n_520), .Y(n_677) );
AND2x2_ASAP7_75t_L g530 ( .A(n_510), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g561 ( .A(n_510), .B(n_520), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_510), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
AND2x2_ASAP7_75t_L g548 ( .A(n_511), .B(n_520), .Y(n_548) );
OR2x2_ASAP7_75t_L g664 ( .A(n_512), .B(n_638), .Y(n_664) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_515), .B(n_644), .Y(n_650) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
OAI32xp33_ASAP7_75t_L g606 ( .A1(n_516), .A2(n_607), .A3(n_609), .B1(n_611), .B2(n_612), .Y(n_606) );
OR2x2_ASAP7_75t_L g623 ( .A(n_516), .B(n_565), .Y(n_623) );
OAI21xp33_ASAP7_75t_SL g648 ( .A1(n_516), .A2(n_526), .B(n_553), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_521), .B1(n_526), .B2(n_529), .Y(n_517) );
INVxp33_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_519), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_520), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g574 ( .A(n_520), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g674 ( .A(n_520), .B(n_615), .Y(n_674) );
OR2x2_ASAP7_75t_L g698 ( .A(n_520), .B(n_592), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_521), .A2(n_580), .B(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g558 ( .A(n_523), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_523), .B(n_528), .Y(n_576) );
AND2x2_ASAP7_75t_L g598 ( .A(n_524), .B(n_571), .Y(n_598) );
INVx1_ASAP7_75t_L g611 ( .A(n_524), .Y(n_611) );
OR2x2_ASAP7_75t_L g616 ( .A(n_524), .B(n_550), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_527), .B(n_565), .Y(n_564) );
OAI22xp33_ASAP7_75t_L g546 ( .A1(n_528), .A2(n_547), .B1(n_552), .B2(n_556), .Y(n_546) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_531), .A2(n_589), .B1(n_596), .B2(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g673 ( .A(n_531), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_533), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g692 ( .A(n_533), .B(n_575), .Y(n_692) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_535), .A2(n_543), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_558), .B1(n_559), .B2(n_564), .C(n_566), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_548), .B(n_550), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_548), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g567 ( .A(n_549), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_549), .A2(n_655), .B(n_656), .C(n_657), .Y(n_654) );
AND2x2_ASAP7_75t_L g659 ( .A(n_549), .B(n_639), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_SL g697 ( .A1(n_549), .A2(n_638), .B(n_698), .C(n_699), .Y(n_697) );
BUFx3_ASAP7_75t_L g589 ( .A(n_550), .Y(n_589) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_553), .B(n_610), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_553), .A2(n_673), .B(n_675), .C(n_681), .Y(n_672) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVxp67_ASAP7_75t_L g633 ( .A(n_555), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_557), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_560), .B(n_562), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AOI211xp5_ASAP7_75t_L g577 ( .A1(n_561), .A2(n_578), .B(n_579), .C(n_587), .Y(n_577) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g662 ( .A(n_565), .Y(n_662) );
OR2x2_ASAP7_75t_L g679 ( .A(n_565), .B(n_609), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_573), .B2(n_576), .Y(n_566) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_568), .A2(n_580), .B1(n_581), .B2(n_582), .Y(n_579) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
OR2x2_ASAP7_75t_L g666 ( .A(n_570), .B(n_610), .Y(n_666) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g621 ( .A(n_571), .B(n_611), .Y(n_621) );
INVx1_ASAP7_75t_L g629 ( .A(n_572), .Y(n_629) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_575), .B(n_589), .Y(n_637) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_585), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g694 ( .A(n_586), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_590), .B(n_593), .Y(n_587) );
INVx1_ASAP7_75t_L g624 ( .A(n_588), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_589), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_589), .B(n_620), .Y(n_619) );
NAND2x1p5_ASAP7_75t_L g640 ( .A(n_589), .B(n_615), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_589), .B(n_636), .Y(n_647) );
OAI211xp5_ASAP7_75t_L g651 ( .A1(n_589), .A2(n_599), .B(n_639), .C(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_599), .B1(n_601), .B2(n_605), .C(n_606), .Y(n_594) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_603), .B(n_611), .Y(n_685) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_605), .A2(n_620), .B(n_622), .C(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_608), .B(n_615), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_609), .B(n_662), .Y(n_699) );
CKINVDCx16_ASAP7_75t_R g609 ( .A(n_610), .Y(n_609) );
INVxp33_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
AOI21xp33_ASAP7_75t_SL g625 ( .A1(n_614), .A2(n_626), .B(n_628), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_614), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_615), .B(n_669), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B1(n_622), .B2(n_624), .C(n_625), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_621), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g655 ( .A(n_627), .Y(n_655) );
NAND5xp2_ASAP7_75t_L g630 ( .A(n_631), .B(n_658), .C(n_672), .D(n_683), .E(n_696), .Y(n_630) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B(n_641), .C(n_654), .Y(n_631) );
INVx2_ASAP7_75t_SL g678 ( .A(n_632), .Y(n_678) );
NAND4xp25_ASAP7_75t_SL g634 ( .A(n_635), .B(n_637), .C(n_638), .D(n_640), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI211xp5_ASAP7_75t_SL g641 ( .A1(n_640), .A2(n_642), .B(n_645), .C(n_651), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_643), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_643), .A2(n_684), .B1(n_686), .B2(n_688), .C(n_690), .Y(n_683) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI221xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_660), .B1(n_663), .B2(n_665), .C(n_667), .Y(n_658) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_666), .A2(n_689), .B1(n_691), .B2(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B1(n_679), .B2(n_680), .Y(n_675) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx3_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_716), .Y(n_711) );
NOR2xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_715), .Y(n_712) );
INVx1_ASAP7_75t_SL g734 ( .A(n_713), .Y(n_734) );
INVx1_ASAP7_75t_L g733 ( .A(n_715), .Y(n_733) );
OA21x2_ASAP7_75t_L g736 ( .A1(n_715), .A2(n_734), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g725 ( .A(n_718), .Y(n_725) );
BUFx2_ASAP7_75t_L g737 ( .A(n_718), .Y(n_737) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_724), .B(n_726), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g728 ( .A(n_725), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
CKINVDCx6p67_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
endmodule