module fake_jpeg_16028_n_354 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_354);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_48),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_0),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_27),
.B(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_25),
.Y(n_65)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_62),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_17),
.B1(n_19),
.B2(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_64),
.B1(n_69),
.B2(n_36),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_42),
.B1(n_38),
.B2(n_17),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_48),
.B1(n_51),
.B2(n_47),
.Y(n_99)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_17),
.B1(n_19),
.B2(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_67),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_25),
.B1(n_34),
.B2(n_32),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_29),
.B1(n_36),
.B2(n_32),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_79),
.A2(n_105),
.B1(n_83),
.B2(n_20),
.Y(n_138)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_92),
.Y(n_123)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_107),
.B1(n_75),
.B2(n_70),
.Y(n_112)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_100),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_54),
.Y(n_97)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_104),
.B1(n_52),
.B2(n_44),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_102),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_59),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_51),
.B1(n_47),
.B2(n_45),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_70),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_40),
.B1(n_44),
.B2(n_41),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_60),
.A2(n_72),
.B1(n_66),
.B2(n_40),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_45),
.B1(n_18),
.B2(n_20),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_108),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_49),
.C(n_39),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_39),
.C(n_49),
.Y(n_134)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_121),
.B1(n_101),
.B2(n_97),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_55),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_125),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_107),
.B1(n_90),
.B2(n_83),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_119),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_124),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_81),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_22),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_52),
.B1(n_63),
.B2(n_74),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_94),
.B1(n_101),
.B2(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_22),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_52),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_74),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_77),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_98),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_138),
.A2(n_108),
.B1(n_86),
.B2(n_105),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_109),
.C(n_99),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_141),
.B(n_154),
.C(n_172),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_143),
.A2(n_18),
.B1(n_16),
.B2(n_15),
.Y(n_198)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_117),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_149),
.A2(n_133),
.B1(n_33),
.B2(n_24),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_151),
.B1(n_137),
.B2(n_111),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_78),
.B1(n_87),
.B2(n_105),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_159),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_89),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_146),
.Y(n_191)
);

NOR2x1_ASAP7_75t_R g155 ( 
.A(n_125),
.B(n_91),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_155),
.A2(n_115),
.B(n_128),
.Y(n_186)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

BUFx24_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_127),
.B(n_13),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_164),
.B(n_135),
.Y(n_195)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_63),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_129),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_110),
.B1(n_11),
.B2(n_12),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_116),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_113),
.A2(n_20),
.B1(n_18),
.B2(n_28),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_20),
.B1(n_18),
.B2(n_23),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_33),
.C(n_23),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_145),
.B(n_127),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_190),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_115),
.Y(n_175)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_185),
.B1(n_147),
.B2(n_149),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_169),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_177),
.B(n_192),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_179),
.B(n_3),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_131),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_181),
.B(n_4),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_116),
.B(n_114),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_182),
.A2(n_184),
.B(n_186),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_155),
.A2(n_136),
.B(n_131),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_116),
.B1(n_114),
.B2(n_111),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_198),
.B1(n_203),
.B2(n_158),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_145),
.B(n_124),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_128),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_24),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_205),
.C(n_133),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_157),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_196),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_156),
.A2(n_133),
.B(n_1),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_172),
.B(n_167),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_142),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_142),
.B(n_0),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_158),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_206),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_209),
.B(n_229),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_214),
.B1(n_219),
.B2(n_222),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_212),
.A2(n_218),
.B(n_204),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_168),
.B1(n_148),
.B2(n_165),
.Y(n_214)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_207),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_170),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_221),
.C(n_223),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_24),
.B(n_33),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_15),
.C(n_14),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_224),
.A2(n_199),
.B1(n_182),
.B2(n_178),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_14),
.C(n_10),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_228),
.C(n_233),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_179),
.C(n_191),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_16),
.B1(n_14),
.B2(n_10),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_174),
.B1(n_208),
.B2(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_177),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_192),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_2),
.C(n_3),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_196),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_234),
.B(n_236),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_235),
.B(n_186),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_173),
.B(n_4),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_189),
.Y(n_255)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_187),
.C(n_180),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_212),
.B(n_224),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_222),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_190),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_245),
.B(n_253),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_249),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_248),
.B(n_223),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_220),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_220),
.A2(n_188),
.B1(n_187),
.B2(n_199),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_258),
.B1(n_261),
.B2(n_216),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_211),
.Y(n_254)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_235),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_189),
.B1(n_197),
.B2(n_201),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_259),
.Y(n_265)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_260),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_214),
.A2(n_201),
.B1(n_5),
.B2(n_6),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_4),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_227),
.C(n_233),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_273),
.Y(n_296)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_232),
.B1(n_217),
.B2(n_221),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_285),
.B1(n_252),
.B2(n_244),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_232),
.B(n_218),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_272),
.A2(n_253),
.B(n_240),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_248),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_256),
.B(n_237),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_282),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_257),
.C(n_262),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_257),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_276),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_300),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_251),
.B1(n_249),
.B2(n_259),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_297),
.B1(n_299),
.B2(n_270),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_246),
.Y(n_290)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_285),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_279),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_295),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_267),
.A2(n_258),
.B1(n_240),
.B2(n_241),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_272),
.A2(n_250),
.B(n_238),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_274),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_302),
.B(n_4),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_277),
.A2(n_263),
.B(n_261),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_283),
.C(n_271),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_306),
.C(n_317),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_305),
.B(n_304),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_282),
.C(n_281),
.Y(n_306)
);

OAI221xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_264),
.B1(n_268),
.B2(n_275),
.C(n_265),
.Y(n_308)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_316),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_289),
.B(n_286),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_273),
.B1(n_280),
.B2(n_269),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_314),
.B1(n_298),
.B2(n_288),
.Y(n_326)
);

XOR2x1_ASAP7_75t_SL g315 ( 
.A(n_301),
.B(n_6),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_7),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_7),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_7),
.C(n_8),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_7),
.C(n_9),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_302),
.C(n_297),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_319),
.B(n_324),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_326),
.C(n_9),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_327),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_312),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_291),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_293),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_321),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_306),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_334),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_315),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_333),
.B(n_339),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_316),
.B(n_317),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_323),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_318),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_330),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_340),
.B(n_342),
.Y(n_348)
);

AOI21x1_ASAP7_75t_L g342 ( 
.A1(n_338),
.A2(n_327),
.B(n_324),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_344),
.B(n_345),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_9),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_341),
.A2(n_338),
.B(n_344),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_336),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_350),
.A2(n_343),
.B(n_331),
.C(n_348),
.Y(n_351)
);

BUFx24_ASAP7_75t_SL g352 ( 
.A(n_351),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_352),
.A2(n_346),
.B(n_9),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);


endmodule