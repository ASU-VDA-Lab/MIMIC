module fake_jpeg_2634_n_78 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_31),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_20),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_34)
);

AO22x2_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_28),
.B1(n_32),
.B2(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_25),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_46),
.B1(n_47),
.B2(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_45),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_29),
.B1(n_32),
.B2(n_21),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_32),
.B1(n_26),
.B2(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_50),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_18),
.B1(n_16),
.B2(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_34),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_29),
.C(n_35),
.Y(n_51)
);

FAx1_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_13),
.CI(n_12),
.CON(n_61),
.SN(n_61)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_0),
.Y(n_58)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_4),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_29),
.B(n_35),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_61),
.B(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_1),
.B(n_3),
.Y(n_59)
);

XNOR2x1_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_55),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

A2O1A1O1Ixp25_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_54),
.B(n_10),
.C(n_7),
.D(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

AO221x1_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_61),
.B1(n_60),
.B2(n_9),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_67),
.B(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

AOI31xp33_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_72),
.A3(n_65),
.B(n_71),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_66),
.B(n_70),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_5),
.C(n_6),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_9),
.Y(n_78)
);


endmodule