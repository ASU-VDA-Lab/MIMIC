module real_jpeg_2154_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_205;
wire n_61;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_167;
wire n_244;
wire n_179;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_45),
.B1(n_58),
.B2(n_60),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_28),
.B1(n_34),
.B2(n_45),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_52),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_2),
.A2(n_52),
.B1(n_58),
.B2(n_60),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_2),
.A2(n_28),
.B1(n_34),
.B2(n_52),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_3),
.A2(n_72),
.B1(n_73),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_3),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_58),
.B1(n_60),
.B2(n_81),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_81),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_28),
.B1(n_34),
.B2(n_81),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_5),
.A2(n_72),
.B1(n_73),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_5),
.A2(n_58),
.B1(n_60),
.B2(n_79),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_79),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_5),
.A2(n_28),
.B1(n_34),
.B2(n_79),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_6),
.B(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_6),
.B(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_6),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_6),
.A2(n_72),
.B(n_136),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_6),
.B(n_62),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_6),
.A2(n_60),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_6),
.B(n_28),
.C(n_48),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_172),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_6),
.B(n_31),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_6),
.B(n_53),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_11),
.A2(n_28),
.B1(n_34),
.B2(n_57),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_13),
.A2(n_72),
.B1(n_73),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_13),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_13),
.A2(n_58),
.B1(n_60),
.B2(n_124),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_124),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_13),
.A2(n_28),
.B1(n_34),
.B2(n_124),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_72),
.B1(n_73),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_14),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_58),
.B1(n_60),
.B2(n_146),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_146),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_14),
.A2(n_28),
.B1(n_34),
.B2(n_146),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_15),
.A2(n_28),
.B1(n_34),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_15),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_16),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_16),
.A2(n_35),
.B1(n_42),
.B2(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_126),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_108),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_21),
.B(n_108),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_54),
.C(n_68),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_23),
.A2(n_24),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_25),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_148)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_27),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_27),
.A2(n_31),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_27),
.A2(n_31),
.B1(n_139),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_27),
.A2(n_31),
.B1(n_176),
.B2(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_27),
.A2(n_31),
.B1(n_172),
.B2(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_27),
.A2(n_31),
.B1(n_225),
.B2(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_28),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_28),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_28),
.B(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_30),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_30),
.A2(n_33),
.B1(n_96),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_30),
.A2(n_96),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_30),
.A2(n_96),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_41),
.A2(n_50),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

AO22x2_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_43),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_42),
.B(n_64),
.Y(n_173)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_43),
.A2(n_60),
.A3(n_63),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_43),
.B(n_213),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_53),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_46),
.A2(n_53),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_46),
.A2(n_53),
.B1(n_168),
.B2(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_46),
.A2(n_53),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_46),
.A2(n_53),
.B1(n_195),
.B2(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_50),
.A2(n_117),
.B1(n_167),
.B2(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_62),
.B1(n_86),
.B2(n_121),
.Y(n_120)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_60),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_58),
.B(n_74),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_58),
.B(n_172),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_60),
.A2(n_73),
.A3(n_75),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_61),
.A2(n_67),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_61),
.A2(n_67),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_61),
.A2(n_67),
.B1(n_142),
.B2(n_158),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_61),
.A2(n_67),
.B1(n_157),
.B2(n_204),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_63),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_69),
.A2(n_76),
.B1(n_80),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_69),
.A2(n_76),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_69),
.A2(n_76),
.B1(n_145),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_70),
.A2(n_78),
.B1(n_123),
.B2(n_125),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_92),
.B1(n_93),
.B2(n_107),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_88),
.B(n_91),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_100),
.B1(n_101),
.B2(n_106),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_113),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_120),
.C(n_122),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_115),
.B(n_118),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_122),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_151),
.B(n_260),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_149),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_130),
.B(n_149),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_148),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_131),
.B(n_148),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_133),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.C(n_144),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_134),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_138),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_141),
.B(n_144),
.Y(n_251)
);

AOI31xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_245),
.A3(n_254),
.B(n_257),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_190),
.B(n_244),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_178),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_154),
.B(n_178),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_165),
.C(n_169),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_155),
.B(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_160),
.C(n_164),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_165),
.B(n_169),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_178),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_178),
.B(n_255),
.Y(n_258)
);

FAx1_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.CI(n_181),
.CON(n_178),
.SN(n_178)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_182),
.B(n_185),
.C(n_189),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_239),
.B(n_243),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_208),
.B(n_238),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_200),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_200),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_197),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_203),
.C(n_206),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_219),
.B(n_237),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_217),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_231),
.B(n_236),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_226),
.B(n_230),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_228),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_235),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_242),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_249),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.C(n_253),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_253),
.Y(n_256)
);


endmodule