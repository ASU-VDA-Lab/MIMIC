module fake_jpeg_1513_n_542 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_542);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx11_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g166 ( 
.A(n_52),
.Y(n_166)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_99),
.Y(n_117)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_90),
.Y(n_104)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_32),
.Y(n_89)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_32),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_18),
.B(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_100),
.Y(n_107)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_98),
.Y(n_156)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_51),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_43),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_23),
.B1(n_43),
.B2(n_51),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_105),
.A2(n_126),
.B1(n_50),
.B2(n_70),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_45),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_121),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_54),
.B(n_30),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_60),
.A2(n_43),
.B1(n_50),
.B2(n_48),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_37),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_130),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_46),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_24),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_87),
.B(n_37),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_56),
.B(n_19),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_19),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_26),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_160),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_26),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_55),
.B(n_34),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_164),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_53),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_72),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_58),
.B(n_25),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVx4_ASAP7_75t_SL g274 ( 
.A(n_167),
.Y(n_274)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_169),
.Y(n_246)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_171),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_131),
.A2(n_65),
.B1(n_20),
.B2(n_46),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_172),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_104),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_174),
.B(n_192),
.Y(n_238)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_175),
.Y(n_268)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_117),
.B(n_24),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_184),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_144),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_144),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_47),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_98),
.B1(n_96),
.B2(n_88),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_188),
.A2(n_220),
.B1(n_125),
.B2(n_152),
.Y(n_249)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_190),
.Y(n_265)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_112),
.Y(n_191)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_191),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_114),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_107),
.B(n_47),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

CKINVDCx12_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_34),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_199),
.Y(n_244)
);

CKINVDCx6p67_ASAP7_75t_R g198 ( 
.A(n_113),
.Y(n_198)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_135),
.B(n_40),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_105),
.A2(n_86),
.B1(n_85),
.B2(n_80),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_200),
.A2(n_152),
.B1(n_151),
.B2(n_122),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_116),
.A2(n_48),
.B1(n_51),
.B2(n_50),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_202),
.A2(n_188),
.B(n_172),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_158),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_203),
.B(n_207),
.Y(n_257)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_136),
.B(n_25),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_40),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_208),
.B(n_209),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_150),
.B(n_36),
.Y(n_209)
);

AOI32xp33_ASAP7_75t_L g210 ( 
.A1(n_131),
.A2(n_41),
.A3(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_210),
.B(n_212),
.Y(n_278)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_129),
.B(n_41),
.Y(n_212)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_138),
.B(n_39),
.Y(n_214)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_214),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_137),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_223),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_129),
.B(n_14),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_217),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_140),
.B(n_14),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_124),
.Y(n_218)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_218),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_126),
.A2(n_78),
.B1(n_77),
.B2(n_75),
.Y(n_220)
);

CKINVDCx6p67_ASAP7_75t_R g221 ( 
.A(n_139),
.Y(n_221)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_221),
.Y(n_277)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_224),
.Y(n_272)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_139),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_157),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_177),
.B(n_142),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_241),
.B(n_254),
.C(n_2),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_146),
.B(n_137),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_242),
.A2(n_227),
.B(n_167),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_194),
.A2(n_66),
.B1(n_71),
.B2(n_68),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_245),
.A2(n_255),
.B1(n_260),
.B2(n_262),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_249),
.A2(n_204),
.B1(n_205),
.B2(n_183),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_251),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_253),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_170),
.B(n_109),
.C(n_142),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_193),
.A2(n_125),
.B1(n_151),
.B2(n_123),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_219),
.A2(n_143),
.B1(n_133),
.B2(n_132),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_200),
.A2(n_123),
.B1(n_132),
.B2(n_143),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_263),
.A2(n_255),
.B1(n_261),
.B2(n_226),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_178),
.A2(n_133),
.B1(n_148),
.B2(n_128),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_270),
.B1(n_279),
.B2(n_245),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_202),
.A2(n_128),
.B1(n_108),
.B2(n_148),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_182),
.A2(n_146),
.B1(n_35),
.B2(n_50),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_273),
.A2(n_167),
.B1(n_2),
.B2(n_4),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_222),
.A2(n_108),
.B1(n_35),
.B2(n_3),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_189),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_280),
.A2(n_291),
.B(n_250),
.Y(n_329)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_231),
.Y(n_281)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_281),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_241),
.B(n_223),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_295),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_283),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_287),
.Y(n_331)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_286),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_238),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_230),
.B(n_198),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_289),
.B(n_294),
.Y(n_327)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_290),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_221),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_292),
.A2(n_297),
.B1(n_306),
.B2(n_318),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_176),
.Y(n_293)
);

NAND2x1p5_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_232),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_266),
.B(n_198),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_257),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_222),
.B1(n_168),
.B2(n_213),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_181),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_299),
.B(n_313),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_244),
.B(n_221),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_300),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_206),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_301),
.B(n_302),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_259),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_270),
.A2(n_175),
.B1(n_171),
.B2(n_201),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_303),
.A2(n_308),
.B1(n_316),
.B2(n_256),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_247),
.B(n_225),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_305),
.B(n_312),
.Y(n_340)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_279),
.A2(n_211),
.B1(n_186),
.B2(n_185),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_309),
.A2(n_319),
.B(n_320),
.Y(n_343)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_236),
.Y(n_310)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_310),
.Y(n_364)
);

INVx11_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_311),
.A2(n_274),
.B1(n_268),
.B2(n_234),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_184),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_229),
.B(n_18),
.Y(n_313)
);

OA22x2_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_264),
.B1(n_234),
.B2(n_240),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_235),
.B(n_17),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_232),
.C(n_268),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_263),
.A2(n_262),
.B1(n_251),
.B2(n_235),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_248),
.B(n_15),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_317),
.B(n_12),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_246),
.A2(n_12),
.B1(n_11),
.B2(n_4),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_248),
.A2(n_246),
.B(n_258),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_272),
.A2(n_0),
.B(n_2),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_258),
.Y(n_322)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_323),
.B(n_233),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_236),
.A2(n_12),
.B1(n_11),
.B2(n_5),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_324),
.A2(n_275),
.B1(n_237),
.B2(n_265),
.Y(n_349)
);

O2A1O1Ixp33_ASAP7_75t_L g325 ( 
.A1(n_259),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_264),
.B(n_250),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_265),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_328),
.A2(n_329),
.B(n_350),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_276),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_326),
.C(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_335),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_321),
.A2(n_240),
.B1(n_239),
.B2(n_243),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_306),
.Y(n_375)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_346),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_304),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_351),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_349),
.A2(n_362),
.B1(n_363),
.B2(n_284),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_291),
.A2(n_275),
.B(n_237),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_280),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_322),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_358),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_310),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_357),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_291),
.A2(n_243),
.B(n_239),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_359),
.A2(n_360),
.B(n_361),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_309),
.A2(n_5),
.B(n_6),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_288),
.A2(n_5),
.B(n_7),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_297),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_292),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_331),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_369),
.B(n_371),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_370),
.B(n_315),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_327),
.Y(n_371)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_365),
.Y(n_373)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

OAI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_375),
.A2(n_349),
.B1(n_314),
.B2(n_334),
.Y(n_429)
);

BUFx24_ASAP7_75t_SL g376 ( 
.A(n_342),
.Y(n_376)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_376),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_381),
.Y(n_427)
);

INVx13_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

OA22x2_ASAP7_75t_L g382 ( 
.A1(n_333),
.A2(n_316),
.B1(n_308),
.B2(n_303),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_SL g425 ( 
.A1(n_382),
.A2(n_293),
.B(n_334),
.C(n_347),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_333),
.A2(n_284),
.B1(n_288),
.B2(n_305),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_383),
.A2(n_332),
.B1(n_293),
.B2(n_363),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_282),
.Y(n_384)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_355),
.Y(n_385)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_386),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_329),
.A2(n_319),
.B(n_302),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_388),
.A2(n_343),
.B(n_350),
.Y(n_406)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_390),
.B(n_392),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_287),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_391),
.B(n_394),
.Y(n_421)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_396),
.C(n_397),
.Y(n_404)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_335),
.Y(n_394)
);

INVx6_ASAP7_75t_SL g395 ( 
.A(n_328),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_SL g409 ( 
.A1(n_395),
.A2(n_398),
.B(n_367),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_330),
.B(n_281),
.C(n_286),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_296),
.C(n_285),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_343),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_357),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_402),
.Y(n_419)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_394),
.B(n_367),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_403),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_406),
.A2(n_407),
.B(n_423),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_387),
.A2(n_359),
.B(n_360),
.Y(n_407)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_409),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_338),
.C(n_344),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_413),
.C(n_417),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_399),
.A2(n_338),
.B(n_344),
.C(n_337),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_425),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_341),
.C(n_337),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_396),
.B(n_341),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_414),
.B(n_383),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_356),
.C(n_300),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_280),
.C(n_323),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_422),
.C(n_392),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_420),
.A2(n_379),
.B1(n_368),
.B2(n_386),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_364),
.C(n_339),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_387),
.A2(n_347),
.B(n_362),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_374),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_428),
.Y(n_454)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_429),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_378),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_377),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_431),
.B(n_294),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_395),
.A2(n_320),
.B(n_361),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_433),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_385),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_441),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_437),
.A2(n_438),
.B1(n_440),
.B2(n_445),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_405),
.A2(n_369),
.B1(n_372),
.B2(n_379),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_416),
.A2(n_368),
.B1(n_399),
.B2(n_398),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_442),
.B(n_449),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_401),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_417),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_410),
.B(n_372),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_444),
.B(n_290),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_421),
.A2(n_375),
.B1(n_382),
.B2(n_400),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_408),
.Y(n_446)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_446),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_407),
.A2(n_382),
.B1(n_400),
.B2(n_389),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_447),
.A2(n_425),
.B1(n_433),
.B2(n_334),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_289),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_455),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_452),
.B(n_453),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_354),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_411),
.B(n_354),
.Y(n_456)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_420),
.A2(n_382),
.B1(n_389),
.B2(n_402),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_457),
.A2(n_423),
.B1(n_425),
.B2(n_427),
.Y(n_472)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_432),
.Y(n_459)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_463),
.C(n_467),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_439),
.A2(n_418),
.B(n_406),
.Y(n_461)
);

AOI21xp33_ASAP7_75t_L g490 ( 
.A1(n_461),
.A2(n_373),
.B(n_440),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_443),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_455),
.Y(n_464)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_464),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_430),
.C(n_422),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_403),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_471),
.Y(n_487)
);

AO22x2_ASAP7_75t_L g470 ( 
.A1(n_457),
.A2(n_425),
.B1(n_403),
.B2(n_412),
.Y(n_470)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_470),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_415),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_472),
.A2(n_445),
.B1(n_458),
.B2(n_435),
.Y(n_488)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_474),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_426),
.C(n_424),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_476),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_419),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_426),
.C(n_364),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_478),
.A2(n_447),
.B1(n_434),
.B2(n_450),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_480),
.A2(n_390),
.B1(n_454),
.B2(n_298),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_482),
.B(n_475),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_466),
.A2(n_451),
.B1(n_450),
.B2(n_301),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_486),
.A2(n_489),
.B1(n_492),
.B2(n_493),
.Y(n_507)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_488),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_470),
.A2(n_435),
.B(n_458),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_490),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_478),
.A2(n_353),
.B(n_381),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_470),
.A2(n_428),
.B1(n_374),
.B2(n_353),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_497),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_470),
.A2(n_374),
.B1(n_307),
.B2(n_324),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_481),
.A2(n_311),
.B1(n_325),
.B2(n_10),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_498),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_468),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_506),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_464),
.C(n_467),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_502),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_460),
.C(n_463),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_494),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_503),
.A2(n_505),
.B1(n_508),
.B2(n_509),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_473),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_491),
.B(n_469),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_494),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_496),
.B(n_479),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_462),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_514),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_501),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_504),
.B(n_477),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_516),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_502),
.B(n_471),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_506),
.B(n_493),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_517),
.B(n_521),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_500),
.B(n_465),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_511),
.B(n_488),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_522),
.B(n_504),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_499),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_524),
.B(n_527),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_520),
.B(n_507),
.C(n_492),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_529),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_515),
.A2(n_489),
.B(n_485),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_519),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_530),
.B(n_523),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_519),
.C(n_514),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_524),
.Y(n_535)
);

OAI21xp33_ASAP7_75t_SL g536 ( 
.A1(n_534),
.A2(n_535),
.B(n_532),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_536),
.B(n_537),
.C(n_530),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_535),
.B(n_513),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_533),
.B(n_510),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_485),
.B1(n_510),
.B2(n_484),
.Y(n_540)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_540),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_495),
.B(n_497),
.Y(n_542)
);


endmodule