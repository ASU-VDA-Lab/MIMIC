module fake_ariane_116_n_4974 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_4974);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_4974;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_2182;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_3765;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_2042;
wire n_1131;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_625;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_559;
wire n_4824;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_561;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_786;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_3482;
wire n_823;
wire n_1900;
wire n_620;
wire n_4268;
wire n_587;
wire n_863;
wire n_3960;
wire n_2433;
wire n_899;
wire n_3975;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_661;
wire n_4227;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_4476;
wire n_579;
wire n_844;
wire n_1267;
wire n_2956;
wire n_2382;
wire n_1213;
wire n_780;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_570;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_575;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3841;
wire n_851;
wire n_3900;
wire n_3413;
wire n_3539;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_555;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_992;
wire n_966;
wire n_3549;
wire n_3914;
wire n_1692;
wire n_2611;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_1178;
wire n_2015;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_619;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_542;
wire n_1087;
wire n_632;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_4367;
wire n_2467;
wire n_4195;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_4254;
wire n_646;
wire n_3438;
wire n_2625;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_670;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_1032;
wire n_1592;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_4588;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_4153;
wire n_1868;
wire n_3601;
wire n_2373;
wire n_3881;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_604;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_4247;
wire n_707;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_688;
wire n_636;
wire n_1490;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_887;
wire n_2125;
wire n_1156;
wire n_2861;
wire n_4344;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_4313;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_4798;
wire n_1500;
wire n_616;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_3337;
wire n_1189;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_655;
wire n_4237;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_951;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_704;
wire n_2958;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_3340;
wire n_1243;
wire n_3486;
wire n_608;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_811;
wire n_791;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_642;
wire n_1406;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_3740;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_1256;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_4882;
wire n_3206;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_3987;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_3380;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_4685;
wire n_565;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_2963;
wire n_2561;
wire n_1056;
wire n_674;
wire n_3168;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_4922;
wire n_629;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_724;
wire n_2931;
wire n_3433;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_875;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_3645;
wire n_793;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_1554;
wire n_3279;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_581;
wire n_3091;
wire n_1024;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_549;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_3633;
wire n_857;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1064;
wire n_633;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_1141;
wire n_3457;
wire n_2324;
wire n_840;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_614;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_2290;
wire n_4398;
wire n_2856;
wire n_3235;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_3628;
wire n_4777;
wire n_3941;
wire n_1915;
wire n_658;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_860;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_774;
wire n_1168;
wire n_4663;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_656;
wire n_4963;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_1581;
wire n_946;
wire n_3058;
wire n_757;
wire n_2047;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_998;
wire n_3592;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_1339;
wire n_1051;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_4622;
wire n_4757;
wire n_1871;
wire n_803;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_548;
wire n_3427;
wire n_3162;
wire n_4591;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_2259;
wire n_849;
wire n_4655;
wire n_1820;
wire n_1233;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_675;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_1169;
wire n_789;
wire n_3181;
wire n_1916;
wire n_610;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_4416;
wire n_4439;
wire n_870;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_645;
wire n_721;
wire n_1084;
wire n_1276;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_3474;
wire n_2458;
wire n_3150;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_4031;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_612;
wire n_4680;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_546;
wire n_1159;
wire n_4498;
wire n_772;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_652;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_3391;
wire n_912;
wire n_4786;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_3240;
wire n_931;
wire n_3362;
wire n_4130;
wire n_967;
wire n_4175;
wire n_1079;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_1226;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_3515;
wire n_2363;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_564;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_552;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_4275;
wire n_3774;
wire n_926;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_855;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_3508;
wire n_4129;
wire n_1105;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_4677;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_2008;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1747;
wire n_3990;
wire n_1171;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_1400;
wire n_3735;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_2137;
wire n_3685;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_595;
wire n_1405;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_1557;
wire n_4744;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_4835;
wire n_1151;
wire n_554;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4559;
wire n_4742;
wire n_3566;
wire n_1133;
wire n_883;
wire n_4372;
wire n_4097;
wire n_4162;
wire n_779;
wire n_4790;
wire n_594;
wire n_4173;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_3738;
wire n_894;
wire n_1380;
wire n_562;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_1023;
wire n_914;
wire n_689;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_588;
wire n_638;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_617;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_2592;
wire n_3490;
wire n_962;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_1968;
wire n_918;
wire n_639;
wire n_673;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_4333;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_2236;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_622;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_1221;
wire n_4217;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_1204;
wire n_994;
wire n_2428;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_856;
wire n_4592;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_679;
wire n_3047;
wire n_3163;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_607;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_4933;
wire n_968;
wire n_4144;
wire n_3278;
wire n_2375;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_1755;
wire n_2212;
wire n_4434;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_831;
wire n_3681;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_550;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_671;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_684;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_4232;
wire n_2097;
wire n_662;
wire n_3461;
wire n_1410;
wire n_2297;
wire n_939;
wire n_4203;
wire n_1325;
wire n_1223;
wire n_2957;
wire n_572;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_3763;
wire n_933;
wire n_3499;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_3590;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_626;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_1264;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_573;
wire n_2823;
wire n_3684;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_589;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_603;
wire n_4259;
wire n_2030;
wire n_850;
wire n_4299;
wire n_2407;
wire n_690;
wire n_2243;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_2731;
wire n_3703;
wire n_1246;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_1196;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_1187;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_568;
wire n_4796;
wire n_1088;
wire n_766;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_665;
wire n_4625;
wire n_2107;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_672;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_3856;
wire n_4038;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_557;
wire n_3419;
wire n_989;
wire n_2233;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_1514;
wire n_2782;
wire n_569;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_4488;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_611;
wire n_2060;
wire n_1295;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_1112;
wire n_700;
wire n_4174;
wire n_2145;
wire n_4801;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_577;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_1253;
wire n_1468;
wire n_762;
wire n_4378;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_2072;
wire n_3852;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_563;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_2762;
wire n_964;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_2261;
wire n_3082;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_1095;
wire n_3078;
wire n_3971;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_3171;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_2308;
wire n_1939;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_547;
wire n_677;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_3788;
wire n_3939;
wire n_590;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_545;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_627;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_3579;
wire n_2379;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_4551;
wire n_551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_1239;
wire n_3417;
wire n_560;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_4328;
wire n_1854;
wire n_666;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1394;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_1078;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_618;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_4766;
wire n_592;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_640;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_643;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_1441;
wire n_682;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_686;
wire n_1154;
wire n_584;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_3976;
wire n_2813;
wire n_2546;
wire n_3381;
wire n_897;
wire n_3736;
wire n_4466;
wire n_891;
wire n_1659;
wire n_3955;
wire n_885;
wire n_1864;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_714;
wire n_3605;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_3840;
wire n_2198;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_2133;
wire n_2497;
wire n_879;
wire n_4561;
wire n_1541;
wire n_597;
wire n_3291;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_1116;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_1549;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_2692;
wire n_683;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_2553;
wire n_1420;
wire n_2645;
wire n_4711;
wire n_2749;
wire n_660;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_571;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_613;
wire n_1022;
wire n_3532;
wire n_2609;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_621;
wire n_1772;
wire n_3106;
wire n_1311;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_697;
wire n_4620;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_880;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_975;
wire n_1645;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_2465;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_4858;
wire n_1445;
wire n_4435;
wire n_3248;
wire n_2387;
wire n_4318;
wire n_830;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_4673;
wire n_2793;
wire n_541;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_663;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2597;
wire n_1077;
wire n_2321;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_1271;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_900;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_2039;
wire n_1285;
wire n_761;
wire n_733;
wire n_3838;
wire n_4059;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_648;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_654;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_539;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_1393;
wire n_723;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_4886;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1982;
wire n_641;
wire n_910;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_4693;
wire n_1043;
wire n_4956;
wire n_2869;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_3112;
wire n_954;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_664;
wire n_1591;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_3779;
wire n_599;
wire n_537;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_583;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_3986;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_1252;
wire n_3045;
wire n_773;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_2135;
wire n_4475;
wire n_1463;
wire n_4626;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_634;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_4702;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_1314;
wire n_1512;
wire n_884;
wire n_3324;
wire n_2192;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_4768;
wire n_1889;
wire n_693;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2769;
wire n_1548;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_2727;
wire n_942;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_3562;
wire n_2281;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_1819;
wire n_3095;
wire n_947;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_1442;
wire n_696;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2549;
wire n_2499;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_4794;
wire n_4843;
wire n_669;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_2462;
wire n_2155;
wire n_615;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_824;
wire n_4272;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_815;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_1627;
wire n_2903;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_965;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_713;
wire n_3179;
wire n_598;
wire n_4836;
wire n_3889;
wire n_3262;
wire n_927;
wire n_3699;
wire n_706;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_3276;
wire n_3682;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_553;
wire n_814;
wire n_578;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_647;
wire n_2027;
wire n_2932;
wire n_600;
wire n_3118;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_1467;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_681;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_920;
wire n_3951;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_861;
wire n_1666;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_3648;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_657;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_1532;
wire n_1030;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_4145;
wire n_624;
wire n_876;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_854;
wire n_2091;
wire n_4312;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_3694;
wire n_771;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_586;
wire n_3543;
wire n_1324;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_605;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_2698;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_3907;
wire n_4603;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_4595;
wire n_960;
wire n_2352;
wire n_790;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_1426;
wire n_4969;
wire n_4641;
wire n_4399;
wire n_4140;
wire n_566;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_4450;
wire n_2934;
wire n_576;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_623;
wire n_3509;
wire n_1403;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_543;
wire n_3456;
wire n_4532;
wire n_601;
wire n_628;
wire n_3790;
wire n_907;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_3101;
wire n_3662;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_593;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_609;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_3533;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_1157;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_540;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_1100;
wire n_585;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_580;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_3470;
wire n_1407;
wire n_2865;
wire n_973;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_3269;
wire n_558;
wire n_4231;
wire n_2591;
wire n_653;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_2550;
wire n_556;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_2169;
wire n_591;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_668;
wire n_2111;
wire n_3743;
wire n_2948;
wire n_3099;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_1003;
wire n_701;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_694;
wire n_4749;
wire n_1845;
wire n_921;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_630;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_741;
wire n_2964;
wire n_865;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_902;
wire n_1723;
wire n_3918;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_596;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_574;
wire n_3593;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_2081;
wire n_1474;
wire n_937;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_1249;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;

INVx1_ASAP7_75t_L g537 ( 
.A(n_175),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_436),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_287),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_109),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_464),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_154),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_26),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_46),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_330),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_360),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_183),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_323),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_327),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_535),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_120),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_227),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_198),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_281),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_216),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_105),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_433),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_475),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_440),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_492),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_412),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_506),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_510),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_67),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_350),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_341),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_457),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_507),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_206),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_382),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_181),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_193),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_238),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_130),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_47),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_183),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_179),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_13),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_502),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_474),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_95),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_301),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_467),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_153),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_471),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_470),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_118),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_392),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_8),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_514),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_104),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_18),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_369),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_25),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_266),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_477),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_488),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_122),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_55),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_288),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_39),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_419),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_186),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_40),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_432),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_348),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_468),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_347),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_528),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_456),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_108),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_182),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_435),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_125),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_523),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_224),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_149),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_111),
.Y(n_619)
);

INVx4_ASAP7_75t_R g620 ( 
.A(n_132),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_495),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_414),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_450),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_465),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_185),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_131),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_305),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_503),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_458),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_479),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_126),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_530),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_353),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_48),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_497),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_330),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_434),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_498),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_352),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_513),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_136),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_454),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_500),
.Y(n_643)
);

CKINVDCx14_ASAP7_75t_R g644 ( 
.A(n_512),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_314),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_136),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_229),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_162),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_483),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_505),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_11),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_15),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_484),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_302),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_194),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_61),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_306),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_532),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_281),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_408),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_158),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_19),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_473),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_104),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_354),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_204),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_189),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_225),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_10),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_231),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_153),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_145),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_302),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_525),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_453),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_66),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_165),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_515),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_352),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_360),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_339),
.Y(n_681)
);

CKINVDCx16_ASAP7_75t_R g682 ( 
.A(n_293),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_184),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_324),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_324),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_129),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_277),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_519),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_124),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_284),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_442),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_40),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_372),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_127),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_364),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_194),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_8),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_485),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_3),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_224),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_160),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_370),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_174),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_348),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_235),
.Y(n_705)
);

CKINVDCx16_ASAP7_75t_R g706 ( 
.A(n_108),
.Y(n_706)
);

CKINVDCx16_ASAP7_75t_R g707 ( 
.A(n_241),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_131),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_162),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_417),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_388),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_460),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_501),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_69),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_381),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_61),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_316),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_127),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_373),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_490),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_280),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_223),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_284),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_289),
.Y(n_724)
);

BUFx2_ASAP7_75t_SL g725 ( 
.A(n_439),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_25),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_240),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_421),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_271),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_232),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_345),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_518),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_378),
.Y(n_733)
);

CKINVDCx16_ASAP7_75t_R g734 ( 
.A(n_466),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_389),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_315),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_58),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_132),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_402),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_249),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_459),
.Y(n_741)
);

BUFx10_ASAP7_75t_L g742 ( 
.A(n_504),
.Y(n_742)
);

CKINVDCx16_ASAP7_75t_R g743 ( 
.A(n_51),
.Y(n_743)
);

BUFx5_ASAP7_75t_L g744 ( 
.A(n_219),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_372),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_260),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_13),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_365),
.Y(n_748)
);

BUFx10_ASAP7_75t_L g749 ( 
.A(n_431),
.Y(n_749)
);

CKINVDCx16_ASAP7_75t_R g750 ( 
.A(n_332),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_349),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_202),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_252),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_487),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_494),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_489),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_203),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_272),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_142),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_524),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_18),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_48),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_337),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_393),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_161),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_496),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_20),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_53),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_10),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_516),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_311),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_91),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_216),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_112),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_42),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_316),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_247),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_422),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_137),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_57),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_118),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_280),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_298),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_461),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_314),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_511),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_399),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_133),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_405),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_391),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_199),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_430),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_86),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_96),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_200),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_20),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_437),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_213),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_290),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_296),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_12),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_298),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_452),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_57),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_325),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_317),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_320),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_154),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_188),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_446),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_120),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_5),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_177),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_182),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_227),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_113),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_493),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_167),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_169),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_24),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_526),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_168),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_520),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_74),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_476),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_373),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_337),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_534),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_139),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_70),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_177),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_531),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_277),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_30),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_110),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_130),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_294),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_323),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_117),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_259),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_133),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_329),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_527),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_521),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_386),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_286),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_359),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_79),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_486),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_283),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_210),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_259),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_33),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_197),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_304),
.Y(n_855)
);

BUFx10_ASAP7_75t_L g856 ( 
.A(n_533),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_60),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_261),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_305),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_258),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_112),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_398),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_383),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_155),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_343),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_426),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_335),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_399),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_370),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_404),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_126),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_100),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_217),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_135),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_438),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_169),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_200),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_58),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_536),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_89),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_408),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_478),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_340),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_94),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_522),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_282),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_141),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_258),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_400),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_394),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_237),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_220),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_32),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_386),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_444),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_205),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_232),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_449),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_411),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_233),
.Y(n_900)
);

CKINVDCx16_ASAP7_75t_R g901 ( 
.A(n_220),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_250),
.Y(n_902)
);

CKINVDCx16_ASAP7_75t_R g903 ( 
.A(n_443),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_413),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_147),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_210),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_203),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_164),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_391),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_38),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_310),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_248),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_413),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_482),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_225),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_174),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_462),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_441),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_144),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_135),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_179),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_429),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_229),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_14),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_371),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_185),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_172),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_366),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_455),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_509),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_77),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_418),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_451),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_215),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_82),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_171),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_66),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_423),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_180),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_508),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_160),
.Y(n_941)
);

BUFx8_ASAP7_75t_SL g942 ( 
.A(n_187),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_269),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_15),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_151),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_178),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_152),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_529),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_41),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_3),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_77),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_134),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_115),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_268),
.Y(n_954)
);

BUFx5_ASAP7_75t_L g955 ( 
.A(n_252),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_152),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_491),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_223),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_218),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_377),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_103),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_481),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_463),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_44),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_499),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_299),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_206),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_390),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_517),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_472),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_400),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_469),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_56),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_251),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_17),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_411),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_238),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_80),
.Y(n_978)
);

BUFx10_ASAP7_75t_L g979 ( 
.A(n_164),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_143),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_6),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_380),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_744),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_609),
.Y(n_984)
);

INVxp33_ASAP7_75t_L g985 ( 
.A(n_718),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_609),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_734),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_609),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_744),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_695),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_695),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_734),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_695),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_700),
.Y(n_994)
);

INVxp67_ASAP7_75t_SL g995 ( 
.A(n_700),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_700),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_722),
.Y(n_997)
);

INVxp33_ASAP7_75t_L g998 ( 
.A(n_942),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_744),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_903),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_963),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_722),
.Y(n_1002)
);

INVxp67_ASAP7_75t_SL g1003 ( 
.A(n_722),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_822),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_822),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_903),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_822),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_560),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_826),
.Y(n_1009)
);

NOR2xp67_ASAP7_75t_L g1010 ( 
.A(n_588),
.B(n_0),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_826),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_560),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_574),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_574),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_826),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_591),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_835),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_835),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_835),
.Y(n_1019)
);

CKINVDCx16_ASAP7_75t_R g1020 ( 
.A(n_682),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_839),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_744),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_839),
.Y(n_1023)
);

CKINVDCx16_ASAP7_75t_R g1024 ( 
.A(n_682),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_839),
.Y(n_1025)
);

BUFx2_ASAP7_75t_SL g1026 ( 
.A(n_675),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_883),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_591),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_744),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_883),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_883),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_935),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_935),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_744),
.Y(n_1034)
);

CKINVDCx16_ASAP7_75t_R g1035 ( 
.A(n_706),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_935),
.Y(n_1036)
);

CKINVDCx14_ASAP7_75t_R g1037 ( 
.A(n_644),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_960),
.Y(n_1038)
);

INVxp67_ASAP7_75t_SL g1039 ( 
.A(n_960),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_756),
.Y(n_1040)
);

INVxp67_ASAP7_75t_SL g1041 ( 
.A(n_960),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_745),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_567),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_756),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_744),
.Y(n_1045)
);

INVxp33_ASAP7_75t_L g1046 ( 
.A(n_874),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_567),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_706),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_567),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_744),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_797),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_797),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_576),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_675),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_707),
.Y(n_1055)
);

INVxp33_ASAP7_75t_SL g1056 ( 
.A(n_874),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_576),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_588),
.B(n_593),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_576),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_707),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_601),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_601),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_743),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_601),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_679),
.Y(n_1065)
);

CKINVDCx16_ASAP7_75t_R g1066 ( 
.A(n_743),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_679),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_675),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_679),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_675),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_724),
.Y(n_1071)
);

INVxp33_ASAP7_75t_L g1072 ( 
.A(n_537),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_724),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_724),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_747),
.Y(n_1075)
);

CKINVDCx14_ASAP7_75t_R g1076 ( 
.A(n_742),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_742),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_848),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_848),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_848),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_744),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_742),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_747),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_955),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_955),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_955),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_750),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_742),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_955),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_955),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_955),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_876),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_955),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_955),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_955),
.Y(n_1095)
);

CKINVDCx16_ASAP7_75t_R g1096 ( 
.A(n_750),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_553),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_749),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_553),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_876),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_564),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_749),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_547),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_749),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_876),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_654),
.Y(n_1106)
);

INVxp33_ASAP7_75t_SL g1107 ( 
.A(n_539),
.Y(n_1107)
);

INVxp67_ASAP7_75t_SL g1108 ( 
.A(n_900),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_540),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_749),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_900),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_900),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_953),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_953),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_953),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_961),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_961),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_961),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_537),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_982),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_982),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_544),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_901),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_544),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_963),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_963),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_810),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_549),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_810),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_540),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_540),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_540),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_549),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_565),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_565),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_572),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_572),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_564),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_589),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_810),
.Y(n_1140)
);

CKINVDCx16_ASAP7_75t_R g1141 ( 
.A(n_901),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_589),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_590),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_810),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_856),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_542),
.Y(n_1146)
);

INVxp33_ASAP7_75t_L g1147 ( 
.A(n_590),
.Y(n_1147)
);

CKINVDCx14_ASAP7_75t_R g1148 ( 
.A(n_856),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_594),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_594),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_856),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_657),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_595),
.Y(n_1153)
);

CKINVDCx14_ASAP7_75t_R g1154 ( 
.A(n_856),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_621),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_564),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_629),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_895),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_970),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_595),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_543),
.Y(n_1161)
);

BUFx2_ASAP7_75t_SL g1162 ( 
.A(n_638),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_596),
.Y(n_1163)
);

BUFx2_ASAP7_75t_SL g1164 ( 
.A(n_638),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_596),
.Y(n_1165)
);

INVxp33_ASAP7_75t_L g1166 ( 
.A(n_602),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_602),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_618),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_618),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_619),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_619),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_626),
.Y(n_1172)
);

BUFx2_ASAP7_75t_SL g1173 ( 
.A(n_638),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_626),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_546),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_548),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_633),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_633),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_634),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_559),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_540),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_634),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_639),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_716),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_639),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_647),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_647),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_662),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_551),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_662),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_665),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_665),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_540),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_667),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_545),
.B(n_562),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_667),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_668),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_552),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_668),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_554),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_559),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_669),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_669),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_555),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_556),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_672),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_570),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_571),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_759),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_573),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_672),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_673),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_790),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_772),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_785),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_673),
.Y(n_1216)
);

INVxp67_ASAP7_75t_SL g1217 ( 
.A(n_790),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_677),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_790),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_790),
.Y(n_1220)
);

INVxp33_ASAP7_75t_SL g1221 ( 
.A(n_575),
.Y(n_1221)
);

INVxp33_ASAP7_75t_L g1222 ( 
.A(n_677),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_584),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_577),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_680),
.Y(n_1225)
);

CKINVDCx16_ASAP7_75t_R g1226 ( 
.A(n_745),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_790),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_963),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_680),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_795),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_578),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_684),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_579),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_582),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_583),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_585),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_684),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_690),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_690),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_693),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_693),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_790),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_811),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_702),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_702),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_704),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_704),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_705),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_830),
.Y(n_1249)
);

CKINVDCx16_ASAP7_75t_R g1250 ( 
.A(n_745),
.Y(n_1250)
);

INVxp33_ASAP7_75t_SL g1251 ( 
.A(n_592),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_599),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_600),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_705),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_709),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_709),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_796),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_796),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_604),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_796),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_710),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_605),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_710),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_584),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_719),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_607),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_719),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_726),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_612),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_608),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_796),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_726),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_727),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_613),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_796),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_727),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_615),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_796),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_608),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_630),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_617),
.Y(n_1281)
);

INVxp67_ASAP7_75t_L g1282 ( 
.A(n_731),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_622),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_731),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_736),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_736),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_593),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_739),
.Y(n_1288)
);

CKINVDCx16_ASAP7_75t_R g1289 ( 
.A(n_745),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_963),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_739),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_740),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_740),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_746),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_746),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_761),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_761),
.Y(n_1297)
);

NOR2xp67_ASAP7_75t_L g1298 ( 
.A(n_681),
.B(n_0),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_630),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_765),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_765),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_767),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_625),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_767),
.Y(n_1304)
);

CKINVDCx16_ASAP7_75t_R g1305 ( 
.A(n_884),
.Y(n_1305)
);

NOR2xp67_ASAP7_75t_L g1306 ( 
.A(n_681),
.B(n_1),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_627),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_779),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_631),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_779),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_781),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_635),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_781),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_782),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_636),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_641),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_645),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_782),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_783),
.Y(n_1319)
);

INVxp33_ASAP7_75t_SL g1320 ( 
.A(n_646),
.Y(n_1320)
);

INVxp33_ASAP7_75t_L g1321 ( 
.A(n_783),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_789),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_789),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_798),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_798),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_648),
.Y(n_1326)
);

INVxp33_ASAP7_75t_SL g1327 ( 
.A(n_652),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_816),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_816),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_819),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_635),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_819),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_640),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_640),
.Y(n_1334)
);

CKINVDCx16_ASAP7_75t_R g1335 ( 
.A(n_884),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_642),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_827),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_833),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_827),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_829),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_655),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_829),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_836),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_836),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_642),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_656),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_659),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_660),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_841),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_913),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_841),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_649),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_661),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_842),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_664),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_666),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_923),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_842),
.Y(n_1358)
);

CKINVDCx16_ASAP7_75t_R g1359 ( 
.A(n_884),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_845),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_845),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_649),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_670),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_946),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1061),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1155),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_1152),
.Y(n_1367)
);

INVxp67_ASAP7_75t_SL g1368 ( 
.A(n_1101),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1069),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1026),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1155),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1092),
.Y(n_1372)
);

CKINVDCx14_ASAP7_75t_R g1373 ( 
.A(n_1076),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1101),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1157),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1152),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1100),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1157),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_1184),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1158),
.Y(n_1380)
);

CKINVDCx16_ASAP7_75t_R g1381 ( 
.A(n_1226),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1108),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1184),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_984),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1209),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1158),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1209),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_986),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1148),
.B(n_658),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_988),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_1054),
.B(n_638),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_990),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1215),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1026),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1215),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_991),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1109),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_993),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1138),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1103),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1159),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_994),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1230),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1159),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1106),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_1138),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_1230),
.Y(n_1407)
);

INVxp33_ASAP7_75t_SL g1408 ( 
.A(n_987),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_996),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1214),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1243),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1054),
.B(n_658),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1243),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_1156),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1109),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1020),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1338),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1037),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_997),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1338),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1002),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1154),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1350),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1156),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1004),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1005),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1048),
.Y(n_1427)
);

CKINVDCx20_ASAP7_75t_R g1428 ( 
.A(n_1350),
.Y(n_1428)
);

INVxp33_ASAP7_75t_L g1429 ( 
.A(n_1060),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_987),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1299),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1357),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1249),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1007),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1009),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1011),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1015),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1017),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1068),
.B(n_691),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1018),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1357),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1048),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1019),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1021),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1364),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1175),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1023),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1025),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1217),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1175),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1176),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_995),
.B(n_691),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1176),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1189),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_992),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1027),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1030),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1189),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1198),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1198),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1055),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1031),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_992),
.Y(n_1463)
);

NOR2xp67_ASAP7_75t_L g1464 ( 
.A(n_1068),
.B(n_538),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1024),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1070),
.B(n_728),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1200),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1032),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1200),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1055),
.Y(n_1470)
);

CKINVDCx20_ASAP7_75t_R g1471 ( 
.A(n_1063),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1063),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1205),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1033),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1087),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1036),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1038),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1227),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1271),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1205),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1081),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1278),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1087),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1097),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1123),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1097),
.Y(n_1486)
);

CKINVDCx20_ASAP7_75t_R g1487 ( 
.A(n_1123),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1035),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1000),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1208),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1099),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1099),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1279),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1279),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1280),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1130),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1280),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1003),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1333),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1039),
.B(n_1041),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1070),
.B(n_728),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1208),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1066),
.Y(n_1503)
);

CKINVDCx16_ASAP7_75t_R g1504 ( 
.A(n_1250),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1333),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1130),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1096),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1141),
.Y(n_1508)
);

NOR2xp67_ASAP7_75t_L g1509 ( 
.A(n_1077),
.B(n_541),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1210),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1334),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1334),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1336),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1210),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1289),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1075),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1075),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1305),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1336),
.Y(n_1519)
);

INVxp67_ASAP7_75t_SL g1520 ( 
.A(n_1180),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1083),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1119),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1224),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1224),
.Y(n_1524)
);

CKINVDCx16_ASAP7_75t_R g1525 ( 
.A(n_1335),
.Y(n_1525)
);

NOR2xp67_ASAP7_75t_L g1526 ( 
.A(n_1077),
.B(n_550),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1231),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1120),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1231),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1233),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1233),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1081),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1121),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_L g1534 ( 
.A(n_1082),
.B(n_558),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1083),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1122),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1234),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1124),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1162),
.B(n_741),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1359),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1234),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1128),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1133),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1235),
.Y(n_1544)
);

NOR2xp67_ASAP7_75t_L g1545 ( 
.A(n_1082),
.B(n_561),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1134),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1235),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1135),
.Y(n_1548)
);

INVxp67_ASAP7_75t_SL g1549 ( 
.A(n_1180),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1236),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1236),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_SL g1552 ( 
.A(n_1042),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1088),
.B(n_741),
.Y(n_1553)
);

CKINVDCx14_ASAP7_75t_R g1554 ( 
.A(n_1000),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_R g1555 ( 
.A(n_1088),
.B(n_563),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1252),
.Y(n_1556)
);

NOR2xp67_ASAP7_75t_L g1557 ( 
.A(n_1098),
.B(n_568),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1136),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1131),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_R g1560 ( 
.A(n_1098),
.B(n_580),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1201),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1252),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1137),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1139),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1253),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1146),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1142),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1006),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1253),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1143),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1161),
.Y(n_1571)
);

CKINVDCx14_ASAP7_75t_R g1572 ( 
.A(n_1006),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1149),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1150),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1259),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1153),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1162),
.B(n_817),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1259),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1262),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1262),
.Y(n_1580)
);

CKINVDCx14_ASAP7_75t_R g1581 ( 
.A(n_1102),
.Y(n_1581)
);

CKINVDCx20_ASAP7_75t_R g1582 ( 
.A(n_1266),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1160),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1163),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1201),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1266),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1269),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1269),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1165),
.Y(n_1589)
);

CKINVDCx20_ASAP7_75t_R g1590 ( 
.A(n_1274),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1223),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1167),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1168),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1169),
.Y(n_1594)
);

CKINVDCx20_ASAP7_75t_R g1595 ( 
.A(n_1274),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1170),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1277),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1171),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1102),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1104),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1104),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1277),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_1281),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1172),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1281),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1110),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1223),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1174),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1177),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1178),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1283),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1264),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1110),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1283),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1182),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1307),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1307),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1183),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1264),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1185),
.Y(n_1620)
);

INVxp67_ASAP7_75t_SL g1621 ( 
.A(n_1270),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1309),
.Y(n_1622)
);

CKINVDCx16_ASAP7_75t_R g1623 ( 
.A(n_1204),
.Y(n_1623)
);

CKINVDCx16_ASAP7_75t_R g1624 ( 
.A(n_1207),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1186),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1187),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1309),
.Y(n_1627)
);

INVxp67_ASAP7_75t_SL g1628 ( 
.A(n_1270),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1188),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1190),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1191),
.Y(n_1631)
);

CKINVDCx16_ASAP7_75t_R g1632 ( 
.A(n_1303),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1315),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1315),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1316),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1192),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1316),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1194),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1317),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1317),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1196),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1131),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1326),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1127),
.B(n_1129),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1326),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1197),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1199),
.Y(n_1647)
);

CKINVDCx20_ASAP7_75t_R g1648 ( 
.A(n_1341),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1341),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1203),
.Y(n_1650)
);

BUFx2_ASAP7_75t_SL g1651 ( 
.A(n_1058),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1346),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1206),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_1346),
.Y(n_1654)
);

INVxp67_ASAP7_75t_SL g1655 ( 
.A(n_1362),
.Y(n_1655)
);

NOR2xp67_ASAP7_75t_L g1656 ( 
.A(n_1127),
.B(n_587),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1164),
.B(n_817),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1211),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_1347),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1347),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1348),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1348),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1216),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1225),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1229),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1353),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1353),
.Y(n_1667)
);

CKINVDCx14_ASAP7_75t_R g1668 ( 
.A(n_1129),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1140),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1355),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1232),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1237),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1140),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1238),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1239),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1355),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1240),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_1356),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1241),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1356),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1244),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1363),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1245),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1246),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1247),
.Y(n_1685)
);

INVxp67_ASAP7_75t_SL g1686 ( 
.A(n_1362),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1449),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1397),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1397),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1400),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1415),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1481),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1415),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1484),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1481),
.Y(n_1695)
);

CKINVDCx20_ASAP7_75t_R g1696 ( 
.A(n_1367),
.Y(n_1696)
);

NOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1464),
.B(n_1287),
.Y(n_1697)
);

INVx4_ASAP7_75t_L g1698 ( 
.A(n_1532),
.Y(n_1698)
);

BUFx8_ASAP7_75t_L g1699 ( 
.A(n_1427),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1520),
.B(n_1042),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1517),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1496),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1486),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1496),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1491),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1532),
.Y(n_1706)
);

CKINVDCx20_ASAP7_75t_R g1707 ( 
.A(n_1367),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1509),
.B(n_1287),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1412),
.A2(n_1012),
.B1(n_1016),
.B2(n_1008),
.Y(n_1709)
);

INVx6_ASAP7_75t_L g1710 ( 
.A(n_1447),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1492),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1493),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1506),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1494),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1549),
.B(n_1072),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1561),
.B(n_1147),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1585),
.B(n_1144),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1506),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1495),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1497),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1559),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1499),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1505),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1591),
.B(n_1166),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1422),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1511),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1607),
.B(n_1179),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1422),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1559),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1642),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1431),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1612),
.B(n_1144),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1642),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1619),
.B(n_1354),
.Y(n_1734)
);

INVx5_ASAP7_75t_L g1735 ( 
.A(n_1431),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1512),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1621),
.B(n_1145),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1513),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1431),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1447),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1628),
.B(n_1202),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1370),
.B(n_1107),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1519),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1581),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1384),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1522),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1478),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1655),
.B(n_1222),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1479),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1686),
.B(n_1321),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1482),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1528),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1388),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1390),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1368),
.B(n_1212),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1392),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1498),
.B(n_1046),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1533),
.B(n_1536),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1396),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1668),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1439),
.B(n_1145),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1398),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1374),
.B(n_1218),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1402),
.Y(n_1764)
);

BUFx8_ASAP7_75t_L g1765 ( 
.A(n_1605),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1409),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1538),
.B(n_985),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1373),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1419),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1542),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1421),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1425),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1426),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1434),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1435),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1436),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1437),
.Y(n_1777)
);

BUFx3_ASAP7_75t_L g1778 ( 
.A(n_1438),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1466),
.B(n_1151),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1543),
.B(n_1299),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1399),
.B(n_1282),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1546),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1548),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1371),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1488),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1440),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1558),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1406),
.B(n_1286),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1443),
.Y(n_1789)
);

CKINVDCx20_ASAP7_75t_R g1790 ( 
.A(n_1376),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1563),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1444),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1564),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1375),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1378),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1567),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1570),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1416),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_R g1799 ( 
.A(n_1554),
.B(n_1151),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_1376),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1573),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1574),
.B(n_1312),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1576),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_1379),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1448),
.Y(n_1805)
);

BUFx2_ASAP7_75t_L g1806 ( 
.A(n_1488),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1405),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1583),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1456),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1503),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1457),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1584),
.Y(n_1812)
);

AND2x6_ASAP7_75t_L g1813 ( 
.A(n_1389),
.B(n_569),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1462),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1468),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1589),
.B(n_1312),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1501),
.B(n_1107),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1592),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1593),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1553),
.B(n_1164),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1594),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1474),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1503),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1596),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1476),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1477),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1598),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1604),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1608),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1465),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1394),
.B(n_1221),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1414),
.B(n_1173),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1609),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1516),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1424),
.B(n_1391),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1521),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1539),
.B(n_1173),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1610),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1644),
.B(n_1221),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1615),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1618),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1577),
.B(n_1008),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1620),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1625),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1626),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1552),
.A2(n_1012),
.B1(n_1028),
.B2(n_1016),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1365),
.B(n_1010),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1629),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1630),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_R g1850 ( 
.A(n_1572),
.B(n_1363),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1410),
.Y(n_1851)
);

CKINVDCx20_ASAP7_75t_R g1852 ( 
.A(n_1379),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1380),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_1685),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1631),
.Y(n_1855)
);

CKINVDCx20_ASAP7_75t_R g1856 ( 
.A(n_1383),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1369),
.B(n_1298),
.Y(n_1857)
);

BUFx6f_ASAP7_75t_L g1858 ( 
.A(n_1636),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1386),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1638),
.B(n_1331),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1641),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1646),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1647),
.Y(n_1863)
);

BUFx2_ASAP7_75t_L g1864 ( 
.A(n_1507),
.Y(n_1864)
);

BUFx2_ASAP7_75t_L g1865 ( 
.A(n_1507),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1433),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1650),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1653),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1658),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1663),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1664),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_SL g1872 ( 
.A(n_1418),
.B(n_1056),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1665),
.B(n_1331),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1671),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1672),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1535),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1674),
.B(n_1345),
.Y(n_1877)
);

INVxp67_ASAP7_75t_L g1878 ( 
.A(n_1445),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1401),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1675),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1684),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1677),
.B(n_1345),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1657),
.B(n_1028),
.Y(n_1883)
);

BUFx8_ASAP7_75t_L g1884 ( 
.A(n_1634),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1651),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1679),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1681),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1683),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1372),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1500),
.B(n_1040),
.Y(n_1890)
);

INVx6_ASAP7_75t_L g1891 ( 
.A(n_1381),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1377),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1404),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1382),
.B(n_1452),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1526),
.B(n_1040),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1508),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1418),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1552),
.B(n_1251),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1442),
.A2(n_1470),
.B1(n_1471),
.B2(n_1461),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1552),
.Y(n_1900)
);

INVx3_ASAP7_75t_L g1901 ( 
.A(n_1446),
.Y(n_1901)
);

XOR2xp5_ASAP7_75t_L g1902 ( 
.A(n_1578),
.B(n_998),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1534),
.B(n_1044),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1450),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1545),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1557),
.B(n_1044),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1566),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1366),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1656),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_1366),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1555),
.B(n_1251),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1571),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1602),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1662),
.Y(n_1914)
);

AND2x6_ASAP7_75t_L g1915 ( 
.A(n_1455),
.B(n_569),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1451),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1463),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1453),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1454),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1458),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1459),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1460),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1560),
.B(n_1051),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1467),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1599),
.B(n_1051),
.Y(n_1925)
);

BUFx8_ASAP7_75t_L g1926 ( 
.A(n_1508),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1469),
.B(n_1306),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1473),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1480),
.B(n_1330),
.Y(n_1929)
);

CKINVDCx20_ASAP7_75t_R g1930 ( 
.A(n_1383),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1490),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1502),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1510),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1514),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1523),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1599),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1600),
.Y(n_1937)
);

NAND2xp33_ASAP7_75t_R g1938 ( 
.A(n_1430),
.B(n_1056),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1524),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1429),
.B(n_1352),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1600),
.A2(n_1052),
.B1(n_1327),
.B2(n_1320),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1527),
.Y(n_1942)
);

INVx3_ASAP7_75t_L g1943 ( 
.A(n_1529),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1601),
.B(n_1352),
.Y(n_1944)
);

INVx5_ASAP7_75t_L g1945 ( 
.A(n_1504),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1530),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1531),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1537),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1601),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1541),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1544),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1547),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1606),
.B(n_1052),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1606),
.B(n_1613),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1613),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1550),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1408),
.B(n_1320),
.Y(n_1957)
);

NAND2x1p5_ASAP7_75t_L g1958 ( 
.A(n_1408),
.B(n_1195),
.Y(n_1958)
);

CKINVDCx14_ASAP7_75t_R g1959 ( 
.A(n_1669),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1551),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1556),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1562),
.Y(n_1962)
);

AND2x2_ASAP7_75t_SL g1963 ( 
.A(n_1525),
.B(n_569),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1669),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1673),
.B(n_1248),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1565),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1569),
.B(n_1254),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1673),
.B(n_1327),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1575),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1580),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1587),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1588),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1597),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_1385),
.Y(n_1974)
);

NOR2x1_ASAP7_75t_L g1975 ( 
.A(n_1578),
.B(n_1195),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1617),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1622),
.B(n_1351),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1627),
.Y(n_1978)
);

INVxp67_ASAP7_75t_L g1979 ( 
.A(n_1633),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1635),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1639),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1640),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1643),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1645),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1623),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1624),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1649),
.B(n_828),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1652),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1661),
.B(n_1255),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1666),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1667),
.B(n_1085),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1676),
.B(n_1013),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1682),
.B(n_1256),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1430),
.B(n_1261),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1489),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1632),
.Y(n_1996)
);

CKINVDCx16_ASAP7_75t_R g1997 ( 
.A(n_1579),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1489),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1579),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_R g2000 ( 
.A(n_1515),
.B(n_597),
.Y(n_2000)
);

OA21x2_ASAP7_75t_L g2001 ( 
.A1(n_1568),
.A2(n_1086),
.B(n_1085),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1582),
.Y(n_2002)
);

BUFx3_ASAP7_75t_L g2003 ( 
.A(n_1582),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1586),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1586),
.Y(n_2005)
);

BUFx6f_ASAP7_75t_L g2006 ( 
.A(n_1590),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1568),
.A2(n_1014),
.B1(n_557),
.B2(n_768),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_L g2008 ( 
.A(n_1590),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1595),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1515),
.B(n_1263),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1595),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1603),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1603),
.B(n_1265),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1611),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1611),
.A2(n_776),
.B1(n_921),
.B2(n_566),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1614),
.Y(n_2016)
);

INVx4_ASAP7_75t_L g2017 ( 
.A(n_1614),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1616),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1616),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1637),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1637),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1648),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1648),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1654),
.B(n_1267),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1654),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1659),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1659),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1660),
.B(n_828),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1660),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1670),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1670),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1678),
.B(n_1086),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1678),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_1680),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1680),
.Y(n_2035)
);

INVx3_ASAP7_75t_L g2036 ( 
.A(n_1518),
.Y(n_2036)
);

BUFx6f_ASAP7_75t_L g2037 ( 
.A(n_1518),
.Y(n_2037)
);

INVx6_ASAP7_75t_L g2038 ( 
.A(n_1540),
.Y(n_2038)
);

BUFx2_ASAP7_75t_L g2039 ( 
.A(n_1540),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1442),
.B(n_1089),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1461),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1715),
.B(n_581),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_SL g2043 ( 
.A1(n_1696),
.A2(n_1790),
.B1(n_1800),
.B2(n_1707),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1700),
.A2(n_813),
.B1(n_866),
.B2(n_844),
.Y(n_2044)
);

OA21x2_ASAP7_75t_L g2045 ( 
.A1(n_1688),
.A2(n_1090),
.B(n_1089),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1688),
.Y(n_2046)
);

INVx4_ASAP7_75t_L g2047 ( 
.A(n_1692),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1701),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1780),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1757),
.B(n_976),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1692),
.B(n_1090),
.Y(n_2051)
);

BUFx3_ASAP7_75t_L g2052 ( 
.A(n_1891),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1692),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1780),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1692),
.B(n_1093),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1802),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1689),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1715),
.B(n_586),
.Y(n_2058)
);

BUFx8_ASAP7_75t_L g2059 ( 
.A(n_1785),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_1761),
.A2(n_801),
.B1(n_676),
.B2(n_683),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1802),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1716),
.B(n_623),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1985),
.B(n_1385),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1689),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1691),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1816),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1816),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1716),
.B(n_674),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1860),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1724),
.B(n_748),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1860),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1873),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1691),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1873),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1877),
.Y(n_2075)
);

HB1xp67_ASAP7_75t_L g2076 ( 
.A(n_2013),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1724),
.B(n_748),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1693),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1877),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1882),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1693),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1882),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1748),
.B(n_857),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_2013),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_1986),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1892),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1892),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1892),
.Y(n_2088)
);

NAND2x1p5_ASAP7_75t_L g2089 ( 
.A(n_1945),
.B(n_1043),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1702),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1892),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1702),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1889),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1704),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1748),
.B(n_857),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_2024),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1889),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1747),
.Y(n_2098)
);

HB1xp67_ASAP7_75t_L g2099 ( 
.A(n_2024),
.Y(n_2099)
);

AND2x6_ASAP7_75t_L g2100 ( 
.A(n_1944),
.B(n_1900),
.Y(n_2100)
);

INVx3_ASAP7_75t_L g2101 ( 
.A(n_1695),
.Y(n_2101)
);

INVxp67_ASAP7_75t_L g2102 ( 
.A(n_1757),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1750),
.B(n_859),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1747),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1940),
.B(n_981),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1747),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1747),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1749),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1749),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1695),
.B(n_1093),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1751),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1704),
.Y(n_2112)
);

NAND2xp33_ASAP7_75t_SL g2113 ( 
.A(n_1799),
.B(n_859),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1750),
.B(n_881),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1945),
.B(n_1268),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_1695),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1713),
.Y(n_2117)
);

BUFx2_ASAP7_75t_L g2118 ( 
.A(n_1996),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_1695),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1751),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1758),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1700),
.A2(n_844),
.B1(n_914),
.B2(n_866),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1758),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1713),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1753),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_1706),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_1731),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1753),
.Y(n_2128)
);

INVxp67_ASAP7_75t_L g2129 ( 
.A(n_1940),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1762),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1721),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1762),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1764),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1764),
.Y(n_2134)
);

HB1xp67_ASAP7_75t_L g2135 ( 
.A(n_1994),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1769),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1769),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1771),
.Y(n_2138)
);

INVx1_ASAP7_75t_SL g2139 ( 
.A(n_1696),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1771),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1721),
.Y(n_2141)
);

INVx3_ASAP7_75t_L g2142 ( 
.A(n_1706),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1772),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1772),
.Y(n_2144)
);

OAI22xp33_ASAP7_75t_SL g2145 ( 
.A1(n_2028),
.A2(n_973),
.B1(n_931),
.B2(n_685),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1773),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_SL g2147 ( 
.A(n_1807),
.B(n_1470),
.Y(n_2147)
);

AOI22xp5_ASAP7_75t_L g2148 ( 
.A1(n_1700),
.A2(n_914),
.B1(n_940),
.B2(n_933),
.Y(n_2148)
);

CKINVDCx8_ASAP7_75t_R g2149 ( 
.A(n_1997),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1773),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1917),
.B(n_1471),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_1945),
.B(n_1272),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1820),
.B(n_881),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1779),
.B(n_1944),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1776),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1894),
.B(n_888),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_1690),
.B(n_1472),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1729),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1776),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1777),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1777),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1789),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1789),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1792),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1792),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1965),
.B(n_1472),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_1817),
.A2(n_686),
.B1(n_687),
.B2(n_671),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1805),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1731),
.Y(n_2169)
);

AND2x2_ASAP7_75t_SL g2170 ( 
.A(n_1963),
.B(n_678),
.Y(n_2170)
);

AOI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_1965),
.A2(n_1987),
.B1(n_1817),
.B2(n_1994),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1729),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1805),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1730),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1994),
.B(n_1094),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1809),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1809),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1811),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1730),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1811),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1718),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_1834),
.Y(n_2182)
);

INVx3_ASAP7_75t_L g2183 ( 
.A(n_1706),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1822),
.Y(n_2184)
);

BUFx6f_ASAP7_75t_L g2185 ( 
.A(n_1731),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1822),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1827),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1718),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1718),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1827),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1840),
.Y(n_2191)
);

AND2x4_ASAP7_75t_L g2192 ( 
.A(n_1945),
.B(n_1273),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1731),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1840),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1843),
.Y(n_2195)
);

NOR2x1_ASAP7_75t_L g2196 ( 
.A(n_1911),
.B(n_1276),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1843),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1733),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1733),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1894),
.B(n_888),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1991),
.B(n_545),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1844),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1844),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1845),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_1739),
.Y(n_2205)
);

INVxp67_ASAP7_75t_L g2206 ( 
.A(n_1989),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1838),
.B(n_562),
.Y(n_2207)
);

NOR2x1_ASAP7_75t_L g2208 ( 
.A(n_1911),
.B(n_1284),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1845),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1838),
.B(n_651),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_1987),
.A2(n_933),
.B1(n_962),
.B2(n_940),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1848),
.Y(n_2212)
);

INVx3_ASAP7_75t_L g2213 ( 
.A(n_1698),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1838),
.B(n_651),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_1739),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1863),
.B(n_868),
.Y(n_2216)
);

BUFx6f_ASAP7_75t_SL g2217 ( 
.A(n_2003),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1848),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1929),
.B(n_1094),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1862),
.Y(n_2220)
);

BUFx6f_ASAP7_75t_L g2221 ( 
.A(n_1739),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_1929),
.B(n_962),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1733),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1698),
.Y(n_2224)
);

BUFx6f_ASAP7_75t_L g2225 ( 
.A(n_1739),
.Y(n_2225)
);

NAND2xp33_ASAP7_75t_SL g2226 ( 
.A(n_1850),
.B(n_868),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_1929),
.B(n_965),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1863),
.B(n_965),
.Y(n_2228)
);

INVx3_ASAP7_75t_L g2229 ( 
.A(n_1698),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1862),
.Y(n_2230)
);

BUFx10_ASAP7_75t_L g2231 ( 
.A(n_1957),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1743),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1880),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1863),
.B(n_969),
.Y(n_2234)
);

AOI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_1989),
.A2(n_969),
.B1(n_725),
.B2(n_603),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1880),
.Y(n_2236)
);

INVx8_ASAP7_75t_L g2237 ( 
.A(n_1945),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1743),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1888),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1888),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_1740),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_1967),
.B(n_678),
.Y(n_2242)
);

NAND2xp33_ASAP7_75t_SL g2243 ( 
.A(n_1920),
.B(n_853),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1743),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_1891),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1694),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1703),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1705),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_1740),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1711),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1886),
.B(n_853),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1886),
.Y(n_2252)
);

OAI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_1842),
.A2(n_689),
.B1(n_694),
.B2(n_692),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1712),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_1754),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1714),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1886),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1719),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_1890),
.B(n_696),
.Y(n_2259)
);

NOR3xp33_ASAP7_75t_L g2260 ( 
.A(n_2032),
.B(n_699),
.C(n_697),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1687),
.B(n_854),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1745),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_1710),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1720),
.Y(n_2264)
);

INVx3_ASAP7_75t_L g2265 ( 
.A(n_1754),
.Y(n_2265)
);

BUFx2_ASAP7_75t_L g2266 ( 
.A(n_1707),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1745),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_1745),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_1710),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_1740),
.Y(n_2270)
);

INVx3_ASAP7_75t_L g2271 ( 
.A(n_1754),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_1935),
.B(n_1901),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_1967),
.B(n_678),
.Y(n_2273)
);

OR2x2_ASAP7_75t_L g2274 ( 
.A(n_1836),
.B(n_1387),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1722),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_SL g2276 ( 
.A(n_2003),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1756),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1723),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_1967),
.B(n_786),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1726),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1736),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_1756),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_1883),
.B(n_701),
.Y(n_2283)
);

INVx3_ASAP7_75t_L g2284 ( 
.A(n_1754),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1738),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_1876),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1746),
.Y(n_2287)
);

AND2x6_ASAP7_75t_L g2288 ( 
.A(n_1993),
.B(n_786),
.Y(n_2288)
);

OAI22xp5_ASAP7_75t_SL g2289 ( 
.A1(n_1790),
.A2(n_1393),
.B1(n_1395),
.B2(n_1387),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_1993),
.B(n_1475),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_1759),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1752),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1770),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1727),
.B(n_1734),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1782),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1756),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1783),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_1740),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1787),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_1710),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1791),
.Y(n_2301)
);

AOI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_1915),
.A2(n_725),
.B1(n_606),
.B2(n_610),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_1710),
.Y(n_2303)
);

OR2x2_ASAP7_75t_L g2304 ( 
.A(n_1851),
.B(n_1393),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1793),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_1767),
.B(n_1475),
.Y(n_2306)
);

AOI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_1915),
.A2(n_611),
.B1(n_614),
.B2(n_598),
.Y(n_2307)
);

BUFx6f_ASAP7_75t_SL g2308 ( 
.A(n_2034),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1796),
.Y(n_2309)
);

BUFx2_ASAP7_75t_L g2310 ( 
.A(n_1800),
.Y(n_2310)
);

AND2x6_ASAP7_75t_L g2311 ( 
.A(n_1977),
.B(n_786),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_1767),
.B(n_1483),
.Y(n_2312)
);

BUFx3_ASAP7_75t_L g2313 ( 
.A(n_1891),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1797),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1801),
.Y(n_2315)
);

INVx8_ASAP7_75t_L g2316 ( 
.A(n_1915),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1774),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_1977),
.B(n_823),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_1759),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1803),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_1759),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1808),
.Y(n_2322)
);

BUFx2_ASAP7_75t_L g2323 ( 
.A(n_1804),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1812),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1727),
.B(n_854),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1818),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1819),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_1774),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1821),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1824),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_1829),
.Y(n_2331)
);

INVx4_ASAP7_75t_L g2332 ( 
.A(n_1829),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1828),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1774),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_SL g2335 ( 
.A(n_1866),
.B(n_1483),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1841),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1727),
.B(n_858),
.Y(n_2337)
);

AOI22xp5_ASAP7_75t_L g2338 ( 
.A1(n_1915),
.A2(n_624),
.B1(n_628),
.B2(n_616),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1849),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_1977),
.B(n_823),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_1855),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1861),
.Y(n_2342)
);

NAND2xp33_ASAP7_75t_SL g2343 ( 
.A(n_1920),
.B(n_858),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1867),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_1868),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_1935),
.B(n_1285),
.Y(n_2346)
);

NAND2xp33_ASAP7_75t_SL g2347 ( 
.A(n_1920),
.B(n_863),
.Y(n_2347)
);

HB1xp67_ASAP7_75t_L g2348 ( 
.A(n_1798),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1814),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1734),
.B(n_863),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_1915),
.A2(n_1763),
.B1(n_1781),
.B2(n_1755),
.Y(n_2351)
);

AND2x6_ASAP7_75t_L g2352 ( 
.A(n_1734),
.B(n_1741),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1814),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1814),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1869),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1870),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_1815),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1871),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_1741),
.B(n_867),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1741),
.B(n_867),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1815),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1815),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_1826),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1874),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_1755),
.B(n_870),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_1878),
.B(n_1485),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1826),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1875),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_1839),
.B(n_703),
.Y(n_2369)
);

INVxp67_ASAP7_75t_L g2370 ( 
.A(n_1907),
.Y(n_2370)
);

HB1xp67_ASAP7_75t_L g2371 ( 
.A(n_1830),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_1826),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_1992),
.B(n_1485),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1887),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1829),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_1759),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_1829),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_1833),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1833),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1833),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_1833),
.Y(n_2381)
);

BUFx6f_ASAP7_75t_L g2382 ( 
.A(n_1854),
.Y(n_2382)
);

OAI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_1839),
.A2(n_711),
.B1(n_714),
.B2(n_708),
.Y(n_2383)
);

INVxp67_ASAP7_75t_L g2384 ( 
.A(n_1907),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1854),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1854),
.Y(n_2386)
);

BUFx6f_ASAP7_75t_L g2387 ( 
.A(n_1854),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1858),
.Y(n_2388)
);

INVx3_ASAP7_75t_L g2389 ( 
.A(n_1766),
.Y(n_2389)
);

OAI22xp5_ASAP7_75t_SL g2390 ( 
.A1(n_1804),
.A2(n_1403),
.B1(n_1407),
.B2(n_1395),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_1766),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_1958),
.Y(n_2392)
);

BUFx6f_ASAP7_75t_L g2393 ( 
.A(n_1858),
.Y(n_2393)
);

BUFx6f_ASAP7_75t_L g2394 ( 
.A(n_1858),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_1920),
.B(n_823),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_1858),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1881),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1881),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_1881),
.Y(n_2399)
);

AND2x6_ASAP7_75t_L g2400 ( 
.A(n_2351),
.B(n_1956),
.Y(n_2400)
);

BUFx2_ASAP7_75t_L g2401 ( 
.A(n_2085),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2294),
.Y(n_2402)
);

INVx2_ASAP7_75t_SL g2403 ( 
.A(n_2118),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2046),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2093),
.Y(n_2405)
);

BUFx3_ASAP7_75t_L g2406 ( 
.A(n_2059),
.Y(n_2406)
);

INVx3_ASAP7_75t_L g2407 ( 
.A(n_2237),
.Y(n_2407)
);

OR2x2_ASAP7_75t_L g2408 ( 
.A(n_2274),
.B(n_2041),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_2237),
.Y(n_2409)
);

INVx1_ASAP7_75t_SL g2410 ( 
.A(n_2139),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_2237),
.Y(n_2411)
);

INVx5_ASAP7_75t_L g2412 ( 
.A(n_2316),
.Y(n_2412)
);

BUFx3_ASAP7_75t_L g2413 ( 
.A(n_2059),
.Y(n_2413)
);

BUFx8_ASAP7_75t_SL g2414 ( 
.A(n_2217),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_2135),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2097),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2050),
.B(n_1958),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2076),
.B(n_1959),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_2149),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2076),
.B(n_1959),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2154),
.B(n_1837),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2102),
.B(n_2001),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2046),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_SL g2424 ( 
.A(n_2272),
.B(n_1956),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2057),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_2053),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2108),
.Y(n_2427)
);

BUFx3_ASAP7_75t_L g2428 ( 
.A(n_2059),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2102),
.B(n_2001),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2109),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2111),
.Y(n_2431)
);

AOI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2352),
.A2(n_1937),
.B1(n_1949),
.B2(n_1936),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2120),
.Y(n_2433)
);

BUFx10_ASAP7_75t_L g2434 ( 
.A(n_2217),
.Y(n_2434)
);

BUFx10_ASAP7_75t_L g2435 ( 
.A(n_2276),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2287),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2057),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2292),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_2272),
.B(n_1956),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2293),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2295),
.Y(n_2441)
);

INVxp67_ASAP7_75t_SL g2442 ( 
.A(n_2331),
.Y(n_2442)
);

INVx1_ASAP7_75t_SL g2443 ( 
.A(n_2157),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2149),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_2206),
.B(n_2040),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_R g2446 ( 
.A(n_2113),
.B(n_1981),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2332),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2297),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2206),
.B(n_1998),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2352),
.B(n_2001),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_2231),
.B(n_1998),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2231),
.B(n_1901),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_2289),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_2053),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2299),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2064),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2084),
.B(n_1936),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2301),
.Y(n_2458)
);

INVx4_ASAP7_75t_L g2459 ( 
.A(n_2052),
.Y(n_2459)
);

BUFx6f_ASAP7_75t_L g2460 ( 
.A(n_2053),
.Y(n_2460)
);

OAI21xp33_ASAP7_75t_SL g2461 ( 
.A1(n_2171),
.A2(n_1708),
.B(n_1697),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2305),
.Y(n_2462)
);

NAND3xp33_ASAP7_75t_L g2463 ( 
.A(n_2369),
.B(n_1981),
.C(n_1949),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2352),
.B(n_1755),
.Y(n_2464)
);

AND2x6_ASAP7_75t_L g2465 ( 
.A(n_2115),
.B(n_2152),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2309),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2352),
.B(n_1763),
.Y(n_2467)
);

OAI21xp33_ASAP7_75t_L g2468 ( 
.A1(n_2259),
.A2(n_1709),
.B(n_1937),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_SL g2469 ( 
.A(n_2272),
.B(n_1956),
.Y(n_2469)
);

INVx5_ASAP7_75t_L g2470 ( 
.A(n_2316),
.Y(n_2470)
);

BUFx6f_ASAP7_75t_L g2471 ( 
.A(n_2053),
.Y(n_2471)
);

BUFx3_ASAP7_75t_L g2472 ( 
.A(n_2052),
.Y(n_2472)
);

HB1xp67_ASAP7_75t_L g2473 ( 
.A(n_2135),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_2231),
.B(n_1901),
.Y(n_2474)
);

AND2x6_ASAP7_75t_L g2475 ( 
.A(n_2115),
.B(n_1971),
.Y(n_2475)
);

BUFx3_ASAP7_75t_L g2476 ( 
.A(n_2245),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_L g2477 ( 
.A(n_2129),
.B(n_1904),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2314),
.Y(n_2478)
);

HB1xp67_ASAP7_75t_L g2479 ( 
.A(n_2048),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2315),
.Y(n_2480)
);

OR2x2_ASAP7_75t_L g2481 ( 
.A(n_2063),
.B(n_2041),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2352),
.B(n_1763),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2320),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2322),
.Y(n_2484)
);

OR2x2_ASAP7_75t_L g2485 ( 
.A(n_2306),
.B(n_2312),
.Y(n_2485)
);

NAND2xp33_ASAP7_75t_L g2486 ( 
.A(n_2252),
.B(n_1971),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2241),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2324),
.Y(n_2488)
);

AOI22xp33_ASAP7_75t_L g2489 ( 
.A1(n_2170),
.A2(n_1915),
.B1(n_1963),
.B2(n_2028),
.Y(n_2489)
);

BUFx3_ASAP7_75t_L g2490 ( 
.A(n_2245),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2313),
.B(n_1971),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2084),
.B(n_2096),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2252),
.B(n_1781),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2326),
.Y(n_2494)
);

INVxp67_ASAP7_75t_SL g2495 ( 
.A(n_2331),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2313),
.B(n_1971),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2064),
.Y(n_2497)
);

OR2x2_ASAP7_75t_L g2498 ( 
.A(n_2048),
.B(n_1785),
.Y(n_2498)
);

AND2x6_ASAP7_75t_L g2499 ( 
.A(n_2115),
.B(n_1973),
.Y(n_2499)
);

INVx2_ASAP7_75t_SL g2500 ( 
.A(n_2346),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2152),
.B(n_1973),
.Y(n_2501)
);

INVx2_ASAP7_75t_SL g2502 ( 
.A(n_2346),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2327),
.Y(n_2503)
);

AND2x4_ASAP7_75t_L g2504 ( 
.A(n_2152),
.B(n_1973),
.Y(n_2504)
);

BUFx6f_ASAP7_75t_L g2505 ( 
.A(n_2241),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2390),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2065),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2065),
.Y(n_2508)
);

INVx2_ASAP7_75t_SL g2509 ( 
.A(n_2346),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2329),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2257),
.B(n_1781),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_SL g2512 ( 
.A(n_2192),
.B(n_1973),
.Y(n_2512)
);

INVx3_ASAP7_75t_L g2513 ( 
.A(n_2332),
.Y(n_2513)
);

BUFx2_ASAP7_75t_L g2514 ( 
.A(n_2151),
.Y(n_2514)
);

INVx8_ASAP7_75t_L g2515 ( 
.A(n_2316),
.Y(n_2515)
);

BUFx6f_ASAP7_75t_L g2516 ( 
.A(n_2241),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2096),
.B(n_1955),
.Y(n_2517)
);

BUFx6f_ASAP7_75t_L g2518 ( 
.A(n_2241),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2330),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2129),
.B(n_1904),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2073),
.Y(n_2521)
);

INVx3_ASAP7_75t_L g2522 ( 
.A(n_2332),
.Y(n_2522)
);

AO22x2_ASAP7_75t_L g2523 ( 
.A1(n_2166),
.A2(n_2011),
.B1(n_2019),
.B2(n_2005),
.Y(n_2523)
);

AOI22xp33_ASAP7_75t_L g2524 ( 
.A1(n_2170),
.A2(n_1881),
.B1(n_1813),
.B2(n_1775),
.Y(n_2524)
);

AND2x4_ASAP7_75t_L g2525 ( 
.A(n_2192),
.B(n_1976),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2266),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2073),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2333),
.Y(n_2528)
);

OR2x2_ASAP7_75t_L g2529 ( 
.A(n_2304),
.B(n_1864),
.Y(n_2529)
);

BUFx2_ASAP7_75t_L g2530 ( 
.A(n_2310),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2336),
.Y(n_2531)
);

BUFx3_ASAP7_75t_L g2532 ( 
.A(n_2323),
.Y(n_2532)
);

OR2x2_ASAP7_75t_L g2533 ( 
.A(n_2099),
.B(n_1864),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_L g2534 ( 
.A(n_2370),
.B(n_1904),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_SL g2535 ( 
.A(n_2192),
.B(n_1976),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_2276),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_L g2537 ( 
.A(n_2370),
.B(n_1943),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2078),
.Y(n_2538)
);

INVx4_ASAP7_75t_L g2539 ( 
.A(n_2331),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_2366),
.Y(n_2540)
);

NOR2xp33_ASAP7_75t_L g2541 ( 
.A(n_2384),
.B(n_1943),
.Y(n_2541)
);

INVx3_ASAP7_75t_L g2542 ( 
.A(n_2047),
.Y(n_2542)
);

INVxp33_ASAP7_75t_L g2543 ( 
.A(n_2290),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2339),
.Y(n_2544)
);

INVx3_ASAP7_75t_L g2545 ( 
.A(n_2047),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2078),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2257),
.B(n_1788),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2262),
.B(n_2267),
.Y(n_2548)
);

OAI22xp33_ASAP7_75t_L g2549 ( 
.A1(n_2122),
.A2(n_1846),
.B1(n_1964),
.B2(n_1955),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2099),
.B(n_1964),
.Y(n_2550)
);

HB1xp67_ASAP7_75t_L g2551 ( 
.A(n_2348),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2081),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2341),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2081),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2105),
.B(n_1912),
.Y(n_2555)
);

OR2x6_ASAP7_75t_L g2556 ( 
.A(n_2043),
.B(n_1891),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_SL g2557 ( 
.A(n_2331),
.B(n_1976),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2373),
.B(n_1912),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2342),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2344),
.Y(n_2560)
);

BUFx6f_ASAP7_75t_L g2561 ( 
.A(n_2249),
.Y(n_2561)
);

INVx8_ASAP7_75t_L g2562 ( 
.A(n_2308),
.Y(n_2562)
);

BUFx3_ASAP7_75t_L g2563 ( 
.A(n_2348),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2345),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2355),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2090),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2090),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2356),
.Y(n_2568)
);

INVxp67_ASAP7_75t_L g2569 ( 
.A(n_2182),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2262),
.B(n_1788),
.Y(n_2570)
);

BUFx6f_ASAP7_75t_L g2571 ( 
.A(n_2249),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2308),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2092),
.Y(n_2573)
);

BUFx3_ASAP7_75t_L g2574 ( 
.A(n_2371),
.Y(n_2574)
);

AOI22xp33_ASAP7_75t_L g2575 ( 
.A1(n_2121),
.A2(n_1813),
.B1(n_1775),
.B2(n_1786),
.Y(n_2575)
);

AOI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2259),
.A2(n_1742),
.B1(n_1831),
.B2(n_1938),
.Y(n_2576)
);

INVx4_ASAP7_75t_L g2577 ( 
.A(n_2382),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2358),
.Y(n_2578)
);

NOR2xp33_ASAP7_75t_L g2579 ( 
.A(n_2384),
.B(n_2392),
.Y(n_2579)
);

NOR2x1p5_ASAP7_75t_L g2580 ( 
.A(n_2123),
.B(n_1744),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2267),
.B(n_1788),
.Y(n_2581)
);

BUFx2_ASAP7_75t_L g2582 ( 
.A(n_2371),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2364),
.Y(n_2583)
);

INVx4_ASAP7_75t_L g2584 ( 
.A(n_2382),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_SL g2585 ( 
.A(n_2382),
.B(n_1976),
.Y(n_2585)
);

INVx3_ASAP7_75t_L g2586 ( 
.A(n_2047),
.Y(n_2586)
);

BUFx10_ASAP7_75t_L g2587 ( 
.A(n_2369),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_SL g2588 ( 
.A(n_2382),
.B(n_1943),
.Y(n_2588)
);

AND2x6_ASAP7_75t_L g2589 ( 
.A(n_2387),
.B(n_1946),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2268),
.B(n_1832),
.Y(n_2590)
);

INVx3_ASAP7_75t_L g2591 ( 
.A(n_2249),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2268),
.B(n_1813),
.Y(n_2592)
);

INVx5_ASAP7_75t_L g2593 ( 
.A(n_2387),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2182),
.B(n_1908),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2286),
.B(n_1908),
.Y(n_2595)
);

INVx3_ASAP7_75t_L g2596 ( 
.A(n_2249),
.Y(n_2596)
);

OR2x2_ASAP7_75t_SL g2597 ( 
.A(n_2392),
.B(n_2006),
.Y(n_2597)
);

INVx3_ASAP7_75t_L g2598 ( 
.A(n_2270),
.Y(n_2598)
);

BUFx3_ASAP7_75t_L g2599 ( 
.A(n_2286),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2270),
.Y(n_2600)
);

CKINVDCx11_ASAP7_75t_R g2601 ( 
.A(n_2147),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2277),
.B(n_1813),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2368),
.Y(n_2603)
);

OR2x2_ASAP7_75t_L g2604 ( 
.A(n_2042),
.B(n_1865),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2335),
.B(n_1910),
.Y(n_2605)
);

BUFx6f_ASAP7_75t_L g2606 ( 
.A(n_2270),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2374),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2277),
.B(n_1813),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2270),
.Y(n_2609)
);

AND2x2_ASAP7_75t_SL g2610 ( 
.A(n_2148),
.B(n_2017),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2092),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2282),
.B(n_1813),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_2113),
.Y(n_2613)
);

INVx4_ASAP7_75t_SL g2614 ( 
.A(n_2311),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2094),
.Y(n_2615)
);

BUFx6f_ASAP7_75t_L g2616 ( 
.A(n_2298),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2175),
.B(n_1946),
.Y(n_2617)
);

AND2x4_ASAP7_75t_L g2618 ( 
.A(n_2219),
.B(n_1946),
.Y(n_2618)
);

AND2x6_ASAP7_75t_L g2619 ( 
.A(n_2387),
.B(n_1982),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2282),
.B(n_2296),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2296),
.B(n_1982),
.Y(n_2621)
);

AND2x6_ASAP7_75t_L g2622 ( 
.A(n_2387),
.B(n_1982),
.Y(n_2622)
);

INVx4_ASAP7_75t_L g2623 ( 
.A(n_2393),
.Y(n_2623)
);

NAND3xp33_ASAP7_75t_SL g2624 ( 
.A(n_2235),
.B(n_1910),
.C(n_1941),
.Y(n_2624)
);

INVx4_ASAP7_75t_L g2625 ( 
.A(n_2393),
.Y(n_2625)
);

BUFx3_ASAP7_75t_L g2626 ( 
.A(n_2049),
.Y(n_2626)
);

AND2x6_ASAP7_75t_L g2627 ( 
.A(n_2393),
.B(n_1990),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2094),
.Y(n_2628)
);

BUFx10_ASAP7_75t_L g2629 ( 
.A(n_2283),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2112),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_L g2631 ( 
.A(n_2175),
.B(n_1990),
.Y(n_2631)
);

AOI22xp33_ASAP7_75t_L g2632 ( 
.A1(n_2288),
.A2(n_1775),
.B1(n_1786),
.B2(n_1766),
.Y(n_2632)
);

NOR2xp33_ASAP7_75t_L g2633 ( 
.A(n_2219),
.B(n_1990),
.Y(n_2633)
);

INVx4_ASAP7_75t_SL g2634 ( 
.A(n_2311),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2112),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2317),
.B(n_1766),
.Y(n_2636)
);

INVx5_ASAP7_75t_L g2637 ( 
.A(n_2393),
.Y(n_2637)
);

OR2x6_ASAP7_75t_L g2638 ( 
.A(n_2089),
.B(n_2038),
.Y(n_2638)
);

INVx4_ASAP7_75t_L g2639 ( 
.A(n_2394),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2058),
.B(n_1954),
.Y(n_2640)
);

AND2x4_ASAP7_75t_L g2641 ( 
.A(n_2222),
.B(n_1778),
.Y(n_2641)
);

INVx4_ASAP7_75t_SL g2642 ( 
.A(n_2311),
.Y(n_2642)
);

BUFx3_ASAP7_75t_L g2643 ( 
.A(n_2054),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2317),
.B(n_1775),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2328),
.B(n_1786),
.Y(n_2645)
);

INVxp67_ASAP7_75t_L g2646 ( 
.A(n_2222),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2298),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_SL g2648 ( 
.A(n_2394),
.B(n_1921),
.Y(n_2648)
);

HB1xp67_ASAP7_75t_L g2649 ( 
.A(n_2232),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2246),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2062),
.B(n_2010),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2247),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2248),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_SL g2654 ( 
.A(n_2394),
.B(n_1921),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2250),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_L g2656 ( 
.A(n_2068),
.B(n_1968),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2227),
.B(n_1778),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2328),
.B(n_1825),
.Y(n_2658)
);

AOI22xp33_ASAP7_75t_L g2659 ( 
.A1(n_2288),
.A2(n_1825),
.B1(n_1786),
.B2(n_1847),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2254),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_R g2661 ( 
.A(n_2226),
.B(n_1744),
.Y(n_2661)
);

AND2x4_ASAP7_75t_L g2662 ( 
.A(n_2227),
.B(n_2056),
.Y(n_2662)
);

INVx4_ASAP7_75t_L g2663 ( 
.A(n_2394),
.Y(n_2663)
);

BUFx6f_ASAP7_75t_L g2664 ( 
.A(n_2298),
.Y(n_2664)
);

NOR2xp33_ASAP7_75t_L g2665 ( 
.A(n_2283),
.B(n_1925),
.Y(n_2665)
);

BUFx2_ASAP7_75t_L g2666 ( 
.A(n_2311),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_2242),
.B(n_1953),
.Y(n_2667)
);

INVx3_ASAP7_75t_L g2668 ( 
.A(n_2298),
.Y(n_2668)
);

INVx4_ASAP7_75t_L g2669 ( 
.A(n_2399),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2256),
.Y(n_2670)
);

INVx2_ASAP7_75t_SL g2671 ( 
.A(n_2196),
.Y(n_2671)
);

INVx3_ASAP7_75t_L g2672 ( 
.A(n_2127),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_2226),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2325),
.B(n_1784),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2258),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_2061),
.Y(n_2676)
);

AOI22xp5_ASAP7_75t_L g2677 ( 
.A1(n_2288),
.A2(n_1931),
.B1(n_1984),
.B2(n_1950),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2264),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2275),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2278),
.Y(n_2680)
);

INVx6_ASAP7_75t_L g2681 ( 
.A(n_2127),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2334),
.B(n_1825),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2399),
.B(n_1924),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2117),
.Y(n_2684)
);

INVxp67_ASAP7_75t_L g2685 ( 
.A(n_2311),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2280),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2337),
.B(n_1784),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2334),
.B(n_1825),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2349),
.B(n_1835),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2281),
.Y(n_2690)
);

INVx4_ASAP7_75t_SL g2691 ( 
.A(n_2288),
.Y(n_2691)
);

INVx4_ASAP7_75t_L g2692 ( 
.A(n_2399),
.Y(n_2692)
);

INVx1_ASAP7_75t_SL g2693 ( 
.A(n_2243),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2117),
.Y(n_2694)
);

INVx1_ASAP7_75t_SL g2695 ( 
.A(n_2243),
.Y(n_2695)
);

NOR2xp33_ASAP7_75t_L g2696 ( 
.A(n_2242),
.B(n_1913),
.Y(n_2696)
);

HB1xp67_ASAP7_75t_L g2697 ( 
.A(n_2232),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2285),
.Y(n_2698)
);

BUFx6f_ASAP7_75t_L g2699 ( 
.A(n_2399),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2125),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2350),
.B(n_1794),
.Y(n_2701)
);

NOR2xp33_ASAP7_75t_SL g2702 ( 
.A(n_2288),
.B(n_1794),
.Y(n_2702)
);

OAI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2349),
.A2(n_1931),
.B1(n_1932),
.B2(n_1924),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2353),
.B(n_1932),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2124),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2128),
.Y(n_2706)
);

INVx2_ASAP7_75t_SL g2707 ( 
.A(n_2208),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_L g2708 ( 
.A(n_2273),
.B(n_1913),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_2066),
.Y(n_2709)
);

INVx4_ASAP7_75t_L g2710 ( 
.A(n_2263),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2124),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_SL g2712 ( 
.A(n_2260),
.B(n_1942),
.Y(n_2712)
);

NAND3xp33_ASAP7_75t_L g2713 ( 
.A(n_2260),
.B(n_1853),
.C(n_1795),
.Y(n_2713)
);

NAND3xp33_ASAP7_75t_L g2714 ( 
.A(n_2060),
.B(n_1853),
.C(n_1795),
.Y(n_2714)
);

BUFx6f_ASAP7_75t_SL g2715 ( 
.A(n_2100),
.Y(n_2715)
);

INVx4_ASAP7_75t_L g2716 ( 
.A(n_2263),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2130),
.Y(n_2717)
);

INVx3_ASAP7_75t_L g2718 ( 
.A(n_2127),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2353),
.B(n_1942),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2132),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2131),
.Y(n_2721)
);

NOR2x1p5_ASAP7_75t_L g2722 ( 
.A(n_2359),
.B(n_1760),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_SL g2723 ( 
.A(n_2044),
.B(n_1950),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2133),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2354),
.B(n_1952),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_L g2726 ( 
.A(n_2127),
.Y(n_2726)
);

AND2x4_ASAP7_75t_L g2727 ( 
.A(n_2067),
.B(n_1952),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2354),
.B(n_1969),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2253),
.Y(n_2729)
);

CKINVDCx5p33_ASAP7_75t_R g2730 ( 
.A(n_2343),
.Y(n_2730)
);

NOR2xp33_ASAP7_75t_L g2731 ( 
.A(n_2273),
.B(n_1969),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2134),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2357),
.B(n_1983),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2136),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2131),
.Y(n_2735)
);

INVx3_ASAP7_75t_L g2736 ( 
.A(n_2169),
.Y(n_2736)
);

AND2x4_ASAP7_75t_L g2737 ( 
.A(n_2069),
.B(n_2071),
.Y(n_2737)
);

INVx1_ASAP7_75t_SL g2738 ( 
.A(n_2343),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2072),
.B(n_1983),
.Y(n_2739)
);

NOR2xp33_ASAP7_75t_L g2740 ( 
.A(n_2279),
.B(n_1984),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2141),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2137),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2141),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2357),
.B(n_1717),
.Y(n_2744)
);

INVx2_ASAP7_75t_SL g2745 ( 
.A(n_2360),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2158),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2255),
.B(n_1916),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2361),
.B(n_1732),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2138),
.Y(n_2749)
);

AND2x4_ASAP7_75t_L g2750 ( 
.A(n_2074),
.B(n_1897),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2361),
.B(n_1737),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2140),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2158),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2172),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2362),
.B(n_1847),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_SL g2756 ( 
.A(n_2255),
.B(n_1918),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2143),
.Y(n_2757)
);

AOI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2468),
.A2(n_1879),
.B1(n_1893),
.B2(n_1859),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2665),
.B(n_2075),
.Y(n_2759)
);

OAI22xp5_ASAP7_75t_L g2760 ( 
.A1(n_2576),
.A2(n_2080),
.B1(n_2082),
.B2(n_2079),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_L g2761 ( 
.A(n_2665),
.B(n_1859),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2421),
.B(n_2362),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2436),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_2656),
.B(n_1879),
.Y(n_2764)
);

OAI221xp5_ASAP7_75t_L g2765 ( 
.A1(n_2432),
.A2(n_1872),
.B1(n_2007),
.B2(n_2015),
.C(n_2011),
.Y(n_2765)
);

INVxp67_ASAP7_75t_L g2766 ( 
.A(n_2401),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2421),
.B(n_2363),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_L g2768 ( 
.A(n_2656),
.B(n_1893),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_SL g2769 ( 
.A(n_2702),
.B(n_2006),
.Y(n_2769)
);

INVx3_ASAP7_75t_L g2770 ( 
.A(n_2515),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2640),
.B(n_2363),
.Y(n_2771)
);

OAI22xp33_ASAP7_75t_L g2772 ( 
.A1(n_2729),
.A2(n_2017),
.B1(n_2006),
.B2(n_2012),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2404),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2640),
.B(n_2367),
.Y(n_2774)
);

OR2x2_ASAP7_75t_L g2775 ( 
.A(n_2485),
.B(n_2009),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2423),
.Y(n_2776)
);

OAI22xp5_ASAP7_75t_L g2777 ( 
.A1(n_2489),
.A2(n_2251),
.B1(n_2211),
.B2(n_2367),
.Y(n_2777)
);

AND2x2_ASAP7_75t_L g2778 ( 
.A(n_2651),
.B(n_1975),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2549),
.B(n_2009),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_SL g2780 ( 
.A(n_2549),
.B(n_2006),
.Y(n_2780)
);

OR2x6_ASAP7_75t_L g2781 ( 
.A(n_2562),
.B(n_2038),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2445),
.B(n_2372),
.Y(n_2782)
);

AND2x6_ASAP7_75t_SL g2783 ( 
.A(n_2605),
.B(n_1999),
.Y(n_2783)
);

NOR2xp33_ASAP7_75t_L g2784 ( 
.A(n_2463),
.B(n_2016),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2425),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2437),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2438),
.Y(n_2787)
);

NOR2xp33_ASAP7_75t_L g2788 ( 
.A(n_2594),
.B(n_2016),
.Y(n_2788)
);

BUFx6f_ASAP7_75t_L g2789 ( 
.A(n_2409),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2446),
.B(n_2008),
.Y(n_2790)
);

INVx1_ASAP7_75t_SL g2791 ( 
.A(n_2582),
.Y(n_2791)
);

INVx2_ASAP7_75t_SL g2792 ( 
.A(n_2562),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2445),
.B(n_2365),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_SL g2794 ( 
.A(n_2446),
.B(n_2008),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2449),
.B(n_2100),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2456),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2440),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_SL g2798 ( 
.A(n_2595),
.B(n_2008),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2441),
.Y(n_2799)
);

INVx2_ASAP7_75t_SL g2800 ( 
.A(n_2562),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2558),
.B(n_2005),
.Y(n_2801)
);

OR2x6_ASAP7_75t_L g2802 ( 
.A(n_2515),
.B(n_2038),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2449),
.B(n_2100),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2448),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2402),
.B(n_2100),
.Y(n_2805)
);

INVx3_ASAP7_75t_L g2806 ( 
.A(n_2515),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2455),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2579),
.B(n_2100),
.Y(n_2808)
);

AOI22xp5_ASAP7_75t_L g2809 ( 
.A1(n_2674),
.A2(n_1979),
.B1(n_1961),
.B2(n_2019),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2458),
.Y(n_2810)
);

OAI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2489),
.A2(n_2372),
.B1(n_2238),
.B2(n_2234),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2462),
.Y(n_2812)
);

NAND2xp33_ASAP7_75t_L g2813 ( 
.A(n_2589),
.B(n_1760),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2466),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2478),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2579),
.B(n_1898),
.Y(n_2816)
);

NOR2xp33_ASAP7_75t_SL g2817 ( 
.A(n_2419),
.B(n_2017),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_SL g2818 ( 
.A(n_2629),
.B(n_2008),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_SL g2819 ( 
.A(n_2629),
.B(n_2012),
.Y(n_2819)
);

INVx3_ASAP7_75t_L g2820 ( 
.A(n_2409),
.Y(n_2820)
);

A2O1A1Ixp33_ASAP7_75t_L g2821 ( 
.A1(n_2667),
.A2(n_2347),
.B(n_2279),
.C(n_2340),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2534),
.B(n_2070),
.Y(n_2822)
);

NAND3xp33_ASAP7_75t_L g2823 ( 
.A(n_2451),
.B(n_1923),
.C(n_1995),
.Y(n_2823)
);

NAND2x1_ASAP7_75t_L g2824 ( 
.A(n_2681),
.B(n_2255),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2497),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2534),
.B(n_2077),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2537),
.B(n_2541),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2537),
.B(n_2083),
.Y(n_2828)
);

NOR2xp33_ASAP7_75t_L g2829 ( 
.A(n_2543),
.B(n_2025),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_SL g2830 ( 
.A(n_2687),
.B(n_2701),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2667),
.B(n_2238),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2403),
.B(n_2012),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2480),
.Y(n_2833)
);

OR2x6_ASAP7_75t_L g2834 ( 
.A(n_2406),
.B(n_2038),
.Y(n_2834)
);

INVxp67_ASAP7_75t_SL g2835 ( 
.A(n_2551),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2541),
.B(n_2744),
.Y(n_2836)
);

INVxp67_ASAP7_75t_L g2837 ( 
.A(n_2551),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_L g2838 ( 
.A(n_2624),
.B(n_2025),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_SL g2839 ( 
.A(n_2451),
.B(n_2012),
.Y(n_2839)
);

INVx2_ASAP7_75t_SL g2840 ( 
.A(n_2434),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2507),
.Y(n_2841)
);

NAND2x1p5_ASAP7_75t_L g2842 ( 
.A(n_2412),
.B(n_2470),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_SL g2843 ( 
.A(n_2457),
.B(n_2023),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_SL g2844 ( 
.A(n_2517),
.B(n_2023),
.Y(n_2844)
);

NAND2xp33_ASAP7_75t_L g2845 ( 
.A(n_2589),
.B(n_1725),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2744),
.B(n_2144),
.Y(n_2846)
);

NOR2xp33_ASAP7_75t_L g2847 ( 
.A(n_2624),
.B(n_2029),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2508),
.Y(n_2848)
);

AOI22xp33_ASAP7_75t_L g2849 ( 
.A1(n_2417),
.A2(n_2022),
.B1(n_2027),
.B2(n_2021),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2748),
.B(n_2146),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2483),
.Y(n_2851)
);

CKINVDCx5p33_ASAP7_75t_R g2852 ( 
.A(n_2414),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2484),
.Y(n_2853)
);

AOI22xp33_ASAP7_75t_L g2854 ( 
.A1(n_2555),
.A2(n_2022),
.B1(n_2027),
.B2(n_2021),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2477),
.B(n_2095),
.Y(n_2855)
);

O2A1O1Ixp5_ASAP7_75t_L g2856 ( 
.A1(n_2712),
.A2(n_2395),
.B(n_2153),
.C(n_2340),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2748),
.B(n_2150),
.Y(n_2857)
);

BUFx3_ASAP7_75t_L g2858 ( 
.A(n_2563),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2488),
.Y(n_2859)
);

INVxp67_ASAP7_75t_L g2860 ( 
.A(n_2479),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2751),
.B(n_2155),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2751),
.B(n_2159),
.Y(n_2862)
);

AOI21xp5_ASAP7_75t_L g2863 ( 
.A1(n_2548),
.A2(n_2228),
.B(n_2244),
.Y(n_2863)
);

NOR2xp33_ASAP7_75t_L g2864 ( 
.A(n_2569),
.B(n_2029),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_SL g2865 ( 
.A(n_2550),
.B(n_2023),
.Y(n_2865)
);

O2A1O1Ixp5_ASAP7_75t_L g2866 ( 
.A1(n_2557),
.A2(n_2395),
.B(n_2318),
.C(n_2207),
.Y(n_2866)
);

NAND2xp33_ASAP7_75t_L g2867 ( 
.A(n_2589),
.B(n_1725),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2477),
.B(n_2103),
.Y(n_2868)
);

CKINVDCx5p33_ASAP7_75t_R g2869 ( 
.A(n_2601),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2520),
.B(n_2114),
.Y(n_2870)
);

OAI22xp33_ASAP7_75t_L g2871 ( 
.A1(n_2533),
.A2(n_2023),
.B1(n_2018),
.B2(n_2004),
.Y(n_2871)
);

INVx2_ASAP7_75t_SL g2872 ( 
.A(n_2434),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2479),
.B(n_2034),
.Y(n_2873)
);

AOI22xp33_ASAP7_75t_L g2874 ( 
.A1(n_2453),
.A2(n_1899),
.B1(n_1487),
.B2(n_1403),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_SL g2875 ( 
.A(n_2610),
.B(n_1919),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2649),
.B(n_2160),
.Y(n_2876)
);

O2A1O1Ixp33_ASAP7_75t_L g2877 ( 
.A1(n_2569),
.A2(n_1928),
.B(n_1933),
.C(n_1922),
.Y(n_2877)
);

INVxp67_ASAP7_75t_L g2878 ( 
.A(n_2574),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2649),
.B(n_2161),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2697),
.B(n_2162),
.Y(n_2880)
);

NOR2xp33_ASAP7_75t_L g2881 ( 
.A(n_2587),
.B(n_2030),
.Y(n_2881)
);

INVx2_ASAP7_75t_SL g2882 ( 
.A(n_2435),
.Y(n_2882)
);

NOR2xp67_ASAP7_75t_L g2883 ( 
.A(n_2714),
.B(n_1897),
.Y(n_2883)
);

OR2x2_ASAP7_75t_L g2884 ( 
.A(n_2498),
.B(n_2030),
.Y(n_2884)
);

BUFx5_ASAP7_75t_L g2885 ( 
.A(n_2589),
.Y(n_2885)
);

BUFx5_ASAP7_75t_L g2886 ( 
.A(n_2589),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_L g2887 ( 
.A(n_2587),
.B(n_2031),
.Y(n_2887)
);

INVx2_ASAP7_75t_SL g2888 ( 
.A(n_2435),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2521),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2610),
.B(n_1934),
.Y(n_2890)
);

NAND2xp33_ASAP7_75t_L g2891 ( 
.A(n_2619),
.B(n_1728),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_SL g2892 ( 
.A(n_2661),
.B(n_1939),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2697),
.B(n_2163),
.Y(n_2893)
);

INVxp67_ASAP7_75t_L g2894 ( 
.A(n_2599),
.Y(n_2894)
);

OR2x2_ASAP7_75t_L g2895 ( 
.A(n_2529),
.B(n_2031),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2443),
.B(n_1852),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_2410),
.B(n_1852),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2494),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2493),
.B(n_2164),
.Y(n_2899)
);

AOI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2418),
.A2(n_1728),
.B1(n_1948),
.B2(n_1947),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_SL g2901 ( 
.A(n_2661),
.B(n_1951),
.Y(n_2901)
);

NOR2xp33_ASAP7_75t_L g2902 ( 
.A(n_2604),
.B(n_1856),
.Y(n_2902)
);

HB1xp67_ASAP7_75t_L g2903 ( 
.A(n_2526),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2503),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2493),
.B(n_2165),
.Y(n_2905)
);

INVx3_ASAP7_75t_L g2906 ( 
.A(n_2409),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2510),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2492),
.B(n_1927),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2520),
.B(n_2156),
.Y(n_2909)
);

INVxp67_ASAP7_75t_SL g2910 ( 
.A(n_2464),
.Y(n_2910)
);

INVx2_ASAP7_75t_SL g2911 ( 
.A(n_2413),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2519),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2452),
.B(n_1856),
.Y(n_2913)
);

CKINVDCx5p33_ASAP7_75t_R g2914 ( 
.A(n_2536),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2745),
.B(n_2200),
.Y(n_2915)
);

AND2x4_ASAP7_75t_L g2916 ( 
.A(n_2504),
.B(n_2318),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2527),
.Y(n_2917)
);

OAI221xp5_ASAP7_75t_L g2918 ( 
.A1(n_2514),
.A2(n_2020),
.B1(n_2026),
.B2(n_2014),
.C(n_2002),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2528),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2548),
.A2(n_2224),
.B(n_2213),
.Y(n_2920)
);

INVx2_ASAP7_75t_SL g2921 ( 
.A(n_2428),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2511),
.B(n_2168),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_SL g2923 ( 
.A(n_2420),
.B(n_1960),
.Y(n_2923)
);

AOI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2500),
.A2(n_1966),
.B1(n_1970),
.B2(n_1962),
.Y(n_2924)
);

INVx8_ASAP7_75t_L g2925 ( 
.A(n_2475),
.Y(n_2925)
);

NAND2x1_ASAP7_75t_L g2926 ( 
.A(n_2681),
.B(n_2265),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2531),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2511),
.B(n_2173),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2547),
.B(n_2570),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_SL g2930 ( 
.A(n_2452),
.B(n_1972),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2474),
.B(n_1930),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2544),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2547),
.B(n_2176),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2553),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2570),
.B(n_2177),
.Y(n_2935)
);

NOR2xp33_ASAP7_75t_L g2936 ( 
.A(n_2474),
.B(n_1930),
.Y(n_2936)
);

NOR2xp33_ASAP7_75t_L g2937 ( 
.A(n_2408),
.B(n_1974),
.Y(n_2937)
);

O2A1O1Ixp5_ASAP7_75t_L g2938 ( 
.A1(n_2585),
.A2(n_2210),
.B(n_2216),
.C(n_2214),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2581),
.B(n_2178),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2559),
.Y(n_2940)
);

NOR2xp33_ASAP7_75t_SL g2941 ( 
.A(n_2506),
.B(n_1768),
.Y(n_2941)
);

AOI22x1_ASAP7_75t_L g2942 ( 
.A1(n_2710),
.A2(n_1909),
.B1(n_1905),
.B2(n_2126),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2560),
.Y(n_2943)
);

BUFx6f_ASAP7_75t_L g2944 ( 
.A(n_2409),
.Y(n_2944)
);

INVx2_ASAP7_75t_SL g2945 ( 
.A(n_2444),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2538),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_SL g2947 ( 
.A(n_2673),
.B(n_1978),
.Y(n_2947)
);

AOI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2620),
.A2(n_2224),
.B(n_2213),
.Y(n_2948)
);

NOR2xp33_ASAP7_75t_L g2949 ( 
.A(n_2481),
.B(n_1974),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2546),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2552),
.Y(n_2951)
);

INVx3_ASAP7_75t_L g2952 ( 
.A(n_2411),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2581),
.B(n_2464),
.Y(n_2953)
);

BUFx12f_ASAP7_75t_L g2954 ( 
.A(n_2572),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2467),
.B(n_2180),
.Y(n_2955)
);

HB1xp67_ASAP7_75t_L g2956 ( 
.A(n_2530),
.Y(n_2956)
);

BUFx6f_ASAP7_75t_L g2957 ( 
.A(n_2411),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2502),
.B(n_1487),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2564),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2646),
.B(n_1980),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2646),
.B(n_1988),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2565),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2568),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_SL g2964 ( 
.A(n_2504),
.B(n_1927),
.Y(n_2964)
);

NAND2xp33_ASAP7_75t_L g2965 ( 
.A(n_2619),
.B(n_2622),
.Y(n_2965)
);

NOR2xp33_ASAP7_75t_L g2966 ( 
.A(n_2509),
.B(n_2033),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2578),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2583),
.Y(n_2968)
);

AND2x2_ASAP7_75t_L g2969 ( 
.A(n_2415),
.B(n_1927),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2415),
.B(n_1847),
.Y(n_2970)
);

NOR2xp67_ASAP7_75t_L g2971 ( 
.A(n_2677),
.B(n_1768),
.Y(n_2971)
);

CKINVDCx20_ASAP7_75t_R g2972 ( 
.A(n_2532),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2603),
.Y(n_2973)
);

AOI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_2467),
.A2(n_1884),
.B1(n_1765),
.B2(n_2035),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2607),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2473),
.B(n_1857),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2473),
.B(n_1857),
.Y(n_2977)
);

OR2x6_ASAP7_75t_L g2978 ( 
.A(n_2638),
.B(n_2556),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2461),
.B(n_1407),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2554),
.Y(n_2980)
);

OR2x2_ASAP7_75t_L g2981 ( 
.A(n_2597),
.B(n_1865),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2737),
.B(n_1857),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2650),
.Y(n_2983)
);

AOI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2482),
.A2(n_1884),
.B1(n_1765),
.B2(n_2633),
.Y(n_2984)
);

INVxp67_ASAP7_75t_SL g2985 ( 
.A(n_2482),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2566),
.Y(n_2986)
);

INVxp67_ASAP7_75t_L g2987 ( 
.A(n_2626),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2567),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2737),
.B(n_2201),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2613),
.B(n_1411),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2652),
.Y(n_2991)
);

INVx8_ASAP7_75t_L g2992 ( 
.A(n_2475),
.Y(n_2992)
);

AOI22x1_ASAP7_75t_L g2993 ( 
.A1(n_2710),
.A2(n_2126),
.B1(n_2229),
.B2(n_2183),
.Y(n_2993)
);

NOR3xp33_ASAP7_75t_L g2994 ( 
.A(n_2713),
.B(n_2018),
.C(n_2004),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2540),
.B(n_2004),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2573),
.Y(n_2996)
);

BUFx6f_ASAP7_75t_L g2997 ( 
.A(n_2411),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2653),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2696),
.B(n_1895),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2696),
.B(n_1903),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_SL g3001 ( 
.A(n_2525),
.B(n_1765),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2525),
.B(n_1884),
.Y(n_3002)
);

OAI22xp33_ASAP7_75t_L g3003 ( 
.A1(n_2730),
.A2(n_2018),
.B1(n_2036),
.B2(n_2037),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2611),
.Y(n_3004)
);

INVx6_ASAP7_75t_L g3005 ( 
.A(n_2459),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2655),
.Y(n_3006)
);

AOI22xp33_ASAP7_75t_L g3007 ( 
.A1(n_2523),
.A2(n_1411),
.B1(n_1417),
.B2(n_1413),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2556),
.B(n_1914),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2615),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2693),
.B(n_2037),
.Y(n_3010)
);

NOR2x1p5_ASAP7_75t_L g3011 ( 
.A(n_2472),
.B(n_2036),
.Y(n_3011)
);

BUFx2_ASAP7_75t_L g3012 ( 
.A(n_2556),
.Y(n_3012)
);

OAI22xp33_ASAP7_75t_L g3013 ( 
.A1(n_2695),
.A2(n_2036),
.B1(n_2037),
.B2(n_2039),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2660),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2708),
.B(n_1906),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2670),
.Y(n_3016)
);

BUFx6f_ASAP7_75t_L g3017 ( 
.A(n_2411),
.Y(n_3017)
);

AOI22xp33_ASAP7_75t_L g3018 ( 
.A1(n_2523),
.A2(n_1413),
.B1(n_1420),
.B2(n_1417),
.Y(n_3018)
);

NOR2xp33_ASAP7_75t_L g3019 ( 
.A(n_2738),
.B(n_1420),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2708),
.B(n_2261),
.Y(n_3020)
);

OAI22xp5_ASAP7_75t_L g3021 ( 
.A1(n_2617),
.A2(n_2142),
.B1(n_2183),
.B2(n_2184),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2675),
.Y(n_3022)
);

OR2x6_ASAP7_75t_L g3023 ( 
.A(n_2638),
.B(n_2037),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2628),
.Y(n_3024)
);

AND2x2_ASAP7_75t_SL g3025 ( 
.A(n_2524),
.B(n_1806),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_SL g3026 ( 
.A(n_2491),
.B(n_2347),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2662),
.B(n_2186),
.Y(n_3027)
);

INVxp67_ASAP7_75t_L g3028 ( 
.A(n_2643),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_L g3029 ( 
.A1(n_2523),
.A2(n_1423),
.B1(n_1432),
.B2(n_1428),
.Y(n_3029)
);

CKINVDCx5p33_ASAP7_75t_R g3030 ( 
.A(n_2580),
.Y(n_3030)
);

INVx2_ASAP7_75t_SL g3031 ( 
.A(n_2476),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2400),
.B(n_2187),
.Y(n_3032)
);

AOI22xp33_ASAP7_75t_L g3033 ( 
.A1(n_2676),
.A2(n_1423),
.B1(n_1432),
.B2(n_1428),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2630),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_SL g3035 ( 
.A(n_2491),
.B(n_2145),
.Y(n_3035)
);

HB1xp67_ASAP7_75t_L g3036 ( 
.A(n_2709),
.Y(n_3036)
);

AOI22xp33_ASAP7_75t_L g3037 ( 
.A1(n_2641),
.A2(n_1441),
.B1(n_2657),
.B2(n_2727),
.Y(n_3037)
);

NAND2x1_ASAP7_75t_L g3038 ( 
.A(n_2681),
.B(n_2265),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_SL g3039 ( 
.A(n_2496),
.B(n_1885),
.Y(n_3039)
);

BUFx12f_ASAP7_75t_L g3040 ( 
.A(n_2722),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_SL g3041 ( 
.A(n_2496),
.B(n_2265),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2635),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_SL g3043 ( 
.A(n_2618),
.B(n_2271),
.Y(n_3043)
);

INVx2_ASAP7_75t_SL g3044 ( 
.A(n_2490),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2400),
.B(n_2190),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2618),
.B(n_1441),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2678),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_SL g3048 ( 
.A(n_2750),
.B(n_2271),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2684),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_2750),
.B(n_2271),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_L g3051 ( 
.A(n_2633),
.B(n_1810),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2694),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2617),
.B(n_2631),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_SL g3054 ( 
.A(n_2631),
.B(n_2641),
.Y(n_3054)
);

INVx1_ASAP7_75t_SL g3055 ( 
.A(n_2727),
.Y(n_3055)
);

INVxp67_ASAP7_75t_L g3056 ( 
.A(n_2739),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2400),
.B(n_2191),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2705),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_SL g3059 ( 
.A(n_2657),
.B(n_2284),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2723),
.B(n_1823),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2679),
.Y(n_3061)
);

BUFx6f_ASAP7_75t_SL g3062 ( 
.A(n_2475),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_SL g3063 ( 
.A(n_2459),
.B(n_2284),
.Y(n_3063)
);

NOR2xp33_ASAP7_75t_L g3064 ( 
.A(n_2731),
.B(n_1896),
.Y(n_3064)
);

NOR2xp33_ASAP7_75t_L g3065 ( 
.A(n_2731),
.B(n_1902),
.Y(n_3065)
);

NOR2xp33_ASAP7_75t_L g3066 ( 
.A(n_2740),
.B(n_1926),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2680),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_2739),
.B(n_2284),
.Y(n_3068)
);

NAND3xp33_ASAP7_75t_L g3069 ( 
.A(n_2740),
.B(n_1926),
.C(n_2383),
.Y(n_3069)
);

AOI22xp5_ASAP7_75t_L g3070 ( 
.A1(n_2400),
.A2(n_2167),
.B1(n_1926),
.B2(n_1699),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_SL g3071 ( 
.A(n_2659),
.B(n_2593),
.Y(n_3071)
);

INVxp67_ASAP7_75t_L g3072 ( 
.A(n_2896),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2764),
.B(n_2662),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2768),
.B(n_2686),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2763),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_2761),
.B(n_884),
.Y(n_3076)
);

INVx5_ASAP7_75t_L g3077 ( 
.A(n_2925),
.Y(n_3077)
);

NOR2xp33_ASAP7_75t_L g3078 ( 
.A(n_2779),
.B(n_2424),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_2788),
.B(n_2469),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2816),
.B(n_2593),
.Y(n_3080)
);

NOR2x1p5_ASAP7_75t_L g3081 ( 
.A(n_2869),
.B(n_2704),
.Y(n_3081)
);

NAND3xp33_ASAP7_75t_SL g3082 ( 
.A(n_2758),
.B(n_2000),
.C(n_717),
.Y(n_3082)
);

INVx3_ASAP7_75t_L g3083 ( 
.A(n_2925),
.Y(n_3083)
);

OAI22xp33_ASAP7_75t_L g3084 ( 
.A1(n_2765),
.A2(n_2638),
.B1(n_2703),
.B2(n_2755),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2778),
.B(n_979),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2787),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2797),
.Y(n_3087)
);

INVxp67_ASAP7_75t_SL g3088 ( 
.A(n_2835),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2836),
.B(n_2929),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2799),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2773),
.Y(n_3091)
);

INVx2_ASAP7_75t_SL g3092 ( 
.A(n_2858),
.Y(n_3092)
);

BUFx6f_ASAP7_75t_L g3093 ( 
.A(n_2925),
.Y(n_3093)
);

AOI22xp33_ASAP7_75t_L g3094 ( 
.A1(n_3007),
.A2(n_2400),
.B1(n_1699),
.B2(n_2422),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2776),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2785),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2786),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2804),
.Y(n_3098)
);

OR2x6_ASAP7_75t_L g3099 ( 
.A(n_2992),
.B(n_2781),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2836),
.B(n_2422),
.Y(n_3100)
);

INVx3_ASAP7_75t_L g3101 ( 
.A(n_2992),
.Y(n_3101)
);

NOR2x1_ASAP7_75t_L g3102 ( 
.A(n_2972),
.B(n_2781),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2801),
.B(n_3065),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2759),
.B(n_2690),
.Y(n_3104)
);

NOR3xp33_ASAP7_75t_SL g3105 ( 
.A(n_3030),
.B(n_721),
.C(n_715),
.Y(n_3105)
);

AOI22xp33_ASAP7_75t_L g3106 ( 
.A1(n_3018),
.A2(n_1699),
.B1(n_2429),
.B2(n_2450),
.Y(n_3106)
);

AND2x6_ASAP7_75t_L g3107 ( 
.A(n_3062),
.B(n_2447),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2793),
.B(n_2698),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2807),
.Y(n_3109)
);

INVx5_ASAP7_75t_L g3110 ( 
.A(n_2992),
.Y(n_3110)
);

INVx1_ASAP7_75t_SL g3111 ( 
.A(n_2791),
.Y(n_3111)
);

AOI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_3064),
.A2(n_2475),
.B1(n_2499),
.B2(n_2465),
.Y(n_3112)
);

AND2x4_ASAP7_75t_L g3113 ( 
.A(n_2978),
.B(n_2614),
.Y(n_3113)
);

AND2x2_ASAP7_75t_SL g3114 ( 
.A(n_3025),
.B(n_2524),
.Y(n_3114)
);

NAND3xp33_ASAP7_75t_L g3115 ( 
.A(n_2838),
.B(n_2486),
.C(n_2302),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2796),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2810),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2812),
.Y(n_3118)
);

BUFx6f_ASAP7_75t_L g3119 ( 
.A(n_2802),
.Y(n_3119)
);

BUFx2_ASAP7_75t_L g3120 ( 
.A(n_2903),
.Y(n_3120)
);

OAI22xp5_ASAP7_75t_SL g3121 ( 
.A1(n_2847),
.A2(n_873),
.B1(n_878),
.B2(n_870),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2825),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2841),
.Y(n_3123)
);

BUFx12f_ASAP7_75t_L g3124 ( 
.A(n_2852),
.Y(n_3124)
);

NOR2xp33_ASAP7_75t_L g3125 ( 
.A(n_3066),
.B(n_2897),
.Y(n_3125)
);

OAI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_2827),
.A2(n_2719),
.B1(n_2725),
.B2(n_2704),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_SL g3127 ( 
.A(n_2913),
.B(n_2593),
.Y(n_3127)
);

O2A1O1Ixp33_ASAP7_75t_L g3128 ( 
.A1(n_2830),
.A2(n_2439),
.B(n_2756),
.C(n_2747),
.Y(n_3128)
);

BUFx3_ASAP7_75t_L g3129 ( 
.A(n_2954),
.Y(n_3129)
);

NAND2x1p5_ASAP7_75t_L g3130 ( 
.A(n_2945),
.B(n_2412),
.Y(n_3130)
);

NOR2x2_ASAP7_75t_L g3131 ( 
.A(n_2781),
.B(n_2834),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_3051),
.B(n_2719),
.Y(n_3132)
);

AOI221xp5_ASAP7_75t_SL g3133 ( 
.A1(n_2760),
.A2(n_2621),
.B1(n_2728),
.B2(n_2733),
.C(n_2725),
.Y(n_3133)
);

AOI21xp5_ASAP7_75t_L g3134 ( 
.A1(n_2965),
.A2(n_2621),
.B(n_2636),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_3055),
.B(n_2728),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2848),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2814),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_SL g3138 ( 
.A(n_2931),
.B(n_2593),
.Y(n_3138)
);

INVx2_ASAP7_75t_SL g3139 ( 
.A(n_3011),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2889),
.Y(n_3140)
);

AOI22xp33_ASAP7_75t_L g3141 ( 
.A1(n_3029),
.A2(n_2429),
.B1(n_2450),
.B2(n_2195),
.Y(n_3141)
);

BUFx6f_ASAP7_75t_L g3142 ( 
.A(n_2802),
.Y(n_3142)
);

AND2x2_ASAP7_75t_L g3143 ( 
.A(n_3037),
.B(n_2873),
.Y(n_3143)
);

O2A1O1Ixp33_ASAP7_75t_L g3144 ( 
.A1(n_2875),
.A2(n_2733),
.B(n_2512),
.C(n_2535),
.Y(n_3144)
);

BUFx2_ASAP7_75t_L g3145 ( 
.A(n_2956),
.Y(n_3145)
);

INVxp67_ASAP7_75t_L g3146 ( 
.A(n_2864),
.Y(n_3146)
);

AOI22xp5_ASAP7_75t_L g3147 ( 
.A1(n_2902),
.A2(n_2475),
.B1(n_2499),
.B2(n_2465),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_SL g3148 ( 
.A(n_2936),
.B(n_2637),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_2917),
.Y(n_3149)
);

INVx3_ASAP7_75t_L g3150 ( 
.A(n_3062),
.Y(n_3150)
);

BUFx2_ASAP7_75t_L g3151 ( 
.A(n_2766),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2815),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2837),
.B(n_2499),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2833),
.Y(n_3154)
);

NAND2x2_ASAP7_75t_L g3155 ( 
.A(n_2884),
.B(n_2671),
.Y(n_3155)
);

NOR2xp33_ASAP7_75t_L g3156 ( 
.A(n_2895),
.B(n_2501),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2851),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2853),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2860),
.B(n_2499),
.Y(n_3159)
);

INVxp67_ASAP7_75t_L g3160 ( 
.A(n_2958),
.Y(n_3160)
);

A2O1A1Ixp33_ASAP7_75t_L g3161 ( 
.A1(n_2821),
.A2(n_2755),
.B(n_2685),
.C(n_2659),
.Y(n_3161)
);

AND2x4_ASAP7_75t_L g3162 ( 
.A(n_2978),
.B(n_2614),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2946),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2950),
.Y(n_3164)
);

NAND2x1p5_ASAP7_75t_L g3165 ( 
.A(n_2792),
.B(n_2412),
.Y(n_3165)
);

AND2x4_ASAP7_75t_L g3166 ( 
.A(n_2978),
.B(n_2614),
.Y(n_3166)
);

AOI22xp5_ASAP7_75t_L g3167 ( 
.A1(n_2890),
.A2(n_2499),
.B1(n_2465),
.B2(n_2715),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2859),
.Y(n_3168)
);

AOI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_2937),
.A2(n_2465),
.B1(n_2715),
.B2(n_2622),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2898),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2904),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2909),
.B(n_2757),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2907),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_3046),
.B(n_979),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_R g3175 ( 
.A(n_2914),
.B(n_2619),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_SL g3176 ( 
.A(n_2772),
.B(n_2637),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2908),
.B(n_2405),
.Y(n_3177)
);

CKINVDCx5p33_ASAP7_75t_R g3178 ( 
.A(n_3040),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_L g3179 ( 
.A(n_2941),
.B(n_2707),
.Y(n_3179)
);

BUFx4f_ASAP7_75t_L g3180 ( 
.A(n_2802),
.Y(n_3180)
);

NAND2x1p5_ASAP7_75t_L g3181 ( 
.A(n_2800),
.B(n_2412),
.Y(n_3181)
);

A2O1A1Ixp33_ASAP7_75t_L g3182 ( 
.A1(n_2999),
.A2(n_3015),
.B(n_3000),
.C(n_2823),
.Y(n_3182)
);

AND2x2_ASAP7_75t_L g3183 ( 
.A(n_3019),
.B(n_979),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_SL g3184 ( 
.A(n_2795),
.B(n_2637),
.Y(n_3184)
);

INVx5_ASAP7_75t_L g3185 ( 
.A(n_2834),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2912),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2919),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2855),
.B(n_2724),
.Y(n_3188)
);

NOR2xp33_ASAP7_75t_R g3189 ( 
.A(n_2817),
.B(n_2619),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_SL g3190 ( 
.A(n_2803),
.B(n_2637),
.Y(n_3190)
);

INVx2_ASAP7_75t_SL g3191 ( 
.A(n_2834),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_L g3192 ( 
.A(n_2829),
.B(n_2588),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2868),
.B(n_2734),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2927),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2932),
.Y(n_3195)
);

NOR2x1p5_ASAP7_75t_L g3196 ( 
.A(n_3069),
.B(n_2407),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2949),
.B(n_2742),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_SL g3198 ( 
.A(n_2808),
.B(n_2447),
.Y(n_3198)
);

AND2x4_ASAP7_75t_L g3199 ( 
.A(n_3023),
.B(n_2634),
.Y(n_3199)
);

BUFx3_ASAP7_75t_L g3200 ( 
.A(n_2911),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2771),
.A2(n_2774),
.B(n_2767),
.Y(n_3201)
);

OR2x2_ASAP7_75t_L g3202 ( 
.A(n_2775),
.B(n_2416),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_2951),
.Y(n_3203)
);

AOI22xp5_ASAP7_75t_L g3204 ( 
.A1(n_3060),
.A2(n_2465),
.B1(n_2622),
.B2(n_2619),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_SL g3205 ( 
.A(n_2871),
.B(n_2513),
.Y(n_3205)
);

NAND2x1p5_ASAP7_75t_L g3206 ( 
.A(n_3031),
.B(n_2470),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_SL g3207 ( 
.A(n_3003),
.B(n_2513),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2934),
.Y(n_3208)
);

INVx3_ASAP7_75t_L g3209 ( 
.A(n_2842),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_L g3210 ( 
.A(n_2990),
.B(n_2749),
.Y(n_3210)
);

NOR2x1_ASAP7_75t_R g3211 ( 
.A(n_3012),
.B(n_2470),
.Y(n_3211)
);

AOI22xp5_ASAP7_75t_L g3212 ( 
.A1(n_2780),
.A2(n_2622),
.B1(n_2627),
.B2(n_2685),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_SL g3213 ( 
.A(n_2822),
.B(n_2826),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2940),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_SL g3215 ( 
.A(n_2828),
.B(n_2522),
.Y(n_3215)
);

BUFx6f_ASAP7_75t_L g3216 ( 
.A(n_2789),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2980),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2986),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2929),
.B(n_2427),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2943),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2959),
.Y(n_3221)
);

NAND3xp33_ASAP7_75t_L g3222 ( 
.A(n_2784),
.B(n_2338),
.C(n_2307),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_2881),
.B(n_2717),
.Y(n_3223)
);

AND2x4_ASAP7_75t_L g3224 ( 
.A(n_3023),
.B(n_2916),
.Y(n_3224)
);

HB1xp67_ASAP7_75t_L g3225 ( 
.A(n_2878),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2962),
.Y(n_3226)
);

BUFx2_ASAP7_75t_L g3227 ( 
.A(n_2894),
.Y(n_3227)
);

BUFx12f_ASAP7_75t_L g3228 ( 
.A(n_2783),
.Y(n_3228)
);

XNOR2xp5_ASAP7_75t_L g3229 ( 
.A(n_3033),
.B(n_2648),
.Y(n_3229)
);

AND2x4_ASAP7_75t_L g3230 ( 
.A(n_3023),
.B(n_2634),
.Y(n_3230)
);

HB1xp67_ASAP7_75t_L g3231 ( 
.A(n_3036),
.Y(n_3231)
);

AOI22xp33_ASAP7_75t_SL g3232 ( 
.A1(n_2979),
.A2(n_2666),
.B1(n_2627),
.B2(n_2622),
.Y(n_3232)
);

AND2x4_ASAP7_75t_L g3233 ( 
.A(n_2916),
.B(n_2634),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_SL g3234 ( 
.A(n_3013),
.B(n_2522),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_2771),
.B(n_2430),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2988),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2774),
.B(n_2431),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2996),
.Y(n_3238)
);

BUFx3_ASAP7_75t_L g3239 ( 
.A(n_2921),
.Y(n_3239)
);

AOI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_2887),
.A2(n_2627),
.B1(n_2632),
.B2(n_2575),
.Y(n_3240)
);

AND2x4_ASAP7_75t_L g3241 ( 
.A(n_3044),
.B(n_2642),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_3020),
.B(n_2433),
.Y(n_3242)
);

NOR2x2_ASAP7_75t_L g3243 ( 
.A(n_2874),
.B(n_620),
.Y(n_3243)
);

AND2x4_ASAP7_75t_L g3244 ( 
.A(n_2971),
.B(n_2642),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_2782),
.B(n_2700),
.Y(n_3245)
);

INVxp67_ASAP7_75t_L g3246 ( 
.A(n_2918),
.Y(n_3246)
);

AND2x4_ASAP7_75t_L g3247 ( 
.A(n_3056),
.B(n_2642),
.Y(n_3247)
);

AOI22xp33_ASAP7_75t_L g3248 ( 
.A1(n_2849),
.A2(n_2197),
.B1(n_2202),
.B2(n_2194),
.Y(n_3248)
);

AOI22xp5_ASAP7_75t_L g3249 ( 
.A1(n_3053),
.A2(n_2627),
.B1(n_2632),
.B2(n_2575),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2870),
.B(n_2720),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_SL g3251 ( 
.A(n_2953),
.B(n_2699),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2963),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_2967),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_2762),
.A2(n_2767),
.B(n_2863),
.Y(n_3254)
);

CKINVDCx5p33_ASAP7_75t_R g3255 ( 
.A(n_2840),
.Y(n_3255)
);

OR2x2_ASAP7_75t_SL g3256 ( 
.A(n_2981),
.B(n_887),
.Y(n_3256)
);

O2A1O1Ixp5_ASAP7_75t_L g3257 ( 
.A1(n_2930),
.A2(n_2683),
.B(n_2654),
.C(n_2577),
.Y(n_3257)
);

AND2x4_ASAP7_75t_SL g3258 ( 
.A(n_2789),
.B(n_2699),
.Y(n_3258)
);

BUFx2_ASAP7_75t_L g3259 ( 
.A(n_2995),
.Y(n_3259)
);

AOI22xp33_ASAP7_75t_L g3260 ( 
.A1(n_2982),
.A2(n_2204),
.B1(n_2209),
.B2(n_2203),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2968),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3004),
.Y(n_3262)
);

CKINVDCx6p67_ASAP7_75t_R g3263 ( 
.A(n_2790),
.Y(n_3263)
);

BUFx6f_ASAP7_75t_L g3264 ( 
.A(n_2789),
.Y(n_3264)
);

INVx3_ASAP7_75t_L g3265 ( 
.A(n_2842),
.Y(n_3265)
);

INVxp67_ASAP7_75t_L g3266 ( 
.A(n_2966),
.Y(n_3266)
);

INVx4_ASAP7_75t_L g3267 ( 
.A(n_2944),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_2854),
.A2(n_3035),
.B1(n_2969),
.B2(n_3002),
.Y(n_3268)
);

INVx2_ASAP7_75t_SL g3269 ( 
.A(n_2872),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2973),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2975),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_2989),
.B(n_2732),
.Y(n_3272)
);

NOR3xp33_ASAP7_75t_L g3273 ( 
.A(n_2994),
.B(n_878),
.C(n_873),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_SL g3274 ( 
.A(n_2953),
.B(n_2699),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_2970),
.B(n_2752),
.Y(n_3275)
);

INVx2_ASAP7_75t_L g3276 ( 
.A(n_3009),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_2976),
.B(n_2706),
.Y(n_3277)
);

CKINVDCx20_ASAP7_75t_R g3278 ( 
.A(n_2900),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2977),
.B(n_2212),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2983),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2991),
.Y(n_3281)
);

NOR2x2_ASAP7_75t_L g3282 ( 
.A(n_2809),
.B(n_620),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2998),
.Y(n_3283)
);

BUFx3_ASAP7_75t_L g3284 ( 
.A(n_2882),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3006),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_SL g3286 ( 
.A(n_2885),
.B(n_2470),
.Y(n_3286)
);

BUFx3_ASAP7_75t_L g3287 ( 
.A(n_2888),
.Y(n_3287)
);

AND2x4_ASAP7_75t_L g3288 ( 
.A(n_2964),
.B(n_2691),
.Y(n_3288)
);

INVx2_ASAP7_75t_SL g3289 ( 
.A(n_3005),
.Y(n_3289)
);

NOR2xp33_ASAP7_75t_L g3290 ( 
.A(n_2987),
.B(n_2716),
.Y(n_3290)
);

BUFx6f_ASAP7_75t_L g3291 ( 
.A(n_2944),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3014),
.Y(n_3292)
);

OAI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_2782),
.A2(n_2220),
.B1(n_2230),
.B2(n_2218),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_3001),
.A2(n_2236),
.B1(n_2239),
.B2(n_2233),
.Y(n_3294)
);

BUFx2_ASAP7_75t_L g3295 ( 
.A(n_3028),
.Y(n_3295)
);

AOI22xp33_ASAP7_75t_L g3296 ( 
.A1(n_3070),
.A2(n_2240),
.B1(n_2086),
.B2(n_2088),
.Y(n_3296)
);

INVxp67_ASAP7_75t_L g3297 ( 
.A(n_2923),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_3008),
.B(n_979),
.Y(n_3298)
);

AND2x4_ASAP7_75t_L g3299 ( 
.A(n_3071),
.B(n_2691),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_2974),
.B(n_1288),
.Y(n_3300)
);

INVx2_ASAP7_75t_SL g3301 ( 
.A(n_3005),
.Y(n_3301)
);

NOR2xp33_ASAP7_75t_R g3302 ( 
.A(n_2813),
.B(n_2627),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_2915),
.B(n_2689),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3024),
.Y(n_3304)
);

INVx3_ASAP7_75t_L g3305 ( 
.A(n_2770),
.Y(n_3305)
);

BUFx2_ASAP7_75t_L g3306 ( 
.A(n_2944),
.Y(n_3306)
);

NOR2x1p5_ASAP7_75t_L g3307 ( 
.A(n_2770),
.B(n_2407),
.Y(n_3307)
);

INVx3_ASAP7_75t_L g3308 ( 
.A(n_2806),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_2960),
.B(n_2689),
.Y(n_3309)
);

BUFx6f_ASAP7_75t_L g3310 ( 
.A(n_2957),
.Y(n_3310)
);

OR2x2_ASAP7_75t_L g3311 ( 
.A(n_2961),
.B(n_3016),
.Y(n_3311)
);

NAND2x1p5_ASAP7_75t_L g3312 ( 
.A(n_2957),
.B(n_2539),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_SL g3313 ( 
.A(n_3125),
.B(n_3021),
.Y(n_3313)
);

NAND2xp33_ASAP7_75t_SL g3314 ( 
.A(n_3175),
.B(n_2806),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_3132),
.B(n_3021),
.Y(n_3315)
);

NAND2xp33_ASAP7_75t_SL g3316 ( 
.A(n_3189),
.B(n_2947),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_SL g3317 ( 
.A(n_3074),
.B(n_2984),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_SL g3318 ( 
.A(n_3223),
.B(n_2883),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_SL g3319 ( 
.A(n_3112),
.B(n_2769),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_SL g3320 ( 
.A(n_3112),
.B(n_2831),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_SL g3321 ( 
.A(n_3073),
.B(n_2831),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_SL g3322 ( 
.A(n_3147),
.B(n_2760),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_SL g3323 ( 
.A(n_3147),
.B(n_2924),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_3204),
.B(n_2846),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_3204),
.B(n_2846),
.Y(n_3325)
);

NAND2xp33_ASAP7_75t_SL g3326 ( 
.A(n_3302),
.B(n_2957),
.Y(n_3326)
);

NAND2xp33_ASAP7_75t_SL g3327 ( 
.A(n_3278),
.B(n_2997),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_SL g3328 ( 
.A(n_3232),
.B(n_2850),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_SL g3329 ( 
.A(n_3240),
.B(n_2850),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_3240),
.B(n_2857),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_SL g3331 ( 
.A(n_3169),
.B(n_2857),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3089),
.B(n_3266),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_SL g3333 ( 
.A(n_3169),
.B(n_2861),
.Y(n_3333)
);

AND2x2_ASAP7_75t_L g3334 ( 
.A(n_3103),
.B(n_3022),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_SL g3335 ( 
.A(n_3197),
.B(n_2861),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_SL g3336 ( 
.A(n_3078),
.B(n_2862),
.Y(n_3336)
);

NAND2xp33_ASAP7_75t_SL g3337 ( 
.A(n_3307),
.B(n_2997),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_SL g3338 ( 
.A(n_3210),
.B(n_2862),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_SL g3339 ( 
.A(n_3089),
.B(n_2885),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_SL g3340 ( 
.A(n_3167),
.B(n_3309),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_SL g3341 ( 
.A(n_3167),
.B(n_2885),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_SL g3342 ( 
.A(n_3084),
.B(n_2885),
.Y(n_3342)
);

AND2x4_ASAP7_75t_L g3343 ( 
.A(n_3113),
.B(n_3054),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3213),
.B(n_3047),
.Y(n_3344)
);

NAND2xp33_ASAP7_75t_SL g3345 ( 
.A(n_3081),
.B(n_2997),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3108),
.B(n_3061),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_SL g3347 ( 
.A(n_3079),
.B(n_2885),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_3182),
.B(n_2885),
.Y(n_3348)
);

NAND2xp33_ASAP7_75t_SL g3349 ( 
.A(n_3255),
.B(n_3017),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3085),
.B(n_3143),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_SL g3351 ( 
.A(n_3146),
.B(n_2886),
.Y(n_3351)
);

NAND2xp33_ASAP7_75t_SL g3352 ( 
.A(n_3076),
.B(n_3017),
.Y(n_3352)
);

NAND2xp33_ASAP7_75t_SL g3353 ( 
.A(n_3202),
.B(n_3017),
.Y(n_3353)
);

AND2x4_ASAP7_75t_L g3354 ( 
.A(n_3113),
.B(n_2820),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_SL g3355 ( 
.A(n_3246),
.B(n_2886),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_3104),
.B(n_2886),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_SL g3357 ( 
.A(n_3179),
.B(n_2886),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_SL g3358 ( 
.A(n_3180),
.B(n_2886),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_3180),
.B(n_2886),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3298),
.B(n_3067),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_SL g3361 ( 
.A(n_3172),
.B(n_2876),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_3188),
.B(n_2876),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3303),
.B(n_2879),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_3111),
.B(n_2879),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_3193),
.B(n_2880),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_SL g3366 ( 
.A(n_3250),
.B(n_2880),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3111),
.B(n_2893),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_3119),
.B(n_2893),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_SL g3369 ( 
.A(n_3119),
.B(n_2762),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_SL g3370 ( 
.A(n_3119),
.B(n_2839),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3088),
.B(n_3027),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_SL g3372 ( 
.A(n_3142),
.B(n_2899),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_SL g3373 ( 
.A(n_3142),
.B(n_2899),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3311),
.B(n_3272),
.Y(n_3374)
);

NAND2xp33_ASAP7_75t_SL g3375 ( 
.A(n_3105),
.B(n_2892),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_SL g3376 ( 
.A(n_3142),
.B(n_2905),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_SL g3377 ( 
.A(n_3242),
.B(n_2905),
.Y(n_3377)
);

NAND2xp33_ASAP7_75t_SL g3378 ( 
.A(n_3178),
.B(n_2901),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_SL g3379 ( 
.A(n_3242),
.B(n_2922),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_SL g3380 ( 
.A(n_3114),
.B(n_3185),
.Y(n_3380)
);

NAND2xp33_ASAP7_75t_SL g3381 ( 
.A(n_3093),
.B(n_2843),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_SL g3382 ( 
.A(n_3185),
.B(n_2922),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_3185),
.B(n_2928),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_SL g3384 ( 
.A(n_3296),
.B(n_2928),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_SL g3385 ( 
.A(n_3219),
.B(n_2933),
.Y(n_3385)
);

AND2x4_ASAP7_75t_L g3386 ( 
.A(n_3162),
.B(n_2820),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3120),
.B(n_2844),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_3219),
.B(n_2933),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_SL g3389 ( 
.A(n_3100),
.B(n_2935),
.Y(n_3389)
);

AND2x2_ASAP7_75t_L g3390 ( 
.A(n_3259),
.B(n_2798),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_SL g3391 ( 
.A(n_3100),
.B(n_2935),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_3115),
.B(n_2939),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_3115),
.B(n_2939),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_SL g3394 ( 
.A(n_3127),
.B(n_2818),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_SL g3395 ( 
.A(n_3138),
.B(n_2819),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_SL g3396 ( 
.A(n_3148),
.B(n_2955),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_SL g3397 ( 
.A(n_3212),
.B(n_2955),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_SL g3398 ( 
.A(n_3212),
.B(n_2726),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_SL g3399 ( 
.A(n_3249),
.B(n_2726),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_SL g3400 ( 
.A(n_3249),
.B(n_2726),
.Y(n_3400)
);

NAND2xp33_ASAP7_75t_SL g3401 ( 
.A(n_3093),
.B(n_2865),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3145),
.B(n_3010),
.Y(n_3402)
);

AND2x4_ASAP7_75t_L g3403 ( 
.A(n_3162),
.B(n_2906),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_SL g3404 ( 
.A(n_3300),
.B(n_2726),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_SL g3405 ( 
.A(n_3192),
.B(n_2877),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3151),
.B(n_2794),
.Y(n_3406)
);

AND2x4_ASAP7_75t_L g3407 ( 
.A(n_3166),
.B(n_2906),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_SL g3408 ( 
.A(n_3222),
.B(n_2426),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3174),
.B(n_3072),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3177),
.B(n_2910),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_SL g3411 ( 
.A(n_3222),
.B(n_2426),
.Y(n_3411)
);

NAND2xp33_ASAP7_75t_SL g3412 ( 
.A(n_3093),
.B(n_2824),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_SL g3413 ( 
.A(n_3133),
.B(n_2426),
.Y(n_3413)
);

AND2x2_ASAP7_75t_L g3414 ( 
.A(n_3183),
.B(n_2832),
.Y(n_3414)
);

AND2x4_ASAP7_75t_L g3415 ( 
.A(n_3166),
.B(n_2952),
.Y(n_3415)
);

NAND2xp33_ASAP7_75t_SL g3416 ( 
.A(n_3121),
.B(n_2926),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_SL g3417 ( 
.A(n_3133),
.B(n_2426),
.Y(n_3417)
);

NAND2xp33_ASAP7_75t_SL g3418 ( 
.A(n_3121),
.B(n_3038),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_SL g3419 ( 
.A(n_3234),
.B(n_2454),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_SL g3420 ( 
.A(n_3290),
.B(n_2454),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_SL g3421 ( 
.A(n_3245),
.B(n_2454),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_3245),
.B(n_2454),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3160),
.B(n_2985),
.Y(n_3423)
);

AND2x4_ASAP7_75t_L g3424 ( 
.A(n_3099),
.B(n_2952),
.Y(n_3424)
);

NAND2xp33_ASAP7_75t_SL g3425 ( 
.A(n_3305),
.B(n_2716),
.Y(n_3425)
);

NAND2xp33_ASAP7_75t_SL g3426 ( 
.A(n_3305),
.B(n_2845),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3135),
.B(n_3034),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3275),
.B(n_3042),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_3153),
.B(n_2460),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_SL g3430 ( 
.A(n_3159),
.B(n_3235),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_SL g3431 ( 
.A(n_3235),
.B(n_2460),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_SL g3432 ( 
.A(n_3237),
.B(n_2460),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_SL g3433 ( 
.A(n_3237),
.B(n_2460),
.Y(n_3433)
);

NAND2xp33_ASAP7_75t_SL g3434 ( 
.A(n_3308),
.B(n_2867),
.Y(n_3434)
);

NAND2xp33_ASAP7_75t_SL g3435 ( 
.A(n_3308),
.B(n_2891),
.Y(n_3435)
);

AND2x4_ASAP7_75t_L g3436 ( 
.A(n_3099),
.B(n_3032),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_3077),
.B(n_2471),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_SL g3438 ( 
.A(n_3077),
.B(n_2471),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_3077),
.B(n_2471),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_SL g3440 ( 
.A(n_3110),
.B(n_2471),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_SL g3441 ( 
.A(n_3110),
.B(n_2487),
.Y(n_3441)
);

XNOR2x2_ASAP7_75t_L g3442 ( 
.A(n_3229),
.B(n_3026),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3277),
.B(n_3049),
.Y(n_3443)
);

NAND2xp33_ASAP7_75t_SL g3444 ( 
.A(n_3269),
.B(n_3048),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_SL g3445 ( 
.A(n_3110),
.B(n_2487),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3156),
.B(n_3052),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_SL g3447 ( 
.A(n_3216),
.B(n_2487),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_SL g3448 ( 
.A(n_3216),
.B(n_2487),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_3216),
.B(n_2505),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_3264),
.B(n_2505),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_SL g3451 ( 
.A(n_3264),
.B(n_2505),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_SL g3452 ( 
.A(n_3264),
.B(n_2505),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3231),
.B(n_3058),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_SL g3454 ( 
.A(n_3291),
.B(n_2516),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_SL g3455 ( 
.A(n_3291),
.B(n_2516),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3227),
.B(n_3225),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_SL g3457 ( 
.A(n_3291),
.B(n_2516),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_SL g3458 ( 
.A(n_3310),
.B(n_2516),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_SL g3459 ( 
.A(n_3310),
.B(n_3279),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3075),
.B(n_3068),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_SL g3461 ( 
.A(n_3310),
.B(n_2518),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_SL g3462 ( 
.A(n_3102),
.B(n_2518),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_SL g3463 ( 
.A(n_3289),
.B(n_2518),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_SL g3464 ( 
.A(n_3301),
.B(n_2518),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_3191),
.B(n_2561),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_SL g3466 ( 
.A(n_3126),
.B(n_2561),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3086),
.B(n_3050),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_SL g3468 ( 
.A(n_3126),
.B(n_2561),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_SL g3469 ( 
.A(n_3244),
.B(n_2561),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_SL g3470 ( 
.A(n_3244),
.B(n_2571),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_3080),
.B(n_2571),
.Y(n_3471)
);

NAND2xp33_ASAP7_75t_SL g3472 ( 
.A(n_3139),
.B(n_3083),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3087),
.B(n_3059),
.Y(n_3473)
);

NAND2xp33_ASAP7_75t_SL g3474 ( 
.A(n_3083),
.B(n_2571),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_3144),
.B(n_2571),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_SL g3476 ( 
.A(n_3209),
.B(n_2600),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3090),
.B(n_3043),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_SL g3478 ( 
.A(n_3209),
.B(n_3265),
.Y(n_3478)
);

NAND2xp33_ASAP7_75t_SL g3479 ( 
.A(n_3101),
.B(n_2600),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_SL g3480 ( 
.A(n_3265),
.B(n_2600),
.Y(n_3480)
);

AND2x2_ASAP7_75t_L g3481 ( 
.A(n_3295),
.B(n_887),
.Y(n_3481)
);

NAND2xp33_ASAP7_75t_SL g3482 ( 
.A(n_3101),
.B(n_2600),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_SL g3483 ( 
.A(n_3299),
.B(n_2606),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_SL g3484 ( 
.A(n_3299),
.B(n_2606),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_SL g3485 ( 
.A(n_3207),
.B(n_3268),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_SL g3486 ( 
.A(n_3293),
.B(n_3150),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_SL g3487 ( 
.A(n_3293),
.B(n_2606),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_SL g3488 ( 
.A(n_3150),
.B(n_3205),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_SL g3489 ( 
.A(n_3273),
.B(n_2606),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_SL g3490 ( 
.A(n_3176),
.B(n_2609),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_SL g3491 ( 
.A(n_3201),
.B(n_2609),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3297),
.B(n_3098),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_SL g3493 ( 
.A(n_3306),
.B(n_3288),
.Y(n_3493)
);

NAND2xp33_ASAP7_75t_SL g3494 ( 
.A(n_3092),
.B(n_2609),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_SL g3495 ( 
.A(n_3288),
.B(n_2609),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3109),
.B(n_3039),
.Y(n_3496)
);

NAND2xp33_ASAP7_75t_SL g3497 ( 
.A(n_3215),
.B(n_3196),
.Y(n_3497)
);

AND2x4_ASAP7_75t_L g3498 ( 
.A(n_3099),
.B(n_3224),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_SL g3499 ( 
.A(n_3294),
.B(n_2616),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_SL g3500 ( 
.A(n_3284),
.B(n_2616),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_SL g3501 ( 
.A(n_3287),
.B(n_2616),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_SL g3502 ( 
.A(n_3267),
.B(n_3224),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_SL g3503 ( 
.A(n_3267),
.B(n_2616),
.Y(n_3503)
);

NAND2xp33_ASAP7_75t_SL g3504 ( 
.A(n_3199),
.B(n_2664),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3117),
.B(n_3118),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_3200),
.B(n_2664),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3239),
.B(n_2664),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_SL g3508 ( 
.A(n_3128),
.B(n_2664),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_SL g3509 ( 
.A(n_3094),
.B(n_3032),
.Y(n_3509)
);

NAND2xp33_ASAP7_75t_SL g3510 ( 
.A(n_3199),
.B(n_2539),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3137),
.B(n_3041),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3152),
.B(n_3154),
.Y(n_3512)
);

NAND2xp33_ASAP7_75t_SL g3513 ( 
.A(n_3230),
.B(n_3241),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_SL g3514 ( 
.A(n_3241),
.B(n_3045),
.Y(n_3514)
);

NAND2xp33_ASAP7_75t_SL g3515 ( 
.A(n_3230),
.B(n_2577),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_3157),
.B(n_3005),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_SL g3517 ( 
.A(n_3161),
.B(n_3045),
.Y(n_3517)
);

NAND2xp33_ASAP7_75t_SL g3518 ( 
.A(n_3198),
.B(n_2584),
.Y(n_3518)
);

AND3x1_ASAP7_75t_L g3519 ( 
.A(n_3124),
.B(n_925),
.C(n_911),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_3247),
.B(n_3057),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_SL g3521 ( 
.A(n_3247),
.B(n_3057),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3158),
.B(n_2711),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_SL g3523 ( 
.A(n_3257),
.B(n_2805),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_SL g3524 ( 
.A(n_3106),
.B(n_2942),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_SL g3525 ( 
.A(n_3134),
.B(n_3254),
.Y(n_3525)
);

OAI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_3323),
.A2(n_3228),
.B1(n_3155),
.B2(n_3082),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_3505),
.Y(n_3527)
);

OR2x6_ASAP7_75t_L g3528 ( 
.A(n_3380),
.B(n_3129),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3512),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3332),
.B(n_3168),
.Y(n_3530)
);

AND2x2_ASAP7_75t_L g3531 ( 
.A(n_3334),
.B(n_3170),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3491),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3473),
.Y(n_3533)
);

NAND2xp33_ASAP7_75t_L g3534 ( 
.A(n_3313),
.B(n_3107),
.Y(n_3534)
);

OR2x2_ASAP7_75t_L g3535 ( 
.A(n_3364),
.B(n_3171),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3367),
.B(n_3173),
.Y(n_3536)
);

A2O1A1Ixp33_ASAP7_75t_L g3537 ( 
.A1(n_3317),
.A2(n_3141),
.B(n_2856),
.C(n_3292),
.Y(n_3537)
);

BUFx6f_ASAP7_75t_L g3538 ( 
.A(n_3354),
.Y(n_3538)
);

BUFx8_ASAP7_75t_SL g3539 ( 
.A(n_3456),
.Y(n_3539)
);

INVx2_ASAP7_75t_SL g3540 ( 
.A(n_3492),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3453),
.Y(n_3541)
);

O2A1O1Ixp5_ASAP7_75t_L g3542 ( 
.A1(n_3313),
.A2(n_3190),
.B(n_3184),
.C(n_3251),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3344),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3477),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3371),
.Y(n_3545)
);

OAI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_3405),
.A2(n_3256),
.B1(n_3263),
.B2(n_3260),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3525),
.A2(n_3315),
.B(n_3466),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3511),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3374),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_3460),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3467),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3338),
.B(n_3186),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3430),
.Y(n_3553)
);

INVx3_ASAP7_75t_L g3554 ( 
.A(n_3424),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_3522),
.Y(n_3555)
);

NAND3xp33_ASAP7_75t_L g3556 ( 
.A(n_3335),
.B(n_3274),
.C(n_968),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3363),
.B(n_3346),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3336),
.B(n_3187),
.Y(n_3558)
);

BUFx3_ASAP7_75t_L g3559 ( 
.A(n_3409),
.Y(n_3559)
);

AOI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_3525),
.A2(n_3286),
.B(n_2811),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3410),
.B(n_3194),
.Y(n_3561)
);

O2A1O1Ixp5_ASAP7_75t_SL g3562 ( 
.A1(n_3318),
.A2(n_3208),
.B(n_3214),
.C(n_3195),
.Y(n_3562)
);

AND2x4_ASAP7_75t_L g3563 ( 
.A(n_3498),
.B(n_3220),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3468),
.Y(n_3564)
);

HB1xp67_ASAP7_75t_L g3565 ( 
.A(n_3423),
.Y(n_3565)
);

INVx3_ASAP7_75t_L g3566 ( 
.A(n_3424),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3427),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_SL g3568 ( 
.A(n_3352),
.B(n_3130),
.Y(n_3568)
);

BUFx6f_ASAP7_75t_L g3569 ( 
.A(n_3354),
.Y(n_3569)
);

AOI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_3315),
.A2(n_3487),
.B(n_3322),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3496),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3402),
.Y(n_3572)
);

BUFx2_ASAP7_75t_L g3573 ( 
.A(n_3349),
.Y(n_3573)
);

AOI22xp5_ASAP7_75t_L g3574 ( 
.A1(n_3416),
.A2(n_3233),
.B1(n_3107),
.B2(n_2777),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_3428),
.Y(n_3575)
);

A2O1A1Ixp33_ASAP7_75t_L g3576 ( 
.A1(n_3316),
.A2(n_3221),
.B(n_3252),
.C(n_3226),
.Y(n_3576)
);

A2O1A1Ixp33_ASAP7_75t_L g3577 ( 
.A1(n_3485),
.A2(n_3270),
.B(n_3271),
.C(n_3261),
.Y(n_3577)
);

OAI21xp33_ASAP7_75t_L g3578 ( 
.A1(n_3524),
.A2(n_925),
.B(n_911),
.Y(n_3578)
);

OR2x2_ASAP7_75t_L g3579 ( 
.A(n_3350),
.B(n_3253),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3443),
.Y(n_3580)
);

CKINVDCx20_ASAP7_75t_R g3581 ( 
.A(n_3378),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3360),
.B(n_3280),
.Y(n_3582)
);

NOR2xp33_ASAP7_75t_L g3583 ( 
.A(n_3406),
.B(n_723),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3387),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3390),
.B(n_3281),
.Y(n_3585)
);

BUFx3_ASAP7_75t_L g3586 ( 
.A(n_3354),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3446),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3361),
.B(n_3283),
.Y(n_3588)
);

AND2x4_ASAP7_75t_L g3589 ( 
.A(n_3498),
.B(n_3285),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3362),
.B(n_3091),
.Y(n_3590)
);

INVx3_ASAP7_75t_L g3591 ( 
.A(n_3424),
.Y(n_3591)
);

INVx2_ASAP7_75t_L g3592 ( 
.A(n_3516),
.Y(n_3592)
);

INVx3_ASAP7_75t_L g3593 ( 
.A(n_3498),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3413),
.Y(n_3594)
);

AND2x4_ASAP7_75t_L g3595 ( 
.A(n_3436),
.B(n_3233),
.Y(n_3595)
);

AND2x4_ASAP7_75t_L g3596 ( 
.A(n_3436),
.B(n_3386),
.Y(n_3596)
);

NOR2xp33_ASAP7_75t_SL g3597 ( 
.A(n_3386),
.B(n_3211),
.Y(n_3597)
);

AND2x4_ASAP7_75t_L g3598 ( 
.A(n_3436),
.B(n_3258),
.Y(n_3598)
);

BUFx6f_ASAP7_75t_L g3599 ( 
.A(n_3386),
.Y(n_3599)
);

AOI21xp5_ASAP7_75t_L g3600 ( 
.A1(n_3426),
.A2(n_3286),
.B(n_2811),
.Y(n_3600)
);

BUFx6f_ASAP7_75t_L g3601 ( 
.A(n_3403),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3417),
.Y(n_3602)
);

OAI22xp33_ASAP7_75t_L g3603 ( 
.A1(n_3329),
.A2(n_2777),
.B1(n_3282),
.B2(n_959),
.Y(n_3603)
);

OAI22xp5_ASAP7_75t_L g3604 ( 
.A1(n_3519),
.A2(n_3489),
.B1(n_3330),
.B2(n_3340),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3365),
.B(n_3095),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3369),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3366),
.B(n_3321),
.Y(n_3607)
);

A2O1A1Ixp33_ASAP7_75t_SL g3608 ( 
.A1(n_3481),
.A2(n_926),
.B(n_944),
.C(n_937),
.Y(n_3608)
);

O2A1O1Ixp33_ASAP7_75t_L g3609 ( 
.A1(n_3392),
.A2(n_926),
.B(n_944),
.C(n_937),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3372),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3421),
.Y(n_3611)
);

BUFx2_ASAP7_75t_L g3612 ( 
.A(n_3345),
.Y(n_3612)
);

HB1xp67_ASAP7_75t_L g3613 ( 
.A(n_3486),
.Y(n_3613)
);

HB1xp67_ASAP7_75t_L g3614 ( 
.A(n_3422),
.Y(n_3614)
);

AOI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3434),
.A2(n_2948),
.B(n_2920),
.Y(n_3615)
);

INVx1_ASAP7_75t_SL g3616 ( 
.A(n_3327),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3373),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3431),
.Y(n_3618)
);

AOI21xp5_ASAP7_75t_L g3619 ( 
.A1(n_3435),
.A2(n_2495),
.B(n_2442),
.Y(n_3619)
);

BUFx2_ASAP7_75t_L g3620 ( 
.A(n_3353),
.Y(n_3620)
);

AOI222xp33_ASAP7_75t_L g3621 ( 
.A1(n_3328),
.A2(n_959),
.B1(n_949),
.B2(n_966),
.C1(n_954),
.C2(n_947),
.Y(n_3621)
);

OAI22xp33_ASAP7_75t_L g3622 ( 
.A1(n_3442),
.A2(n_980),
.B1(n_949),
.B2(n_954),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3377),
.B(n_3096),
.Y(n_3623)
);

INVx4_ASAP7_75t_L g3624 ( 
.A(n_3403),
.Y(n_3624)
);

BUFx6f_ASAP7_75t_L g3625 ( 
.A(n_3403),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_SL g3626 ( 
.A(n_3497),
.B(n_3206),
.Y(n_3626)
);

OR2x6_ASAP7_75t_L g3627 ( 
.A(n_3343),
.B(n_3312),
.Y(n_3627)
);

BUFx3_ASAP7_75t_L g3628 ( 
.A(n_3407),
.Y(n_3628)
);

BUFx6f_ASAP7_75t_L g3629 ( 
.A(n_3407),
.Y(n_3629)
);

HB1xp67_ASAP7_75t_L g3630 ( 
.A(n_3432),
.Y(n_3630)
);

BUFx3_ASAP7_75t_L g3631 ( 
.A(n_3407),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_3376),
.Y(n_3632)
);

INVx4_ASAP7_75t_L g3633 ( 
.A(n_3415),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3433),
.Y(n_3634)
);

NOR2x1_ASAP7_75t_L g3635 ( 
.A(n_3393),
.B(n_3420),
.Y(n_3635)
);

AOI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_3418),
.A2(n_3107),
.B1(n_2691),
.B2(n_3248),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3339),
.Y(n_3637)
);

OR2x6_ASAP7_75t_L g3638 ( 
.A(n_3343),
.B(n_3165),
.Y(n_3638)
);

CKINVDCx5p33_ASAP7_75t_R g3639 ( 
.A(n_3375),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_3494),
.B(n_3181),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3517),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3379),
.B(n_3097),
.Y(n_3642)
);

BUFx3_ASAP7_75t_L g3643 ( 
.A(n_3415),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3385),
.B(n_3116),
.Y(n_3644)
);

CKINVDCx5p33_ASAP7_75t_R g3645 ( 
.A(n_3415),
.Y(n_3645)
);

AOI22xp5_ASAP7_75t_L g3646 ( 
.A1(n_3414),
.A2(n_3107),
.B1(n_730),
.B2(n_733),
.Y(n_3646)
);

CKINVDCx5p33_ASAP7_75t_R g3647 ( 
.A(n_3472),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_3459),
.Y(n_3648)
);

INVx3_ASAP7_75t_L g3649 ( 
.A(n_3343),
.Y(n_3649)
);

CKINVDCx20_ASAP7_75t_R g3650 ( 
.A(n_3513),
.Y(n_3650)
);

OAI22xp5_ASAP7_75t_L g3651 ( 
.A1(n_3324),
.A2(n_2993),
.B1(n_2736),
.B2(n_2672),
.Y(n_3651)
);

O2A1O1Ixp33_ASAP7_75t_L g3652 ( 
.A1(n_3394),
.A2(n_947),
.B(n_968),
.C(n_966),
.Y(n_3652)
);

OAI21xp5_ASAP7_75t_L g3653 ( 
.A1(n_3508),
.A2(n_2866),
.B(n_2938),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3368),
.Y(n_3654)
);

INVx2_ASAP7_75t_SL g3655 ( 
.A(n_3502),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3356),
.Y(n_3656)
);

A2O1A1Ixp33_ASAP7_75t_L g3657 ( 
.A1(n_3384),
.A2(n_3333),
.B(n_3331),
.C(n_3325),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3514),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3404),
.B(n_980),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3408),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_3444),
.B(n_729),
.Y(n_3661)
);

BUFx6f_ASAP7_75t_L g3662 ( 
.A(n_3469),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3411),
.Y(n_3663)
);

O2A1O1Ixp33_ASAP7_75t_L g3664 ( 
.A1(n_3395),
.A2(n_1292),
.B(n_1293),
.C(n_1291),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3320),
.B(n_1047),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3429),
.Y(n_3666)
);

NAND2x2_ASAP7_75t_L g3667 ( 
.A(n_3314),
.B(n_1),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3388),
.B(n_3122),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3520),
.Y(n_3669)
);

AOI22xp5_ASAP7_75t_L g3670 ( 
.A1(n_3319),
.A2(n_737),
.B1(n_738),
.B2(n_735),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3389),
.B(n_3123),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3419),
.Y(n_3672)
);

NOR2xp33_ASAP7_75t_SL g3673 ( 
.A(n_3326),
.B(n_3211),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3488),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3521),
.Y(n_3675)
);

AOI21xp5_ASAP7_75t_L g3676 ( 
.A1(n_3391),
.A2(n_2495),
.B(n_2442),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3382),
.Y(n_3677)
);

BUFx2_ASAP7_75t_SL g3678 ( 
.A(n_3462),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3396),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3383),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3397),
.Y(n_3681)
);

OR2x6_ASAP7_75t_L g3682 ( 
.A(n_3493),
.B(n_3131),
.Y(n_3682)
);

OAI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_3348),
.A2(n_2089),
.B(n_2055),
.Y(n_3683)
);

OAI22xp5_ASAP7_75t_L g3684 ( 
.A1(n_3347),
.A2(n_2736),
.B1(n_2672),
.B2(n_2718),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3506),
.B(n_751),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3399),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3400),
.Y(n_3687)
);

A2O1A1Ixp33_ASAP7_75t_SL g3688 ( 
.A1(n_3425),
.A2(n_1295),
.B(n_1296),
.C(n_1294),
.Y(n_3688)
);

A2O1A1Ixp33_ASAP7_75t_L g3689 ( 
.A1(n_3342),
.A2(n_3243),
.B(n_1300),
.C(n_1301),
.Y(n_3689)
);

NOR2xp33_ASAP7_75t_L g3690 ( 
.A(n_3507),
.B(n_752),
.Y(n_3690)
);

INVx4_ASAP7_75t_L g3691 ( 
.A(n_3337),
.Y(n_3691)
);

INVx5_ASAP7_75t_L g3692 ( 
.A(n_3504),
.Y(n_3692)
);

OR2x6_ASAP7_75t_L g3693 ( 
.A(n_3358),
.B(n_3359),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3465),
.Y(n_3694)
);

INVx5_ASAP7_75t_L g3695 ( 
.A(n_3510),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3370),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3509),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3471),
.Y(n_3698)
);

BUFx8_ASAP7_75t_L g3699 ( 
.A(n_3412),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3351),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3357),
.B(n_3136),
.Y(n_3701)
);

BUFx6f_ASAP7_75t_L g3702 ( 
.A(n_3470),
.Y(n_3702)
);

INVx3_ASAP7_75t_L g3703 ( 
.A(n_3474),
.Y(n_3703)
);

O2A1O1Ixp5_ASAP7_75t_L g3704 ( 
.A1(n_3355),
.A2(n_3063),
.B(n_2623),
.C(n_2625),
.Y(n_3704)
);

NOR2xp33_ASAP7_75t_L g3705 ( 
.A(n_3500),
.B(n_753),
.Y(n_3705)
);

INVxp67_ASAP7_75t_L g3706 ( 
.A(n_3501),
.Y(n_3706)
);

OAI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_3475),
.A2(n_2718),
.B1(n_2291),
.B2(n_2545),
.Y(n_3707)
);

CKINVDCx20_ASAP7_75t_R g3708 ( 
.A(n_3381),
.Y(n_3708)
);

A2O1A1Ixp33_ASAP7_75t_L g3709 ( 
.A1(n_3401),
.A2(n_3341),
.B(n_3515),
.C(n_3499),
.Y(n_3709)
);

BUFx6f_ASAP7_75t_L g3710 ( 
.A(n_3483),
.Y(n_3710)
);

AND2x2_ASAP7_75t_SL g3711 ( 
.A(n_3479),
.B(n_843),
.Y(n_3711)
);

O2A1O1Ixp33_ASAP7_75t_SL g3712 ( 
.A1(n_3503),
.A2(n_843),
.B(n_879),
.C(n_1297),
.Y(n_3712)
);

INVxp67_ASAP7_75t_SL g3713 ( 
.A(n_3523),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3478),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_SL g3715 ( 
.A(n_3482),
.B(n_2584),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3490),
.Y(n_3716)
);

O2A1O1Ixp33_ASAP7_75t_L g3717 ( 
.A1(n_3463),
.A2(n_3464),
.B(n_1304),
.C(n_1308),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3495),
.B(n_3140),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_3398),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_SL g3720 ( 
.A(n_3518),
.B(n_2623),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3476),
.Y(n_3721)
);

O2A1O1Ixp33_ASAP7_75t_L g3722 ( 
.A1(n_3447),
.A2(n_1310),
.B(n_1311),
.C(n_1302),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3480),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3484),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3448),
.A2(n_2644),
.B(n_2636),
.Y(n_3725)
);

INVx3_ASAP7_75t_L g3726 ( 
.A(n_3437),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3449),
.Y(n_3727)
);

AOI22xp5_ASAP7_75t_L g3728 ( 
.A1(n_3438),
.A2(n_758),
.B1(n_762),
.B2(n_757),
.Y(n_3728)
);

NOR2xp33_ASAP7_75t_L g3729 ( 
.A(n_3450),
.B(n_763),
.Y(n_3729)
);

O2A1O1Ixp33_ASAP7_75t_L g3730 ( 
.A1(n_3461),
.A2(n_1314),
.B(n_1318),
.C(n_1313),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3451),
.Y(n_3731)
);

INVx3_ASAP7_75t_L g3732 ( 
.A(n_3439),
.Y(n_3732)
);

AOI21x1_ASAP7_75t_L g3733 ( 
.A1(n_3452),
.A2(n_1053),
.B(n_1049),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_SL g3734 ( 
.A(n_3440),
.B(n_2625),
.Y(n_3734)
);

INVx2_ASAP7_75t_L g3735 ( 
.A(n_3454),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3455),
.Y(n_3736)
);

OAI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_3441),
.A2(n_2291),
.B1(n_2545),
.B2(n_2542),
.Y(n_3737)
);

CKINVDCx20_ASAP7_75t_R g3738 ( 
.A(n_3458),
.Y(n_3738)
);

AND2x4_ASAP7_75t_L g3739 ( 
.A(n_3445),
.B(n_3149),
.Y(n_3739)
);

INVx1_ASAP7_75t_SL g3740 ( 
.A(n_3457),
.Y(n_3740)
);

INVx3_ASAP7_75t_SL g3741 ( 
.A(n_3334),
.Y(n_3741)
);

INVx4_ASAP7_75t_L g3742 ( 
.A(n_3424),
.Y(n_3742)
);

AOI21xp5_ASAP7_75t_L g3743 ( 
.A1(n_3313),
.A2(n_2645),
.B(n_2644),
.Y(n_3743)
);

BUFx10_ASAP7_75t_L g3744 ( 
.A(n_3354),
.Y(n_3744)
);

INVxp67_ASAP7_75t_L g3745 ( 
.A(n_3456),
.Y(n_3745)
);

HB1xp67_ASAP7_75t_L g3746 ( 
.A(n_3364),
.Y(n_3746)
);

OAI21x1_ASAP7_75t_L g3747 ( 
.A1(n_3615),
.A2(n_2602),
.B(n_2592),
.Y(n_3747)
);

OAI21xp5_ASAP7_75t_SL g3748 ( 
.A1(n_3622),
.A2(n_843),
.B(n_1319),
.Y(n_3748)
);

AOI21xp5_ASAP7_75t_L g3749 ( 
.A1(n_3600),
.A2(n_2658),
.B(n_2645),
.Y(n_3749)
);

OA21x2_ASAP7_75t_L g3750 ( 
.A1(n_3547),
.A2(n_1059),
.B(n_1057),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3565),
.B(n_1062),
.Y(n_3751)
);

BUFx2_ASAP7_75t_L g3752 ( 
.A(n_3573),
.Y(n_3752)
);

AOI22xp5_ASAP7_75t_L g3753 ( 
.A1(n_3546),
.A2(n_3603),
.B1(n_3604),
.B2(n_3534),
.Y(n_3753)
);

AOI21xp5_ASAP7_75t_L g3754 ( 
.A1(n_3560),
.A2(n_3657),
.B(n_3570),
.Y(n_3754)
);

OAI21x1_ASAP7_75t_L g3755 ( 
.A1(n_3562),
.A2(n_2602),
.B(n_2592),
.Y(n_3755)
);

CKINVDCx5p33_ASAP7_75t_R g3756 ( 
.A(n_3539),
.Y(n_3756)
);

HB1xp67_ASAP7_75t_L g3757 ( 
.A(n_3613),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3543),
.Y(n_3758)
);

HB1xp67_ASAP7_75t_L g3759 ( 
.A(n_3553),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_3695),
.A2(n_2682),
.B(n_2658),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3557),
.B(n_1064),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3741),
.B(n_1322),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3527),
.Y(n_3763)
);

AO22x2_ASAP7_75t_L g3764 ( 
.A1(n_3545),
.A2(n_3164),
.B1(n_3203),
.B2(n_3163),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3529),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3548),
.Y(n_3766)
);

BUFx3_ASAP7_75t_L g3767 ( 
.A(n_3559),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3533),
.Y(n_3768)
);

OAI22xp33_ASAP7_75t_L g3769 ( 
.A1(n_3574),
.A2(n_3667),
.B1(n_3636),
.B2(n_3646),
.Y(n_3769)
);

NAND3xp33_ASAP7_75t_L g3770 ( 
.A(n_3641),
.B(n_1067),
.C(n_1065),
.Y(n_3770)
);

OAI21x1_ASAP7_75t_L g3771 ( 
.A1(n_3653),
.A2(n_2612),
.B(n_2608),
.Y(n_3771)
);

OAI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3661),
.A2(n_3578),
.B(n_3537),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3544),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3745),
.B(n_1071),
.Y(n_3774)
);

AOI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_3695),
.A2(n_2688),
.B(n_2682),
.Y(n_3775)
);

O2A1O1Ixp5_ASAP7_75t_SL g3776 ( 
.A1(n_3594),
.A2(n_1074),
.B(n_1078),
.C(n_1073),
.Y(n_3776)
);

OAI21x1_ASAP7_75t_L g3777 ( 
.A1(n_3619),
.A2(n_2612),
.B(n_2608),
.Y(n_3777)
);

OAI21x1_ASAP7_75t_L g3778 ( 
.A1(n_3542),
.A2(n_3733),
.B(n_3703),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3746),
.B(n_1079),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3540),
.B(n_1323),
.Y(n_3780)
);

OAI21x1_ASAP7_75t_L g3781 ( 
.A1(n_3703),
.A2(n_2688),
.B(n_2620),
.Y(n_3781)
);

NOR2xp67_ASAP7_75t_L g3782 ( 
.A(n_3695),
.B(n_1080),
.Y(n_3782)
);

INVx2_ASAP7_75t_SL g3783 ( 
.A(n_3645),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3592),
.Y(n_3784)
);

AOI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_3711),
.A2(n_2590),
.B(n_2586),
.Y(n_3785)
);

OAI21x1_ASAP7_75t_L g3786 ( 
.A1(n_3651),
.A2(n_2116),
.B(n_2101),
.Y(n_3786)
);

OAI21x1_ASAP7_75t_L g3787 ( 
.A1(n_3743),
.A2(n_2116),
.B(n_2101),
.Y(n_3787)
);

INVx1_ASAP7_75t_SL g3788 ( 
.A(n_3582),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3550),
.Y(n_3789)
);

OAI21xp5_ASAP7_75t_L g3790 ( 
.A1(n_3670),
.A2(n_879),
.B(n_1324),
.Y(n_3790)
);

CKINVDCx6p67_ASAP7_75t_R g3791 ( 
.A(n_3528),
.Y(n_3791)
);

AOI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3692),
.A2(n_2590),
.B(n_2586),
.Y(n_3792)
);

CKINVDCx8_ASAP7_75t_R g3793 ( 
.A(n_3639),
.Y(n_3793)
);

AOI21xp5_ASAP7_75t_L g3794 ( 
.A1(n_3692),
.A2(n_2542),
.B(n_2591),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3530),
.B(n_1105),
.Y(n_3795)
);

AOI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_3692),
.A2(n_2596),
.B(n_2591),
.Y(n_3796)
);

OAI21x1_ASAP7_75t_L g3797 ( 
.A1(n_3635),
.A2(n_2119),
.B(n_2375),
.Y(n_3797)
);

AOI221xp5_ASAP7_75t_SL g3798 ( 
.A1(n_3609),
.A2(n_1329),
.B1(n_1332),
.B2(n_1328),
.C(n_1325),
.Y(n_3798)
);

OR2x2_ASAP7_75t_L g3799 ( 
.A(n_3579),
.B(n_1111),
.Y(n_3799)
);

AOI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_3626),
.A2(n_2598),
.B(n_2596),
.Y(n_3800)
);

OAI21x1_ASAP7_75t_L g3801 ( 
.A1(n_3707),
.A2(n_2119),
.B(n_2375),
.Y(n_3801)
);

OAI22xp5_ASAP7_75t_L g3802 ( 
.A1(n_3581),
.A2(n_2647),
.B1(n_2668),
.B2(n_2598),
.Y(n_3802)
);

OAI21x1_ASAP7_75t_L g3803 ( 
.A1(n_3594),
.A2(n_2381),
.B(n_2378),
.Y(n_3803)
);

CKINVDCx5p33_ASAP7_75t_R g3804 ( 
.A(n_3647),
.Y(n_3804)
);

AO31x2_ASAP7_75t_L g3805 ( 
.A1(n_3687),
.A2(n_3641),
.A3(n_3719),
.B(n_3602),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3532),
.Y(n_3806)
);

A2O1A1Ixp33_ASAP7_75t_L g3807 ( 
.A1(n_3689),
.A2(n_1113),
.B(n_1114),
.C(n_1112),
.Y(n_3807)
);

NAND3x1_ASAP7_75t_L g3808 ( 
.A(n_3531),
.B(n_3585),
.C(n_3607),
.Y(n_3808)
);

OAI21x1_ASAP7_75t_L g3809 ( 
.A1(n_3602),
.A2(n_2381),
.B(n_2378),
.Y(n_3809)
);

OR2x2_ASAP7_75t_L g3810 ( 
.A(n_3572),
.B(n_1115),
.Y(n_3810)
);

OAI21xp5_ASAP7_75t_SL g3811 ( 
.A1(n_3621),
.A2(n_1339),
.B(n_1337),
.Y(n_3811)
);

OR2x2_ASAP7_75t_L g3812 ( 
.A(n_3584),
.B(n_1116),
.Y(n_3812)
);

OAI21x1_ASAP7_75t_L g3813 ( 
.A1(n_3532),
.A2(n_2396),
.B(n_2388),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3551),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3567),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3596),
.B(n_1340),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3709),
.A2(n_2668),
.B(n_2647),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3713),
.A2(n_2663),
.B(n_2639),
.Y(n_3818)
);

INVx1_ASAP7_75t_SL g3819 ( 
.A(n_3708),
.Y(n_3819)
);

OAI22x1_ASAP7_75t_L g3820 ( 
.A1(n_3571),
.A2(n_1118),
.B1(n_1117),
.B2(n_769),
.Y(n_3820)
);

OAI21x1_ASAP7_75t_L g3821 ( 
.A1(n_3676),
.A2(n_2396),
.B(n_2388),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3720),
.A2(n_2663),
.B(n_2639),
.Y(n_3822)
);

O2A1O1Ixp33_ASAP7_75t_L g3823 ( 
.A1(n_3608),
.A2(n_1343),
.B(n_1344),
.C(n_1342),
.Y(n_3823)
);

INVx1_ASAP7_75t_SL g3824 ( 
.A(n_3616),
.Y(n_3824)
);

AOI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_3640),
.A2(n_2692),
.B(n_2669),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3660),
.Y(n_3826)
);

AOI21xp5_ASAP7_75t_L g3827 ( 
.A1(n_3612),
.A2(n_2692),
.B(n_2669),
.Y(n_3827)
);

INVx3_ASAP7_75t_L g3828 ( 
.A(n_3742),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3568),
.A2(n_2055),
.B(n_2051),
.Y(n_3829)
);

O2A1O1Ixp33_ASAP7_75t_SL g3830 ( 
.A1(n_3526),
.A2(n_1358),
.B(n_1360),
.C(n_1349),
.Y(n_3830)
);

OAI21xp5_ASAP7_75t_SL g3831 ( 
.A1(n_3652),
.A2(n_1361),
.B(n_2),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3681),
.B(n_2),
.Y(n_3832)
);

OAI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3576),
.A2(n_771),
.B(n_764),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_3593),
.B(n_3217),
.Y(n_3834)
);

OAI21xp33_ASAP7_75t_L g3835 ( 
.A1(n_3564),
.A2(n_805),
.B(n_775),
.Y(n_3835)
);

AOI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3688),
.A2(n_2110),
.B(n_2051),
.Y(n_3836)
);

AO21x2_ASAP7_75t_L g3837 ( 
.A1(n_3701),
.A2(n_3236),
.B(n_3218),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3555),
.Y(n_3838)
);

AOI211xp5_ASAP7_75t_L g3839 ( 
.A1(n_3583),
.A2(n_774),
.B(n_777),
.C(n_773),
.Y(n_3839)
);

AND2x4_ASAP7_75t_L g3840 ( 
.A(n_3593),
.B(n_3238),
.Y(n_3840)
);

NAND2x1p5_ASAP7_75t_L g3841 ( 
.A(n_3691),
.B(n_3262),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3620),
.B(n_3276),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3541),
.Y(n_3843)
);

OAI22x1_ASAP7_75t_L g3844 ( 
.A1(n_3587),
.A2(n_787),
.B1(n_788),
.B2(n_780),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_3715),
.A2(n_2110),
.B(n_2291),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3561),
.B(n_4),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3549),
.B(n_4),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3596),
.B(n_1132),
.Y(n_3848)
);

AO31x2_ASAP7_75t_L g3849 ( 
.A1(n_3686),
.A2(n_3304),
.A3(n_2735),
.B(n_2741),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3535),
.Y(n_3850)
);

AOI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3673),
.A2(n_2321),
.B(n_2319),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3679),
.B(n_3552),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3624),
.B(n_5),
.Y(n_3853)
);

BUFx3_ASAP7_75t_L g3854 ( 
.A(n_3699),
.Y(n_3854)
);

OAI22xp5_ASAP7_75t_L g3855 ( 
.A1(n_3556),
.A2(n_793),
.B1(n_794),
.B2(n_791),
.Y(n_3855)
);

BUFx2_ASAP7_75t_SL g3856 ( 
.A(n_3650),
.Y(n_3856)
);

OAI21x1_ASAP7_75t_L g3857 ( 
.A1(n_3725),
.A2(n_2321),
.B(n_2319),
.Y(n_3857)
);

AOI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_3691),
.A2(n_2389),
.B(n_2376),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3554),
.B(n_1132),
.Y(n_3859)
);

OAI221xp5_ASAP7_75t_L g3860 ( 
.A1(n_3577),
.A2(n_802),
.B1(n_804),
.B2(n_800),
.C(n_799),
.Y(n_3860)
);

AOI21xp5_ASAP7_75t_L g3861 ( 
.A1(n_3597),
.A2(n_2389),
.B(n_2376),
.Y(n_3861)
);

AOI21xp5_ASAP7_75t_L g3862 ( 
.A1(n_3712),
.A2(n_2391),
.B(n_2385),
.Y(n_3862)
);

NOR2x1_ASAP7_75t_R g3863 ( 
.A(n_3742),
.B(n_806),
.Y(n_3863)
);

OAI21xp5_ASAP7_75t_L g3864 ( 
.A1(n_3729),
.A2(n_808),
.B(n_807),
.Y(n_3864)
);

NOR2xp33_ASAP7_75t_SL g3865 ( 
.A(n_3699),
.B(n_2087),
.Y(n_3865)
);

AOI21xp5_ASAP7_75t_L g3866 ( 
.A1(n_3734),
.A2(n_2391),
.B(n_2398),
.Y(n_3866)
);

A2O1A1Ixp33_ASAP7_75t_L g3867 ( 
.A1(n_3685),
.A2(n_812),
.B(n_815),
.C(n_814),
.Y(n_3867)
);

OAI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3690),
.A2(n_818),
.B(n_809),
.Y(n_3868)
);

AOI21xp5_ASAP7_75t_L g3869 ( 
.A1(n_3564),
.A2(n_2379),
.B(n_2377),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3660),
.Y(n_3870)
);

OAI22xp5_ASAP7_75t_L g3871 ( 
.A1(n_3738),
.A2(n_824),
.B1(n_831),
.B2(n_820),
.Y(n_3871)
);

AND2x4_ASAP7_75t_L g3872 ( 
.A(n_3554),
.B(n_1181),
.Y(n_3872)
);

BUFx6f_ASAP7_75t_L g3873 ( 
.A(n_3538),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_3588),
.Y(n_3874)
);

OAI21x1_ASAP7_75t_L g3875 ( 
.A1(n_3683),
.A2(n_2386),
.B(n_2380),
.Y(n_3875)
);

BUFx2_ASAP7_75t_L g3876 ( 
.A(n_3624),
.Y(n_3876)
);

OAI21x1_ASAP7_75t_L g3877 ( 
.A1(n_3697),
.A2(n_2397),
.B(n_2098),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3575),
.Y(n_3878)
);

NOR2x1_ASAP7_75t_SL g3879 ( 
.A(n_3693),
.B(n_3682),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3566),
.B(n_1181),
.Y(n_3880)
);

AOI21x1_ASAP7_75t_L g3881 ( 
.A1(n_3665),
.A2(n_1213),
.B(n_1193),
.Y(n_3881)
);

AOI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3663),
.A2(n_2104),
.B(n_2091),
.Y(n_3882)
);

NAND3xp33_ASAP7_75t_L g3883 ( 
.A(n_3674),
.B(n_1213),
.C(n_1193),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3536),
.B(n_6),
.Y(n_3884)
);

AO31x2_ASAP7_75t_L g3885 ( 
.A1(n_3663),
.A2(n_3672),
.A3(n_3666),
.B(n_3611),
.Y(n_3885)
);

OA21x2_ASAP7_75t_L g3886 ( 
.A1(n_3656),
.A2(n_3637),
.B(n_3618),
.Y(n_3886)
);

OAI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_3705),
.A2(n_837),
.B(n_834),
.Y(n_3887)
);

NOR2xp67_ASAP7_75t_L g3888 ( 
.A(n_3558),
.B(n_1219),
.Y(n_3888)
);

INVxp67_ASAP7_75t_L g3889 ( 
.A(n_3614),
.Y(n_3889)
);

AND2x4_ASAP7_75t_L g3890 ( 
.A(n_3566),
.B(n_1219),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3637),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3580),
.B(n_7),
.Y(n_3892)
);

O2A1O1Ixp33_ASAP7_75t_L g3893 ( 
.A1(n_3664),
.A2(n_1242),
.B(n_1257),
.C(n_1220),
.Y(n_3893)
);

A2O1A1Ixp33_ASAP7_75t_L g3894 ( 
.A1(n_3659),
.A2(n_840),
.B(n_846),
.C(n_838),
.Y(n_3894)
);

AOI22xp5_ASAP7_75t_L g3895 ( 
.A1(n_3563),
.A2(n_850),
.B1(n_851),
.B2(n_847),
.Y(n_3895)
);

INVx2_ASAP7_75t_SL g3896 ( 
.A(n_3538),
.Y(n_3896)
);

OAI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3706),
.A2(n_855),
.B(n_852),
.Y(n_3897)
);

BUFx2_ASAP7_75t_L g3898 ( 
.A(n_3633),
.Y(n_3898)
);

NAND3xp33_ASAP7_75t_L g3899 ( 
.A(n_3716),
.B(n_1242),
.C(n_1220),
.Y(n_3899)
);

NAND3xp33_ASAP7_75t_L g3900 ( 
.A(n_3700),
.B(n_1258),
.C(n_1257),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_SL g3901 ( 
.A(n_3710),
.B(n_1258),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3648),
.B(n_7),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3669),
.B(n_9),
.Y(n_3903)
);

NOR2xp67_ASAP7_75t_SL g3904 ( 
.A(n_3678),
.B(n_963),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_3675),
.B(n_9),
.Y(n_3905)
);

AOI21xp5_ASAP7_75t_L g3906 ( 
.A1(n_3656),
.A2(n_2107),
.B(n_2106),
.Y(n_3906)
);

CKINVDCx5p33_ASAP7_75t_R g3907 ( 
.A(n_3528),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_3737),
.A2(n_2185),
.B(n_2169),
.Y(n_3908)
);

OA21x2_ASAP7_75t_L g3909 ( 
.A1(n_3611),
.A2(n_1275),
.B(n_1260),
.Y(n_3909)
);

BUFx3_ASAP7_75t_L g3910 ( 
.A(n_3538),
.Y(n_3910)
);

A2O1A1Ixp33_ASAP7_75t_L g3911 ( 
.A1(n_3728),
.A2(n_861),
.B(n_862),
.C(n_860),
.Y(n_3911)
);

BUFx6f_ASAP7_75t_L g3912 ( 
.A(n_3569),
.Y(n_3912)
);

OAI21x1_ASAP7_75t_L g3913 ( 
.A1(n_3704),
.A2(n_2743),
.B(n_2721),
.Y(n_3913)
);

OAI21x1_ASAP7_75t_L g3914 ( 
.A1(n_3727),
.A2(n_2753),
.B(n_2746),
.Y(n_3914)
);

INVx8_ASAP7_75t_L g3915 ( 
.A(n_3682),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3618),
.Y(n_3916)
);

OAI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3727),
.A2(n_3736),
.B(n_3731),
.Y(n_3917)
);

OAI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3731),
.A2(n_3736),
.B(n_3634),
.Y(n_3918)
);

O2A1O1Ixp33_ASAP7_75t_SL g3919 ( 
.A1(n_3655),
.A2(n_14),
.B(n_11),
.C(n_12),
.Y(n_3919)
);

AO31x2_ASAP7_75t_L g3920 ( 
.A1(n_3634),
.A2(n_3606),
.A3(n_3721),
.B(n_3698),
.Y(n_3920)
);

AOI22xp33_ASAP7_75t_L g3921 ( 
.A1(n_3696),
.A2(n_2754),
.B1(n_2172),
.B2(n_2179),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3684),
.A2(n_2185),
.B(n_2169),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_3740),
.A2(n_2185),
.B(n_2169),
.Y(n_3923)
);

AO31x2_ASAP7_75t_L g3924 ( 
.A1(n_3677),
.A2(n_3714),
.A3(n_3617),
.B(n_3632),
.Y(n_3924)
);

AO31x2_ASAP7_75t_L g3925 ( 
.A1(n_3610),
.A2(n_1275),
.A3(n_1260),
.B(n_2174),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3590),
.Y(n_3926)
);

AOI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_3630),
.A2(n_2193),
.B(n_2185),
.Y(n_3927)
);

A2O1A1Ixp33_ASAP7_75t_L g3928 ( 
.A1(n_3717),
.A2(n_865),
.B(n_871),
.C(n_864),
.Y(n_3928)
);

AOI21x1_ASAP7_75t_L g3929 ( 
.A1(n_3723),
.A2(n_989),
.B(n_983),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3605),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_3693),
.A2(n_2205),
.B(n_2193),
.Y(n_3931)
);

A2O1A1Ixp33_ASAP7_75t_L g3932 ( 
.A1(n_3658),
.A2(n_872),
.B(n_877),
.C(n_869),
.Y(n_3932)
);

OAI21xp5_ASAP7_75t_L g3933 ( 
.A1(n_3680),
.A2(n_886),
.B(n_880),
.Y(n_3933)
);

INVx1_ASAP7_75t_SL g3934 ( 
.A(n_3586),
.Y(n_3934)
);

NAND2x1p5_ASAP7_75t_L g3935 ( 
.A(n_3633),
.B(n_2269),
.Y(n_3935)
);

AO31x2_ASAP7_75t_L g3936 ( 
.A1(n_3724),
.A2(n_2179),
.A3(n_2174),
.B(n_2181),
.Y(n_3936)
);

OAI21x1_ASAP7_75t_L g3937 ( 
.A1(n_3735),
.A2(n_3732),
.B(n_3726),
.Y(n_3937)
);

BUFx2_ASAP7_75t_L g3938 ( 
.A(n_3628),
.Y(n_3938)
);

A2O1A1Ixp33_ASAP7_75t_L g3939 ( 
.A1(n_3563),
.A2(n_890),
.B(n_891),
.C(n_889),
.Y(n_3939)
);

NOR2xp33_ASAP7_75t_L g3940 ( 
.A(n_3569),
.B(n_16),
.Y(n_3940)
);

INVx3_ASAP7_75t_L g3941 ( 
.A(n_3591),
.Y(n_3941)
);

NAND3x1_ASAP7_75t_L g3942 ( 
.A(n_3591),
.B(n_16),
.C(n_17),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3644),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3589),
.B(n_19),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3726),
.A2(n_2205),
.B(n_2193),
.Y(n_3945)
);

AOI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_3732),
.A2(n_2205),
.B(n_2193),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3668),
.Y(n_3947)
);

AO21x1_ASAP7_75t_L g3948 ( 
.A1(n_3589),
.A2(n_21),
.B(n_22),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_SL g3949 ( 
.A(n_3710),
.B(n_2205),
.Y(n_3949)
);

OAI21x1_ASAP7_75t_L g3950 ( 
.A1(n_3623),
.A2(n_2045),
.B(n_2126),
.Y(n_3950)
);

A2O1A1Ixp33_ASAP7_75t_L g3951 ( 
.A1(n_3654),
.A2(n_893),
.B(n_894),
.C(n_892),
.Y(n_3951)
);

CKINVDCx5p33_ASAP7_75t_R g3952 ( 
.A(n_3569),
.Y(n_3952)
);

BUFx12f_ASAP7_75t_L g3953 ( 
.A(n_3599),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3671),
.B(n_21),
.Y(n_3954)
);

OAI21x1_ASAP7_75t_L g3955 ( 
.A1(n_3642),
.A2(n_2045),
.B(n_2181),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3694),
.Y(n_3956)
);

AO31x2_ASAP7_75t_L g3957 ( 
.A1(n_3718),
.A2(n_2189),
.A3(n_2198),
.B(n_2188),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3649),
.Y(n_3958)
);

O2A1O1Ixp5_ASAP7_75t_SL g3959 ( 
.A1(n_3649),
.A2(n_2142),
.B(n_2300),
.C(n_2269),
.Y(n_3959)
);

INVx2_ASAP7_75t_L g3960 ( 
.A(n_3739),
.Y(n_3960)
);

AO31x2_ASAP7_75t_L g3961 ( 
.A1(n_3739),
.A2(n_2189),
.A3(n_2198),
.B(n_2188),
.Y(n_3961)
);

O2A1O1Ixp33_ASAP7_75t_L g3962 ( 
.A1(n_3722),
.A2(n_2223),
.B(n_2199),
.C(n_2300),
.Y(n_3962)
);

BUFx2_ASAP7_75t_L g3963 ( 
.A(n_3631),
.Y(n_3963)
);

OAI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_3730),
.A2(n_897),
.B(n_896),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3710),
.Y(n_3965)
);

INVx4_ASAP7_75t_L g3966 ( 
.A(n_3662),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3643),
.B(n_22),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3662),
.Y(n_3968)
);

AOI21x1_ASAP7_75t_L g3969 ( 
.A1(n_3598),
.A2(n_989),
.B(n_983),
.Y(n_3969)
);

HB1xp67_ASAP7_75t_L g3970 ( 
.A(n_3662),
.Y(n_3970)
);

INVx4_ASAP7_75t_L g3971 ( 
.A(n_3702),
.Y(n_3971)
);

BUFx12f_ASAP7_75t_L g3972 ( 
.A(n_3599),
.Y(n_3972)
);

OAI21x1_ASAP7_75t_L g3973 ( 
.A1(n_3778),
.A2(n_3927),
.B(n_3923),
.Y(n_3973)
);

A2O1A1Ixp33_ASAP7_75t_L g3974 ( 
.A1(n_3772),
.A2(n_3754),
.B(n_3753),
.C(n_3831),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3891),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3920),
.Y(n_3976)
);

NOR2xp33_ASAP7_75t_L g3977 ( 
.A(n_3793),
.B(n_3599),
.Y(n_3977)
);

CKINVDCx11_ASAP7_75t_R g3978 ( 
.A(n_3819),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3891),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3920),
.Y(n_3980)
);

BUFx10_ASAP7_75t_L g3981 ( 
.A(n_3756),
.Y(n_3981)
);

OAI21x1_ASAP7_75t_L g3982 ( 
.A1(n_3781),
.A2(n_3744),
.B(n_2223),
.Y(n_3982)
);

OAI21x1_ASAP7_75t_L g3983 ( 
.A1(n_3803),
.A2(n_3744),
.B(n_2199),
.Y(n_3983)
);

OAI21x1_ASAP7_75t_L g3984 ( 
.A1(n_3809),
.A2(n_3702),
.B(n_2045),
.Y(n_3984)
);

NOR2x1_ASAP7_75t_SL g3985 ( 
.A(n_3842),
.B(n_3601),
.Y(n_3985)
);

BUFx2_ASAP7_75t_L g3986 ( 
.A(n_3752),
.Y(n_3986)
);

NOR2xp33_ASAP7_75t_L g3987 ( 
.A(n_3824),
.B(n_3601),
.Y(n_3987)
);

OR2x6_ASAP7_75t_SL g3988 ( 
.A(n_3907),
.B(n_899),
.Y(n_3988)
);

OAI22xp33_ASAP7_75t_L g3989 ( 
.A1(n_3769),
.A2(n_3638),
.B1(n_3627),
.B2(n_3702),
.Y(n_3989)
);

AO31x2_ASAP7_75t_L g3990 ( 
.A1(n_3956),
.A2(n_1022),
.A3(n_1029),
.B(n_999),
.Y(n_3990)
);

OAI21x1_ASAP7_75t_L g3991 ( 
.A1(n_3937),
.A2(n_2303),
.B(n_3627),
.Y(n_3991)
);

OAI21x1_ASAP7_75t_L g3992 ( 
.A1(n_3931),
.A2(n_2303),
.B(n_2229),
.Y(n_3992)
);

OAI21x1_ASAP7_75t_SL g3993 ( 
.A1(n_3879),
.A2(n_23),
.B(n_24),
.Y(n_3993)
);

AO21x2_ASAP7_75t_L g3994 ( 
.A1(n_3888),
.A2(n_3598),
.B(n_3595),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3767),
.B(n_3788),
.Y(n_3995)
);

AOI21xp33_ASAP7_75t_L g3996 ( 
.A1(n_3820),
.A2(n_3638),
.B(n_3595),
.Y(n_3996)
);

OAI21x1_ASAP7_75t_L g3997 ( 
.A1(n_3929),
.A2(n_3625),
.B(n_3601),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_SL g3998 ( 
.A(n_3917),
.B(n_3625),
.Y(n_3998)
);

AND2x4_ASAP7_75t_L g3999 ( 
.A(n_3941),
.B(n_3625),
.Y(n_3999)
);

OAI22xp33_ASAP7_75t_L g4000 ( 
.A1(n_3915),
.A2(n_3629),
.B1(n_904),
.B2(n_905),
.Y(n_4000)
);

AO21x2_ASAP7_75t_L g4001 ( 
.A1(n_3918),
.A2(n_1022),
.B(n_999),
.Y(n_4001)
);

AOI21xp33_ASAP7_75t_SL g4002 ( 
.A1(n_3804),
.A2(n_23),
.B(n_26),
.Y(n_4002)
);

OAI21x1_ASAP7_75t_L g4003 ( 
.A1(n_3786),
.A2(n_3629),
.B(n_1034),
.Y(n_4003)
);

NOR2xp33_ASAP7_75t_L g4004 ( 
.A(n_3854),
.B(n_3629),
.Y(n_4004)
);

BUFx2_ASAP7_75t_L g4005 ( 
.A(n_3757),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3826),
.Y(n_4006)
);

AO31x2_ASAP7_75t_L g4007 ( 
.A1(n_3806),
.A2(n_1034),
.A3(n_1045),
.B(n_1029),
.Y(n_4007)
);

BUFx6f_ASAP7_75t_L g4008 ( 
.A(n_3873),
.Y(n_4008)
);

OA21x2_ASAP7_75t_L g4009 ( 
.A1(n_3806),
.A2(n_906),
.B(n_902),
.Y(n_4009)
);

OAI21x1_ASAP7_75t_L g4010 ( 
.A1(n_3945),
.A2(n_1050),
.B(n_1045),
.Y(n_4010)
);

OAI21x1_ASAP7_75t_L g4011 ( 
.A1(n_3946),
.A2(n_1084),
.B(n_1050),
.Y(n_4011)
);

BUFx6f_ASAP7_75t_L g4012 ( 
.A(n_3873),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3826),
.Y(n_4013)
);

INVx6_ASAP7_75t_SL g4014 ( 
.A(n_3834),
.Y(n_4014)
);

CKINVDCx11_ASAP7_75t_R g4015 ( 
.A(n_3791),
.Y(n_4015)
);

AOI21xp33_ASAP7_75t_L g4016 ( 
.A1(n_3916),
.A2(n_908),
.B(n_907),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_3920),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_3948),
.A2(n_2221),
.B1(n_2225),
.B2(n_2215),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3870),
.Y(n_4019)
);

OAI21x1_ASAP7_75t_L g4020 ( 
.A1(n_3813),
.A2(n_1091),
.B(n_1084),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3870),
.Y(n_4021)
);

OAI22xp5_ASAP7_75t_SL g4022 ( 
.A1(n_3856),
.A2(n_910),
.B1(n_912),
.B2(n_909),
.Y(n_4022)
);

OAI21x1_ASAP7_75t_L g4023 ( 
.A1(n_3869),
.A2(n_1095),
.B(n_1091),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3759),
.Y(n_4024)
);

OR2x2_ASAP7_75t_L g4025 ( 
.A(n_3850),
.B(n_3889),
.Y(n_4025)
);

OAI21x1_ASAP7_75t_L g4026 ( 
.A1(n_3950),
.A2(n_1095),
.B(n_27),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3766),
.Y(n_4027)
);

INVx8_ASAP7_75t_L g4028 ( 
.A(n_3915),
.Y(n_4028)
);

BUFx6f_ASAP7_75t_L g4029 ( 
.A(n_3873),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3885),
.Y(n_4030)
);

INVx2_ASAP7_75t_L g4031 ( 
.A(n_3885),
.Y(n_4031)
);

OAI21x1_ASAP7_75t_L g4032 ( 
.A1(n_3776),
.A2(n_27),
.B(n_28),
.Y(n_4032)
);

BUFx4f_ASAP7_75t_L g4033 ( 
.A(n_3841),
.Y(n_4033)
);

A2O1A1Ixp33_ASAP7_75t_SL g4034 ( 
.A1(n_3853),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_4034)
);

AO21x2_ASAP7_75t_L g4035 ( 
.A1(n_3751),
.A2(n_916),
.B(n_915),
.Y(n_4035)
);

NOR2xp33_ASAP7_75t_L g4036 ( 
.A(n_3762),
.B(n_29),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3885),
.Y(n_4037)
);

AOI22xp33_ASAP7_75t_L g4038 ( 
.A1(n_3960),
.A2(n_2221),
.B1(n_2225),
.B2(n_2215),
.Y(n_4038)
);

OAI21x1_ASAP7_75t_SL g4039 ( 
.A1(n_3852),
.A2(n_31),
.B(n_32),
.Y(n_4039)
);

OAI21x1_ASAP7_75t_L g4040 ( 
.A1(n_3747),
.A2(n_31),
.B(n_33),
.Y(n_4040)
);

NAND2xp33_ASAP7_75t_SL g4041 ( 
.A(n_3876),
.B(n_919),
.Y(n_4041)
);

OAI21xp5_ASAP7_75t_L g4042 ( 
.A1(n_3942),
.A2(n_924),
.B(n_920),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3947),
.Y(n_4043)
);

AOI21xp5_ASAP7_75t_L g4044 ( 
.A1(n_3792),
.A2(n_3749),
.B(n_3908),
.Y(n_4044)
);

NOR2xp67_ASAP7_75t_L g4045 ( 
.A(n_3774),
.B(n_34),
.Y(n_4045)
);

HB1xp67_ASAP7_75t_L g4046 ( 
.A(n_3805),
.Y(n_4046)
);

OAI21xp5_ASAP7_75t_L g4047 ( 
.A1(n_3833),
.A2(n_928),
.B(n_927),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3924),
.Y(n_4048)
);

O2A1O1Ixp33_ASAP7_75t_L g4049 ( 
.A1(n_3830),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_3924),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3947),
.Y(n_4051)
);

AO21x1_ASAP7_75t_L g4052 ( 
.A1(n_3846),
.A2(n_35),
.B(n_36),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3758),
.Y(n_4053)
);

OAI21x1_ASAP7_75t_L g4054 ( 
.A1(n_3797),
.A2(n_37),
.B(n_38),
.Y(n_4054)
);

OAI21x1_ASAP7_75t_L g4055 ( 
.A1(n_3881),
.A2(n_37),
.B(n_39),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3874),
.Y(n_4056)
);

AOI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3808),
.A2(n_934),
.B1(n_936),
.B2(n_932),
.Y(n_4057)
);

OAI22xp5_ASAP7_75t_L g4058 ( 
.A1(n_3860),
.A2(n_941),
.B1(n_943),
.B2(n_939),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_3924),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_3941),
.B(n_41),
.Y(n_4060)
);

NOR2xp33_ASAP7_75t_SL g4061 ( 
.A(n_3863),
.B(n_945),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_3805),
.Y(n_4062)
);

AOI21xp5_ASAP7_75t_L g4063 ( 
.A1(n_3760),
.A2(n_2221),
.B(n_2215),
.Y(n_4063)
);

OR2x2_ASAP7_75t_L g4064 ( 
.A(n_3843),
.B(n_42),
.Y(n_4064)
);

AND2x4_ASAP7_75t_L g4065 ( 
.A(n_3958),
.B(n_43),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3943),
.Y(n_4066)
);

OAI21x1_ASAP7_75t_L g4067 ( 
.A1(n_3882),
.A2(n_43),
.B(n_44),
.Y(n_4067)
);

NAND3xp33_ASAP7_75t_L g4068 ( 
.A(n_3832),
.B(n_951),
.C(n_950),
.Y(n_4068)
);

AND2x2_ASAP7_75t_L g4069 ( 
.A(n_3938),
.B(n_45),
.Y(n_4069)
);

OR2x6_ASAP7_75t_L g4070 ( 
.A(n_3953),
.B(n_3972),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_SL g4071 ( 
.A(n_3966),
.B(n_952),
.Y(n_4071)
);

OAI21x1_ASAP7_75t_L g4072 ( 
.A1(n_3955),
.A2(n_45),
.B(n_46),
.Y(n_4072)
);

OAI21x1_ASAP7_75t_L g4073 ( 
.A1(n_3877),
.A2(n_47),
.B(n_49),
.Y(n_4073)
);

OAI21x1_ASAP7_75t_L g4074 ( 
.A1(n_3787),
.A2(n_49),
.B(n_50),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3926),
.B(n_956),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3930),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3805),
.Y(n_4077)
);

AOI221xp5_ASAP7_75t_L g4078 ( 
.A1(n_3919),
.A2(n_967),
.B1(n_971),
.B2(n_964),
.C(n_958),
.Y(n_4078)
);

OAI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_3897),
.A2(n_975),
.B(n_974),
.Y(n_4079)
);

AOI21xp5_ASAP7_75t_L g4080 ( 
.A1(n_3775),
.A2(n_2221),
.B(n_2215),
.Y(n_4080)
);

OAI21x1_ASAP7_75t_L g4081 ( 
.A1(n_3886),
.A2(n_50),
.B(n_51),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3780),
.B(n_977),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3886),
.Y(n_4083)
);

CKINVDCx5p33_ASAP7_75t_R g4084 ( 
.A(n_3783),
.Y(n_4084)
);

BUFx2_ASAP7_75t_L g4085 ( 
.A(n_3963),
.Y(n_4085)
);

AOI221xp5_ASAP7_75t_L g4086 ( 
.A1(n_3871),
.A2(n_3864),
.B1(n_3887),
.B2(n_3868),
.C(n_3844),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3849),
.Y(n_4087)
);

CKINVDCx20_ASAP7_75t_R g4088 ( 
.A(n_3952),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3849),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3849),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3884),
.B(n_978),
.Y(n_4091)
);

OAI21x1_ASAP7_75t_L g4092 ( 
.A1(n_3959),
.A2(n_52),
.B(n_53),
.Y(n_4092)
);

AND2x2_ASAP7_75t_L g4093 ( 
.A(n_3898),
.B(n_52),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3768),
.Y(n_4094)
);

OA21x2_ASAP7_75t_L g4095 ( 
.A1(n_3779),
.A2(n_637),
.B(n_632),
.Y(n_4095)
);

OA21x2_ASAP7_75t_L g4096 ( 
.A1(n_3968),
.A2(n_650),
.B(n_643),
.Y(n_4096)
);

OAI21x1_ASAP7_75t_L g4097 ( 
.A1(n_3906),
.A2(n_3821),
.B(n_3909),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3773),
.Y(n_4098)
);

INVx2_ASAP7_75t_SL g4099 ( 
.A(n_3910),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3789),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3814),
.Y(n_4101)
);

AND2x4_ASAP7_75t_L g4102 ( 
.A(n_3828),
.B(n_54),
.Y(n_4102)
);

OAI221xp5_ASAP7_75t_L g4103 ( 
.A1(n_3839),
.A2(n_688),
.B1(n_698),
.B2(n_663),
.C(n_653),
.Y(n_4103)
);

OA21x2_ASAP7_75t_L g4104 ( 
.A1(n_3968),
.A2(n_713),
.B(n_712),
.Y(n_4104)
);

BUFx3_ASAP7_75t_L g4105 ( 
.A(n_3944),
.Y(n_4105)
);

OAI222xp33_ASAP7_75t_L g4106 ( 
.A1(n_3763),
.A2(n_755),
.B1(n_732),
.B2(n_760),
.C1(n_754),
.C2(n_720),
.Y(n_4106)
);

OAI21x1_ASAP7_75t_L g4107 ( 
.A1(n_3909),
.A2(n_54),
.B(n_55),
.Y(n_4107)
);

OAI21x1_ASAP7_75t_L g4108 ( 
.A1(n_3777),
.A2(n_56),
.B(n_59),
.Y(n_4108)
);

AOI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_3922),
.A2(n_2225),
.B(n_1735),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3765),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3810),
.Y(n_4111)
);

OAI22xp33_ASAP7_75t_L g4112 ( 
.A1(n_3865),
.A2(n_770),
.B1(n_778),
.B2(n_766),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3812),
.Y(n_4113)
);

BUFx3_ASAP7_75t_L g4114 ( 
.A(n_3834),
.Y(n_4114)
);

HB1xp67_ASAP7_75t_L g4115 ( 
.A(n_3970),
.Y(n_4115)
);

A2O1A1Ixp33_ASAP7_75t_L g4116 ( 
.A1(n_3835),
.A2(n_792),
.B(n_803),
.C(n_784),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_SL g4117 ( 
.A(n_3966),
.B(n_2225),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3784),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3838),
.Y(n_4119)
);

OAI22xp5_ASAP7_75t_L g4120 ( 
.A1(n_3967),
.A2(n_825),
.B1(n_832),
.B2(n_821),
.Y(n_4120)
);

OA21x2_ASAP7_75t_L g4121 ( 
.A1(n_3795),
.A2(n_875),
.B(n_849),
.Y(n_4121)
);

BUFx3_ASAP7_75t_L g4122 ( 
.A(n_3840),
.Y(n_4122)
);

OAI21x1_ASAP7_75t_SL g4123 ( 
.A1(n_3902),
.A2(n_59),
.B(n_60),
.Y(n_4123)
);

AND2x4_ASAP7_75t_L g4124 ( 
.A(n_3828),
.B(n_62),
.Y(n_4124)
);

AND2x4_ASAP7_75t_L g4125 ( 
.A(n_3965),
.B(n_3934),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_L g4126 ( 
.A1(n_3764),
.A2(n_1735),
.B1(n_885),
.B2(n_898),
.Y(n_4126)
);

OA21x2_ASAP7_75t_L g4127 ( 
.A1(n_3954),
.A2(n_917),
.B(n_882),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3799),
.B(n_62),
.Y(n_4128)
);

AOI22xp33_ASAP7_75t_L g4129 ( 
.A1(n_3764),
.A2(n_1735),
.B1(n_922),
.B2(n_929),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3815),
.Y(n_4130)
);

OAI21x1_ASAP7_75t_L g4131 ( 
.A1(n_3857),
.A2(n_3914),
.B(n_3750),
.Y(n_4131)
);

AND2x4_ASAP7_75t_L g4132 ( 
.A(n_3971),
.B(n_63),
.Y(n_4132)
);

A2O1A1Ixp33_ASAP7_75t_L g4133 ( 
.A1(n_3748),
.A2(n_930),
.B(n_938),
.C(n_918),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3878),
.Y(n_4134)
);

OAI22xp5_ASAP7_75t_L g4135 ( 
.A1(n_3782),
.A2(n_957),
.B1(n_972),
.B2(n_948),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_3837),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_3847),
.B(n_63),
.Y(n_4137)
);

OAI21x1_ASAP7_75t_L g4138 ( 
.A1(n_3750),
.A2(n_64),
.B(n_65),
.Y(n_4138)
);

INVx5_ASAP7_75t_L g4139 ( 
.A(n_3872),
.Y(n_4139)
);

OAI22xp5_ASAP7_75t_L g4140 ( 
.A1(n_3802),
.A2(n_1735),
.B1(n_67),
.B2(n_64),
.Y(n_4140)
);

BUFx3_ASAP7_75t_L g4141 ( 
.A(n_3840),
.Y(n_4141)
);

OA21x2_ASAP7_75t_L g4142 ( 
.A1(n_3903),
.A2(n_65),
.B(n_68),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3837),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_3961),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_3816),
.B(n_68),
.Y(n_4145)
);

OAI21x1_ASAP7_75t_L g4146 ( 
.A1(n_3969),
.A2(n_3801),
.B(n_3949),
.Y(n_4146)
);

OR2x6_ASAP7_75t_L g4147 ( 
.A(n_3896),
.B(n_1001),
.Y(n_4147)
);

O2A1O1Ixp33_ASAP7_75t_SL g4148 ( 
.A1(n_3867),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_4148)
);

INVx4_ASAP7_75t_SL g4149 ( 
.A(n_3912),
.Y(n_4149)
);

OAI21x1_ASAP7_75t_L g4150 ( 
.A1(n_3827),
.A2(n_71),
.B(n_72),
.Y(n_4150)
);

AOI22xp33_ASAP7_75t_L g4151 ( 
.A1(n_3848),
.A2(n_1735),
.B1(n_1125),
.B2(n_1126),
.Y(n_4151)
);

OR2x2_ASAP7_75t_L g4152 ( 
.A(n_3761),
.B(n_72),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_4024),
.B(n_4005),
.Y(n_4153)
);

INVx4_ASAP7_75t_L g4154 ( 
.A(n_4028),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_4043),
.Y(n_4155)
);

AOI21x1_ASAP7_75t_L g4156 ( 
.A1(n_4083),
.A2(n_3904),
.B(n_3892),
.Y(n_4156)
);

INVx4_ASAP7_75t_L g4157 ( 
.A(n_4028),
.Y(n_4157)
);

CKINVDCx5p33_ASAP7_75t_R g4158 ( 
.A(n_3978),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3975),
.Y(n_4159)
);

INVxp33_ASAP7_75t_SL g4160 ( 
.A(n_4015),
.Y(n_4160)
);

NAND2xp33_ASAP7_75t_R g4161 ( 
.A(n_4127),
.B(n_3905),
.Y(n_4161)
);

AND2x4_ASAP7_75t_L g4162 ( 
.A(n_3986),
.B(n_3971),
.Y(n_4162)
);

HB1xp67_ASAP7_75t_L g4163 ( 
.A(n_4115),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_4043),
.Y(n_4164)
);

AND2x2_ASAP7_75t_L g4165 ( 
.A(n_4085),
.B(n_3912),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3975),
.Y(n_4166)
);

OAI22xp5_ASAP7_75t_L g4167 ( 
.A1(n_3974),
.A2(n_3940),
.B1(n_3895),
.B2(n_3894),
.Y(n_4167)
);

AND2x4_ASAP7_75t_L g4168 ( 
.A(n_3995),
.B(n_3912),
.Y(n_4168)
);

INVx3_ASAP7_75t_L g4169 ( 
.A(n_3999),
.Y(n_4169)
);

AOI22xp33_ASAP7_75t_L g4170 ( 
.A1(n_4127),
.A2(n_3933),
.B1(n_3790),
.B2(n_3770),
.Y(n_4170)
);

AOI211xp5_ASAP7_75t_L g4171 ( 
.A1(n_4002),
.A2(n_3939),
.B(n_3951),
.C(n_3932),
.Y(n_4171)
);

AOI21xp33_ASAP7_75t_L g4172 ( 
.A1(n_3989),
.A2(n_3880),
.B(n_3859),
.Y(n_4172)
);

HB1xp67_ASAP7_75t_L g4173 ( 
.A(n_4051),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_SL g4174 ( 
.A1(n_4009),
.A2(n_3890),
.B1(n_3872),
.B2(n_3964),
.Y(n_4174)
);

OAI22xp5_ASAP7_75t_L g4175 ( 
.A1(n_4057),
.A2(n_3817),
.B1(n_3935),
.B2(n_3911),
.Y(n_4175)
);

BUFx2_ASAP7_75t_L g4176 ( 
.A(n_4014),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3979),
.Y(n_4177)
);

INVx2_ASAP7_75t_SL g4178 ( 
.A(n_4125),
.Y(n_4178)
);

AOI22xp5_ASAP7_75t_L g4179 ( 
.A1(n_4052),
.A2(n_3798),
.B1(n_3811),
.B2(n_3855),
.Y(n_4179)
);

OAI221xp5_ASAP7_75t_L g4180 ( 
.A1(n_4086),
.A2(n_3928),
.B1(n_3807),
.B2(n_3823),
.C(n_3901),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4051),
.Y(n_4181)
);

CKINVDCx9p33_ASAP7_75t_R g4182 ( 
.A(n_3977),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_SL g4183 ( 
.A1(n_4009),
.A2(n_3890),
.B1(n_3900),
.B2(n_3899),
.Y(n_4183)
);

AOI22xp33_ASAP7_75t_SL g4184 ( 
.A1(n_4121),
.A2(n_3883),
.B1(n_3771),
.B2(n_3875),
.Y(n_4184)
);

INVx3_ASAP7_75t_L g4185 ( 
.A(n_3999),
.Y(n_4185)
);

AOI211xp5_ASAP7_75t_L g4186 ( 
.A1(n_4036),
.A2(n_3800),
.B(n_3818),
.C(n_3825),
.Y(n_4186)
);

OAI22xp5_ASAP7_75t_L g4187 ( 
.A1(n_4018),
.A2(n_3858),
.B1(n_3822),
.B2(n_3794),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_3979),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4056),
.B(n_3961),
.Y(n_4189)
);

AOI22xp33_ASAP7_75t_L g4190 ( 
.A1(n_4121),
.A2(n_4095),
.B1(n_4035),
.B2(n_4096),
.Y(n_4190)
);

CKINVDCx5p33_ASAP7_75t_R g4191 ( 
.A(n_3981),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4056),
.B(n_3961),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4019),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_4066),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4019),
.Y(n_4195)
);

OR2x2_ASAP7_75t_L g4196 ( 
.A(n_4025),
.B(n_3957),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4125),
.B(n_3957),
.Y(n_4197)
);

OAI22xp33_ASAP7_75t_L g4198 ( 
.A1(n_4033),
.A2(n_3785),
.B1(n_3861),
.B2(n_3851),
.Y(n_4198)
);

AOI22xp33_ASAP7_75t_L g4199 ( 
.A1(n_4095),
.A2(n_3921),
.B1(n_3829),
.B2(n_3836),
.Y(n_4199)
);

CKINVDCx5p33_ASAP7_75t_R g4200 ( 
.A(n_3981),
.Y(n_4200)
);

AOI22xp33_ASAP7_75t_L g4201 ( 
.A1(n_4035),
.A2(n_3755),
.B1(n_3845),
.B2(n_3913),
.Y(n_4201)
);

AOI21x1_ASAP7_75t_L g4202 ( 
.A1(n_4083),
.A2(n_3796),
.B(n_3862),
.Y(n_4202)
);

A2O1A1Ixp33_ASAP7_75t_L g4203 ( 
.A1(n_4045),
.A2(n_3962),
.B(n_3893),
.C(n_3866),
.Y(n_4203)
);

NAND2xp33_ASAP7_75t_SL g4204 ( 
.A(n_4088),
.B(n_73),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_4099),
.B(n_3957),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4006),
.Y(n_4206)
);

INVx4_ASAP7_75t_L g4207 ( 
.A(n_4132),
.Y(n_4207)
);

OAI22xp33_ASAP7_75t_L g4208 ( 
.A1(n_4033),
.A2(n_3936),
.B1(n_3925),
.B2(n_1125),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4013),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_4105),
.B(n_3936),
.Y(n_4210)
);

AOI22xp33_ASAP7_75t_L g4211 ( 
.A1(n_4096),
.A2(n_1125),
.B1(n_1126),
.B2(n_1001),
.Y(n_4211)
);

AO21x2_ASAP7_75t_L g4212 ( 
.A1(n_4030),
.A2(n_4037),
.B(n_4077),
.Y(n_4212)
);

AND2x4_ASAP7_75t_L g4213 ( 
.A(n_4114),
.B(n_3925),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_4066),
.B(n_3936),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_4076),
.B(n_3925),
.Y(n_4215)
);

CKINVDCx11_ASAP7_75t_R g4216 ( 
.A(n_3988),
.Y(n_4216)
);

BUFx6f_ASAP7_75t_L g4217 ( 
.A(n_4147),
.Y(n_4217)
);

AOI221xp5_ASAP7_75t_L g4218 ( 
.A1(n_4148),
.A2(n_1126),
.B1(n_1228),
.B2(n_1125),
.C(n_1001),
.Y(n_4218)
);

OR2x6_ASAP7_75t_L g4219 ( 
.A(n_4070),
.B(n_1001),
.Y(n_4219)
);

AOI21xp5_ASAP7_75t_L g4220 ( 
.A1(n_4044),
.A2(n_73),
.B(n_74),
.Y(n_4220)
);

INVx3_ASAP7_75t_L g4221 ( 
.A(n_4008),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4021),
.Y(n_4222)
);

OAI221xp5_ASAP7_75t_L g4223 ( 
.A1(n_4042),
.A2(n_1126),
.B1(n_1228),
.B2(n_1125),
.C(n_1001),
.Y(n_4223)
);

OR2x2_ASAP7_75t_L g4224 ( 
.A(n_4111),
.B(n_4113),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4053),
.Y(n_4225)
);

NOR3xp33_ASAP7_75t_SL g4226 ( 
.A(n_4084),
.B(n_75),
.C(n_76),
.Y(n_4226)
);

CKINVDCx5p33_ASAP7_75t_R g4227 ( 
.A(n_4004),
.Y(n_4227)
);

AOI21xp33_ASAP7_75t_L g4228 ( 
.A1(n_4034),
.A2(n_75),
.B(n_76),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_4122),
.B(n_4141),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4053),
.Y(n_4230)
);

NOR2xp33_ASAP7_75t_L g4231 ( 
.A(n_4091),
.B(n_78),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4094),
.Y(n_4232)
);

AOI22xp33_ASAP7_75t_L g4233 ( 
.A1(n_4104),
.A2(n_1228),
.B1(n_1290),
.B2(n_1126),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_4027),
.B(n_78),
.Y(n_4234)
);

INVx1_ASAP7_75t_SL g4235 ( 
.A(n_4041),
.Y(n_4235)
);

NAND2xp33_ASAP7_75t_R g4236 ( 
.A(n_4132),
.B(n_4102),
.Y(n_4236)
);

OA21x2_ASAP7_75t_L g4237 ( 
.A1(n_4030),
.A2(n_79),
.B(n_80),
.Y(n_4237)
);

NOR2xp33_ASAP7_75t_SL g4238 ( 
.A(n_3987),
.B(n_3996),
.Y(n_4238)
);

INVx4_ASAP7_75t_L g4239 ( 
.A(n_4102),
.Y(n_4239)
);

BUFx12f_ASAP7_75t_L g4240 ( 
.A(n_4152),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_SL g4241 ( 
.A(n_4065),
.B(n_1228),
.Y(n_4241)
);

INVx1_ASAP7_75t_SL g4242 ( 
.A(n_4014),
.Y(n_4242)
);

OR2x6_ASAP7_75t_L g4243 ( 
.A(n_4070),
.B(n_1228),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4111),
.B(n_81),
.Y(n_4244)
);

AND2x2_ASAP7_75t_L g4245 ( 
.A(n_4149),
.B(n_81),
.Y(n_4245)
);

A2O1A1Ixp33_ASAP7_75t_L g4246 ( 
.A1(n_4049),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_4246)
);

OAI22xp5_ASAP7_75t_L g4247 ( 
.A1(n_4124),
.A2(n_4065),
.B1(n_4142),
.B2(n_4064),
.Y(n_4247)
);

NOR2xp33_ASAP7_75t_L g4248 ( 
.A(n_4137),
.B(n_83),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4094),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4098),
.Y(n_4250)
);

AND2x6_ASAP7_75t_L g4251 ( 
.A(n_4124),
.B(n_1290),
.Y(n_4251)
);

NOR2xp33_ASAP7_75t_L g4252 ( 
.A(n_4068),
.B(n_84),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4113),
.B(n_85),
.Y(n_4253)
);

INVx4_ASAP7_75t_L g4254 ( 
.A(n_4142),
.Y(n_4254)
);

INVx4_ASAP7_75t_R g4255 ( 
.A(n_4093),
.Y(n_4255)
);

BUFx4f_ASAP7_75t_SL g4256 ( 
.A(n_4069),
.Y(n_4256)
);

CKINVDCx11_ASAP7_75t_R g4257 ( 
.A(n_4008),
.Y(n_4257)
);

AOI22xp33_ASAP7_75t_L g4258 ( 
.A1(n_4104),
.A2(n_1290),
.B1(n_87),
.B2(n_85),
.Y(n_4258)
);

OAI211xp5_ASAP7_75t_SL g4259 ( 
.A1(n_4078),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_4063),
.A2(n_4080),
.B(n_4117),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_4149),
.B(n_88),
.Y(n_4261)
);

AOI22xp33_ASAP7_75t_SL g4262 ( 
.A1(n_3985),
.A2(n_1290),
.B1(n_91),
.B2(n_89),
.Y(n_4262)
);

NOR2x1_ASAP7_75t_SL g4263 ( 
.A(n_3998),
.B(n_1290),
.Y(n_4263)
);

NAND3xp33_ASAP7_75t_SL g4264 ( 
.A(n_4082),
.B(n_90),
.C(n_92),
.Y(n_4264)
);

OAI22xp5_ASAP7_75t_SL g4265 ( 
.A1(n_4022),
.A2(n_4145),
.B1(n_4128),
.B2(n_4047),
.Y(n_4265)
);

CKINVDCx5p33_ASAP7_75t_R g4266 ( 
.A(n_4008),
.Y(n_4266)
);

AOI22xp33_ASAP7_75t_L g4267 ( 
.A1(n_4126),
.A2(n_93),
.B1(n_90),
.B2(n_92),
.Y(n_4267)
);

INVx4_ASAP7_75t_L g4268 ( 
.A(n_4060),
.Y(n_4268)
);

A2O1A1Ixp33_ASAP7_75t_L g4269 ( 
.A1(n_4081),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_4269)
);

BUFx6f_ASAP7_75t_L g4270 ( 
.A(n_4147),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4031),
.Y(n_4271)
);

INVx3_ASAP7_75t_SL g4272 ( 
.A(n_4012),
.Y(n_4272)
);

BUFx3_ASAP7_75t_L g4273 ( 
.A(n_3993),
.Y(n_4273)
);

AOI22xp33_ASAP7_75t_L g4274 ( 
.A1(n_4129),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4098),
.Y(n_4275)
);

CKINVDCx5p33_ASAP7_75t_R g4276 ( 
.A(n_4012),
.Y(n_4276)
);

BUFx3_ASAP7_75t_L g4277 ( 
.A(n_4101),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4100),
.Y(n_4278)
);

HB1xp67_ASAP7_75t_L g4279 ( 
.A(n_4100),
.Y(n_4279)
);

AO21x2_ASAP7_75t_L g4280 ( 
.A1(n_4037),
.A2(n_97),
.B(n_98),
.Y(n_4280)
);

AOI22xp33_ASAP7_75t_SL g4281 ( 
.A1(n_4039),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_4281)
);

OR2x6_ASAP7_75t_L g4282 ( 
.A(n_4012),
.B(n_99),
.Y(n_4282)
);

AOI22xp33_ASAP7_75t_L g4283 ( 
.A1(n_3994),
.A2(n_4110),
.B1(n_4123),
.B2(n_4119),
.Y(n_4283)
);

CKINVDCx5p33_ASAP7_75t_R g4284 ( 
.A(n_4029),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4110),
.Y(n_4285)
);

BUFx6f_ASAP7_75t_L g4286 ( 
.A(n_4150),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4075),
.B(n_101),
.Y(n_4287)
);

AND2x4_ASAP7_75t_L g4288 ( 
.A(n_4139),
.B(n_102),
.Y(n_4288)
);

INVx2_ASAP7_75t_L g4289 ( 
.A(n_4062),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_4118),
.B(n_102),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_4130),
.B(n_103),
.Y(n_4291)
);

AOI21x1_ASAP7_75t_L g4292 ( 
.A1(n_4046),
.A2(n_105),
.B(n_106),
.Y(n_4292)
);

OAI222xp33_ASAP7_75t_L g4293 ( 
.A1(n_4134),
.A2(n_4143),
.B1(n_4048),
.B2(n_4059),
.C1(n_4050),
.C2(n_3976),
.Y(n_4293)
);

OAI22xp33_ASAP7_75t_L g4294 ( 
.A1(n_4139),
.A2(n_109),
.B1(n_106),
.B2(n_107),
.Y(n_4294)
);

OAI22xp33_ASAP7_75t_L g4295 ( 
.A1(n_4254),
.A2(n_4139),
.B1(n_4061),
.B2(n_4140),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4225),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_SL g4297 ( 
.A(n_4247),
.B(n_4029),
.Y(n_4297)
);

OAI211xp5_ASAP7_75t_L g4298 ( 
.A1(n_4226),
.A2(n_4079),
.B(n_4071),
.C(n_4016),
.Y(n_4298)
);

BUFx12f_ASAP7_75t_L g4299 ( 
.A(n_4216),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4194),
.Y(n_4300)
);

INVx3_ASAP7_75t_L g4301 ( 
.A(n_4207),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_4254),
.B(n_3973),
.Y(n_4302)
);

AOI22xp33_ASAP7_75t_L g4303 ( 
.A1(n_4190),
.A2(n_3994),
.B1(n_4058),
.B2(n_4143),
.Y(n_4303)
);

OAI22xp33_ASAP7_75t_L g4304 ( 
.A1(n_4161),
.A2(n_4029),
.B1(n_4000),
.B2(n_4017),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4169),
.B(n_4026),
.Y(n_4305)
);

NAND3xp33_ASAP7_75t_L g4306 ( 
.A(n_4220),
.B(n_4120),
.C(n_3980),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4230),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_4224),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_4163),
.B(n_4007),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4279),
.Y(n_4310)
);

AOI22xp33_ASAP7_75t_L g4311 ( 
.A1(n_4265),
.A2(n_4001),
.B1(n_4144),
.B2(n_4089),
.Y(n_4311)
);

AOI22xp33_ASAP7_75t_L g4312 ( 
.A1(n_4167),
.A2(n_4001),
.B1(n_4089),
.B2(n_4087),
.Y(n_4312)
);

OA21x2_ASAP7_75t_L g4313 ( 
.A1(n_4293),
.A2(n_4136),
.B(n_4090),
.Y(n_4313)
);

CKINVDCx6p67_ASAP7_75t_R g4314 ( 
.A(n_4282),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4277),
.B(n_4007),
.Y(n_4315)
);

AOI21xp5_ASAP7_75t_L g4316 ( 
.A1(n_4198),
.A2(n_4109),
.B(n_4133),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4232),
.Y(n_4317)
);

AOI211xp5_ASAP7_75t_L g4318 ( 
.A1(n_4204),
.A2(n_4112),
.B(n_4116),
.C(n_4106),
.Y(n_4318)
);

CKINVDCx20_ASAP7_75t_R g4319 ( 
.A(n_4158),
.Y(n_4319)
);

AOI22xp33_ASAP7_75t_L g4320 ( 
.A1(n_4237),
.A2(n_4087),
.B1(n_4090),
.B2(n_4138),
.Y(n_4320)
);

INVxp67_ASAP7_75t_L g4321 ( 
.A(n_4236),
.Y(n_4321)
);

AND2x2_ASAP7_75t_L g4322 ( 
.A(n_4169),
.B(n_3982),
.Y(n_4322)
);

OAI221xp5_ASAP7_75t_L g4323 ( 
.A1(n_4174),
.A2(n_4135),
.B1(n_4103),
.B2(n_4038),
.C(n_4151),
.Y(n_4323)
);

CKINVDCx20_ASAP7_75t_R g4324 ( 
.A(n_4257),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4173),
.B(n_4007),
.Y(n_4325)
);

AOI22xp33_ASAP7_75t_L g4326 ( 
.A1(n_4237),
.A2(n_4107),
.B1(n_4055),
.B2(n_4067),
.Y(n_4326)
);

AND2x4_ASAP7_75t_L g4327 ( 
.A(n_4239),
.B(n_3991),
.Y(n_4327)
);

INVx2_ASAP7_75t_SL g4328 ( 
.A(n_4255),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4249),
.Y(n_4329)
);

BUFx3_ASAP7_75t_L g4330 ( 
.A(n_4160),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_4206),
.B(n_4072),
.Y(n_4331)
);

OA21x2_ASAP7_75t_L g4332 ( 
.A1(n_4271),
.A2(n_4097),
.B(n_4131),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4209),
.B(n_4108),
.Y(n_4333)
);

OAI22xp5_ASAP7_75t_SL g4334 ( 
.A1(n_4256),
.A2(n_4040),
.B1(n_4074),
.B2(n_4073),
.Y(n_4334)
);

AO21x2_ASAP7_75t_L g4335 ( 
.A1(n_4212),
.A2(n_4291),
.B(n_4290),
.Y(n_4335)
);

AOI22xp33_ASAP7_75t_L g4336 ( 
.A1(n_4280),
.A2(n_4054),
.B1(n_3997),
.B2(n_4146),
.Y(n_4336)
);

INVx2_ASAP7_75t_L g4337 ( 
.A(n_4155),
.Y(n_4337)
);

AOI22xp33_ASAP7_75t_SL g4338 ( 
.A1(n_4280),
.A2(n_4003),
.B1(n_3992),
.B2(n_3983),
.Y(n_4338)
);

OR2x6_ASAP7_75t_L g4339 ( 
.A(n_4288),
.B(n_3984),
.Y(n_4339)
);

BUFx8_ASAP7_75t_L g4340 ( 
.A(n_4245),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_4222),
.B(n_4092),
.Y(n_4341)
);

AOI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_4241),
.A2(n_4032),
.B(n_4011),
.Y(n_4342)
);

OAI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_4248),
.A2(n_4010),
.B(n_4023),
.Y(n_4343)
);

OAI211xp5_ASAP7_75t_L g4344 ( 
.A1(n_4281),
.A2(n_111),
.B(n_107),
.C(n_110),
.Y(n_4344)
);

AOI22xp33_ASAP7_75t_L g4345 ( 
.A1(n_4286),
.A2(n_4020),
.B1(n_3990),
.B2(n_115),
.Y(n_4345)
);

O2A1O1Ixp33_ASAP7_75t_L g4346 ( 
.A1(n_4246),
.A2(n_116),
.B(n_113),
.C(n_114),
.Y(n_4346)
);

AO21x2_ASAP7_75t_L g4347 ( 
.A1(n_4212),
.A2(n_3990),
.B(n_114),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4164),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4250),
.Y(n_4349)
);

AO21x2_ASAP7_75t_L g4350 ( 
.A1(n_4244),
.A2(n_3990),
.B(n_116),
.Y(n_4350)
);

AOI21xp5_ASAP7_75t_L g4351 ( 
.A1(n_4260),
.A2(n_4288),
.B(n_4243),
.Y(n_4351)
);

OR2x2_ASAP7_75t_L g4352 ( 
.A(n_4153),
.B(n_117),
.Y(n_4352)
);

AOI22xp33_ASAP7_75t_L g4353 ( 
.A1(n_4286),
.A2(n_122),
.B1(n_119),
.B2(n_121),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_4207),
.A2(n_123),
.B1(n_119),
.B2(n_121),
.Y(n_4354)
);

OAI221xp5_ASAP7_75t_L g4355 ( 
.A1(n_4283),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.C(n_128),
.Y(n_4355)
);

OAI22xp5_ASAP7_75t_L g4356 ( 
.A1(n_4239),
.A2(n_134),
.B1(n_128),
.B2(n_129),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4275),
.Y(n_4357)
);

INVx2_ASAP7_75t_L g4358 ( 
.A(n_4181),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4185),
.B(n_137),
.Y(n_4359)
);

AOI22xp5_ASAP7_75t_L g4360 ( 
.A1(n_4179),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_4278),
.B(n_138),
.Y(n_4361)
);

OR2x6_ASAP7_75t_L g4362 ( 
.A(n_4282),
.B(n_140),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4285),
.Y(n_4363)
);

AND2x2_ASAP7_75t_L g4364 ( 
.A(n_4185),
.B(n_141),
.Y(n_4364)
);

OAI22xp5_ASAP7_75t_L g4365 ( 
.A1(n_4268),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4205),
.Y(n_4366)
);

OAI211xp5_ASAP7_75t_SL g4367 ( 
.A1(n_4171),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_4367)
);

AOI221xp5_ASAP7_75t_L g4368 ( 
.A1(n_4264),
.A2(n_149),
.B1(n_146),
.B2(n_148),
.C(n_150),
.Y(n_4368)
);

INVx1_ASAP7_75t_SL g4369 ( 
.A(n_4182),
.Y(n_4369)
);

OAI22xp5_ASAP7_75t_L g4370 ( 
.A1(n_4268),
.A2(n_151),
.B1(n_148),
.B2(n_150),
.Y(n_4370)
);

CKINVDCx5p33_ASAP7_75t_R g4371 ( 
.A(n_4191),
.Y(n_4371)
);

OR2x2_ASAP7_75t_L g4372 ( 
.A(n_4178),
.B(n_155),
.Y(n_4372)
);

OAI221xp5_ASAP7_75t_L g4373 ( 
.A1(n_4258),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.C(n_159),
.Y(n_4373)
);

AOI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_4219),
.A2(n_4243),
.B(n_4186),
.Y(n_4374)
);

OA21x2_ASAP7_75t_L g4375 ( 
.A1(n_4289),
.A2(n_156),
.B(n_157),
.Y(n_4375)
);

BUFx12f_ASAP7_75t_L g4376 ( 
.A(n_4200),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4286),
.A2(n_4184),
.B1(n_4170),
.B2(n_4183),
.Y(n_4377)
);

AOI21xp5_ASAP7_75t_L g4378 ( 
.A1(n_4219),
.A2(n_159),
.B(n_161),
.Y(n_4378)
);

NAND4xp25_ASAP7_75t_L g4379 ( 
.A(n_4273),
.B(n_166),
.C(n_163),
.D(n_165),
.Y(n_4379)
);

OR3x1_ASAP7_75t_L g4380 ( 
.A(n_4255),
.B(n_4228),
.C(n_4231),
.Y(n_4380)
);

BUFx2_ASAP7_75t_L g4381 ( 
.A(n_4162),
.Y(n_4381)
);

AOI22xp5_ASAP7_75t_L g4382 ( 
.A1(n_4179),
.A2(n_167),
.B1(n_163),
.B2(n_166),
.Y(n_4382)
);

AND2x2_ASAP7_75t_L g4383 ( 
.A(n_4165),
.B(n_168),
.Y(n_4383)
);

AND2x4_ASAP7_75t_L g4384 ( 
.A(n_4176),
.B(n_170),
.Y(n_4384)
);

AND2x4_ASAP7_75t_L g4385 ( 
.A(n_4162),
.B(n_170),
.Y(n_4385)
);

AOI222xp33_ASAP7_75t_L g4386 ( 
.A1(n_4287),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.C1(n_175),
.C2(n_176),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_SL g4387 ( 
.A1(n_4240),
.A2(n_178),
.B1(n_173),
.B2(n_176),
.Y(n_4387)
);

AO31x2_ASAP7_75t_L g4388 ( 
.A1(n_4189),
.A2(n_184),
.A3(n_180),
.B(n_181),
.Y(n_4388)
);

OAI221xp5_ASAP7_75t_L g4389 ( 
.A1(n_4269),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.C(n_189),
.Y(n_4389)
);

AND2x2_ASAP7_75t_L g4390 ( 
.A(n_4168),
.B(n_190),
.Y(n_4390)
);

AO21x2_ASAP7_75t_L g4391 ( 
.A1(n_4253),
.A2(n_190),
.B(n_191),
.Y(n_4391)
);

CKINVDCx5p33_ASAP7_75t_R g4392 ( 
.A(n_4154),
.Y(n_4392)
);

BUFx6f_ASAP7_75t_L g4393 ( 
.A(n_4217),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_4294),
.A2(n_191),
.B(n_192),
.Y(n_4394)
);

OAI211xp5_ASAP7_75t_L g4395 ( 
.A1(n_4252),
.A2(n_195),
.B(n_192),
.C(n_193),
.Y(n_4395)
);

A2O1A1Ixp33_ASAP7_75t_L g4396 ( 
.A1(n_4261),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_L g4397 ( 
.A(n_4159),
.B(n_196),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4166),
.Y(n_4398)
);

AOI22xp33_ASAP7_75t_L g4399 ( 
.A1(n_4259),
.A2(n_201),
.B1(n_198),
.B2(n_199),
.Y(n_4399)
);

CKINVDCx6p67_ASAP7_75t_R g4400 ( 
.A(n_4154),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_4177),
.B(n_201),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_4188),
.B(n_4193),
.Y(n_4402)
);

OAI221xp5_ASAP7_75t_SL g4403 ( 
.A1(n_4267),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.C(n_207),
.Y(n_4403)
);

OAI221xp5_ASAP7_75t_SL g4404 ( 
.A1(n_4274),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.C(n_211),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4195),
.Y(n_4405)
);

AOI22xp33_ASAP7_75t_L g4406 ( 
.A1(n_4199),
.A2(n_4218),
.B1(n_4180),
.B2(n_4172),
.Y(n_4406)
);

BUFx3_ASAP7_75t_L g4407 ( 
.A(n_4227),
.Y(n_4407)
);

AOI22xp33_ASAP7_75t_SL g4408 ( 
.A1(n_4238),
.A2(n_211),
.B1(n_208),
.B2(n_209),
.Y(n_4408)
);

INVx2_ASAP7_75t_L g4409 ( 
.A(n_4197),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4234),
.Y(n_4410)
);

HB1xp67_ASAP7_75t_L g4411 ( 
.A(n_4196),
.Y(n_4411)
);

INVx3_ASAP7_75t_L g4412 ( 
.A(n_4168),
.Y(n_4412)
);

OAI22xp33_ASAP7_75t_L g4413 ( 
.A1(n_4156),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_4413)
);

AOI221xp5_ASAP7_75t_L g4414 ( 
.A1(n_4192),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.C(n_217),
.Y(n_4414)
);

AOI22xp33_ASAP7_75t_L g4415 ( 
.A1(n_4211),
.A2(n_221),
.B1(n_218),
.B2(n_219),
.Y(n_4415)
);

A2O1A1Ixp33_ASAP7_75t_L g4416 ( 
.A1(n_4235),
.A2(n_226),
.B(n_221),
.C(n_222),
.Y(n_4416)
);

AOI22xp33_ASAP7_75t_L g4417 ( 
.A1(n_4233),
.A2(n_228),
.B1(n_222),
.B2(n_226),
.Y(n_4417)
);

OAI22xp5_ASAP7_75t_L g4418 ( 
.A1(n_4242),
.A2(n_231),
.B1(n_228),
.B2(n_230),
.Y(n_4418)
);

BUFx3_ASAP7_75t_L g4419 ( 
.A(n_4157),
.Y(n_4419)
);

OAI22xp5_ASAP7_75t_L g4420 ( 
.A1(n_4262),
.A2(n_234),
.B1(n_230),
.B2(n_233),
.Y(n_4420)
);

INVx4_ASAP7_75t_SL g4421 ( 
.A(n_4251),
.Y(n_4421)
);

OAI22xp33_ASAP7_75t_L g4422 ( 
.A1(n_4217),
.A2(n_4270),
.B1(n_4292),
.B2(n_4272),
.Y(n_4422)
);

OAI22xp5_ASAP7_75t_L g4423 ( 
.A1(n_4266),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_4423)
);

OAI211xp5_ASAP7_75t_SL g4424 ( 
.A1(n_4175),
.A2(n_239),
.B(n_236),
.C(n_237),
.Y(n_4424)
);

AND2x2_ASAP7_75t_L g4425 ( 
.A(n_4229),
.B(n_239),
.Y(n_4425)
);

OAI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_4210),
.A2(n_240),
.B(n_241),
.Y(n_4426)
);

NAND2xp33_ASAP7_75t_R g4427 ( 
.A(n_4362),
.B(n_4276),
.Y(n_4427)
);

AND2x2_ASAP7_75t_L g4428 ( 
.A(n_4381),
.B(n_4284),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_4335),
.B(n_4251),
.Y(n_4429)
);

NOR2xp33_ASAP7_75t_R g4430 ( 
.A(n_4299),
.B(n_4157),
.Y(n_4430)
);

AND2x4_ASAP7_75t_L g4431 ( 
.A(n_4328),
.B(n_4251),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_SL g4432 ( 
.A(n_4369),
.B(n_4217),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_4335),
.B(n_4251),
.Y(n_4433)
);

BUFx3_ASAP7_75t_L g4434 ( 
.A(n_4324),
.Y(n_4434)
);

NOR2xp33_ASAP7_75t_R g4435 ( 
.A(n_4319),
.B(n_4221),
.Y(n_4435)
);

NAND2xp33_ASAP7_75t_R g4436 ( 
.A(n_4362),
.B(n_4221),
.Y(n_4436)
);

CKINVDCx5p33_ASAP7_75t_R g4437 ( 
.A(n_4376),
.Y(n_4437)
);

NOR2xp33_ASAP7_75t_R g4438 ( 
.A(n_4392),
.B(n_242),
.Y(n_4438)
);

NAND2xp33_ASAP7_75t_SL g4439 ( 
.A(n_4385),
.B(n_4270),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4296),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4301),
.B(n_4270),
.Y(n_4441)
);

NOR2xp33_ASAP7_75t_R g4442 ( 
.A(n_4371),
.B(n_242),
.Y(n_4442)
);

AND2x4_ASAP7_75t_L g4443 ( 
.A(n_4301),
.B(n_4202),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_4375),
.Y(n_4444)
);

OR2x6_ASAP7_75t_L g4445 ( 
.A(n_4384),
.B(n_4203),
.Y(n_4445)
);

NAND2xp33_ASAP7_75t_R g4446 ( 
.A(n_4384),
.B(n_4213),
.Y(n_4446)
);

NOR2xp33_ASAP7_75t_R g4447 ( 
.A(n_4330),
.B(n_243),
.Y(n_4447)
);

NOR2xp33_ASAP7_75t_R g4448 ( 
.A(n_4400),
.B(n_243),
.Y(n_4448)
);

NAND2xp33_ASAP7_75t_R g4449 ( 
.A(n_4385),
.B(n_4213),
.Y(n_4449)
);

AND2x4_ASAP7_75t_L g4450 ( 
.A(n_4321),
.B(n_4215),
.Y(n_4450)
);

NAND2x1p5_ASAP7_75t_L g4451 ( 
.A(n_4407),
.B(n_4263),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4307),
.Y(n_4452)
);

INVx2_ASAP7_75t_L g4453 ( 
.A(n_4375),
.Y(n_4453)
);

AND2x4_ASAP7_75t_L g4454 ( 
.A(n_4327),
.B(n_4214),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4305),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_SL g4456 ( 
.A(n_4351),
.B(n_4187),
.Y(n_4456)
);

INVxp67_ASAP7_75t_L g4457 ( 
.A(n_4391),
.Y(n_4457)
);

OR2x6_ASAP7_75t_L g4458 ( 
.A(n_4425),
.B(n_4201),
.Y(n_4458)
);

NAND2xp33_ASAP7_75t_R g4459 ( 
.A(n_4359),
.B(n_244),
.Y(n_4459)
);

NAND2xp33_ASAP7_75t_R g4460 ( 
.A(n_4364),
.B(n_244),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_4410),
.B(n_4208),
.Y(n_4461)
);

NAND2xp33_ASAP7_75t_R g4462 ( 
.A(n_4390),
.B(n_4383),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_L g4463 ( 
.A(n_4391),
.B(n_4388),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4388),
.B(n_4223),
.Y(n_4464)
);

AND2x4_ASAP7_75t_L g4465 ( 
.A(n_4327),
.B(n_245),
.Y(n_4465)
);

NAND2xp33_ASAP7_75t_R g4466 ( 
.A(n_4372),
.B(n_245),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4388),
.B(n_246),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4317),
.Y(n_4468)
);

INVx2_ASAP7_75t_SL g4469 ( 
.A(n_4340),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4329),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_SL g4471 ( 
.A(n_4304),
.B(n_246),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4349),
.Y(n_4472)
);

BUFx3_ASAP7_75t_L g4473 ( 
.A(n_4340),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_SL g4474 ( 
.A(n_4422),
.B(n_247),
.Y(n_4474)
);

NOR2xp33_ASAP7_75t_L g4475 ( 
.A(n_4314),
.B(n_248),
.Y(n_4475)
);

XNOR2xp5_ASAP7_75t_L g4476 ( 
.A(n_4380),
.B(n_249),
.Y(n_4476)
);

XNOR2xp5_ASAP7_75t_L g4477 ( 
.A(n_4379),
.B(n_250),
.Y(n_4477)
);

CKINVDCx20_ASAP7_75t_R g4478 ( 
.A(n_4419),
.Y(n_4478)
);

OR2x2_ASAP7_75t_L g4479 ( 
.A(n_4308),
.B(n_251),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4310),
.B(n_253),
.Y(n_4480)
);

NOR2xp33_ASAP7_75t_R g4481 ( 
.A(n_4352),
.B(n_4361),
.Y(n_4481)
);

HB1xp67_ASAP7_75t_L g4482 ( 
.A(n_4357),
.Y(n_4482)
);

AND2x2_ASAP7_75t_L g4483 ( 
.A(n_4412),
.B(n_4297),
.Y(n_4483)
);

AND2x4_ASAP7_75t_L g4484 ( 
.A(n_4412),
.B(n_253),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_4322),
.B(n_254),
.Y(n_4485)
);

NAND2xp33_ASAP7_75t_R g4486 ( 
.A(n_4374),
.B(n_254),
.Y(n_4486)
);

AND2x4_ASAP7_75t_L g4487 ( 
.A(n_4339),
.B(n_255),
.Y(n_4487)
);

OR2x6_ASAP7_75t_L g4488 ( 
.A(n_4426),
.B(n_255),
.Y(n_4488)
);

AND2x4_ASAP7_75t_L g4489 ( 
.A(n_4339),
.B(n_256),
.Y(n_4489)
);

XNOR2xp5_ASAP7_75t_L g4490 ( 
.A(n_4360),
.B(n_256),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_SL g4491 ( 
.A(n_4295),
.B(n_4393),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4331),
.B(n_4333),
.Y(n_4492)
);

OR2x6_ASAP7_75t_L g4493 ( 
.A(n_4316),
.B(n_257),
.Y(n_4493)
);

NAND2xp33_ASAP7_75t_R g4494 ( 
.A(n_4313),
.B(n_257),
.Y(n_4494)
);

XNOR2xp5_ASAP7_75t_L g4495 ( 
.A(n_4360),
.B(n_260),
.Y(n_4495)
);

NAND2xp33_ASAP7_75t_SL g4496 ( 
.A(n_4377),
.B(n_261),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4363),
.Y(n_4497)
);

INVxp67_ASAP7_75t_L g4498 ( 
.A(n_4393),
.Y(n_4498)
);

NAND2x1p5_ASAP7_75t_L g4499 ( 
.A(n_4393),
.B(n_262),
.Y(n_4499)
);

INVxp67_ASAP7_75t_L g4500 ( 
.A(n_4397),
.Y(n_4500)
);

NAND2xp33_ASAP7_75t_R g4501 ( 
.A(n_4313),
.B(n_262),
.Y(n_4501)
);

AND2x4_ASAP7_75t_L g4502 ( 
.A(n_4421),
.B(n_263),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4300),
.Y(n_4503)
);

NAND2xp33_ASAP7_75t_R g4504 ( 
.A(n_4401),
.B(n_263),
.Y(n_4504)
);

OR2x4_ASAP7_75t_L g4505 ( 
.A(n_4302),
.B(n_264),
.Y(n_4505)
);

INVxp67_ASAP7_75t_L g4506 ( 
.A(n_4334),
.Y(n_4506)
);

AND2x4_ASAP7_75t_L g4507 ( 
.A(n_4421),
.B(n_264),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4398),
.B(n_4405),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4341),
.B(n_265),
.Y(n_4509)
);

AND2x2_ASAP7_75t_L g4510 ( 
.A(n_4409),
.B(n_265),
.Y(n_4510)
);

NAND2xp33_ASAP7_75t_R g4511 ( 
.A(n_4315),
.B(n_266),
.Y(n_4511)
);

NAND2xp33_ASAP7_75t_R g4512 ( 
.A(n_4309),
.B(n_267),
.Y(n_4512)
);

XNOR2xp5_ASAP7_75t_L g4513 ( 
.A(n_4382),
.B(n_267),
.Y(n_4513)
);

BUFx3_ASAP7_75t_L g4514 ( 
.A(n_4382),
.Y(n_4514)
);

AND2x2_ASAP7_75t_L g4515 ( 
.A(n_4402),
.B(n_268),
.Y(n_4515)
);

NAND2xp33_ASAP7_75t_R g4516 ( 
.A(n_4394),
.B(n_269),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4406),
.B(n_270),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_L g4518 ( 
.A(n_4350),
.B(n_270),
.Y(n_4518)
);

OR2x6_ASAP7_75t_L g4519 ( 
.A(n_4378),
.B(n_271),
.Y(n_4519)
);

BUFx3_ASAP7_75t_L g4520 ( 
.A(n_4334),
.Y(n_4520)
);

NOR2xp33_ASAP7_75t_R g4521 ( 
.A(n_4353),
.B(n_272),
.Y(n_4521)
);

NOR2xp33_ASAP7_75t_R g4522 ( 
.A(n_4399),
.B(n_273),
.Y(n_4522)
);

AND2x2_ASAP7_75t_L g4523 ( 
.A(n_4366),
.B(n_4337),
.Y(n_4523)
);

CKINVDCx20_ASAP7_75t_R g4524 ( 
.A(n_4418),
.Y(n_4524)
);

NAND2xp33_ASAP7_75t_R g4525 ( 
.A(n_4343),
.B(n_273),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_4348),
.B(n_274),
.Y(n_4526)
);

BUFx10_ASAP7_75t_L g4527 ( 
.A(n_4387),
.Y(n_4527)
);

NOR2xp33_ASAP7_75t_R g4528 ( 
.A(n_4298),
.B(n_274),
.Y(n_4528)
);

NAND2xp33_ASAP7_75t_R g4529 ( 
.A(n_4325),
.B(n_275),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4350),
.B(n_275),
.Y(n_4530)
);

HB1xp67_ASAP7_75t_L g4531 ( 
.A(n_4482),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4440),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4514),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4452),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_4444),
.Y(n_4535)
);

HB1xp67_ASAP7_75t_L g4536 ( 
.A(n_4500),
.Y(n_4536)
);

NOR2xp67_ASAP7_75t_L g4537 ( 
.A(n_4506),
.B(n_4469),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_4453),
.Y(n_4538)
);

OAI22xp33_ASAP7_75t_L g4539 ( 
.A1(n_4505),
.A2(n_4355),
.B1(n_4306),
.B2(n_4411),
.Y(n_4539)
);

INVxp67_ASAP7_75t_SL g4540 ( 
.A(n_4520),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4515),
.B(n_4457),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4483),
.B(n_4358),
.Y(n_4542)
);

AND2x2_ASAP7_75t_L g4543 ( 
.A(n_4431),
.B(n_4311),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_4527),
.Y(n_4544)
);

BUFx3_ASAP7_75t_L g4545 ( 
.A(n_4473),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4468),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4470),
.Y(n_4547)
);

AND2x2_ASAP7_75t_L g4548 ( 
.A(n_4431),
.B(n_4303),
.Y(n_4548)
);

OR2x2_ASAP7_75t_L g4549 ( 
.A(n_4508),
.B(n_4326),
.Y(n_4549)
);

NOR2x1_ASAP7_75t_L g4550 ( 
.A(n_4493),
.B(n_4424),
.Y(n_4550)
);

HB1xp67_ASAP7_75t_L g4551 ( 
.A(n_4472),
.Y(n_4551)
);

INVx2_ASAP7_75t_L g4552 ( 
.A(n_4493),
.Y(n_4552)
);

NOR2xp33_ASAP7_75t_L g4553 ( 
.A(n_4434),
.B(n_4395),
.Y(n_4553)
);

AOI221xp5_ASAP7_75t_L g4554 ( 
.A1(n_4463),
.A2(n_4413),
.B1(n_4346),
.B2(n_4389),
.C(n_4367),
.Y(n_4554)
);

OR2x2_ASAP7_75t_L g4555 ( 
.A(n_4497),
.B(n_4336),
.Y(n_4555)
);

OR2x2_ASAP7_75t_L g4556 ( 
.A(n_4492),
.B(n_4320),
.Y(n_4556)
);

AND2x2_ASAP7_75t_L g4557 ( 
.A(n_4441),
.B(n_4365),
.Y(n_4557)
);

OR2x2_ASAP7_75t_L g4558 ( 
.A(n_4509),
.B(n_4312),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4487),
.B(n_4414),
.Y(n_4559)
);

OR2x2_ASAP7_75t_L g4560 ( 
.A(n_4467),
.B(n_4332),
.Y(n_4560)
);

INVx2_ASAP7_75t_L g4561 ( 
.A(n_4445),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4518),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_4445),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_4530),
.Y(n_4564)
);

INVx3_ASAP7_75t_L g4565 ( 
.A(n_4443),
.Y(n_4565)
);

AND2x2_ASAP7_75t_L g4566 ( 
.A(n_4428),
.B(n_4370),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4479),
.Y(n_4567)
);

AND2x4_ASAP7_75t_SL g4568 ( 
.A(n_4465),
.B(n_4345),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4480),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_4465),
.B(n_4332),
.Y(n_4570)
);

OR2x2_ASAP7_75t_L g4571 ( 
.A(n_4458),
.B(n_4356),
.Y(n_4571)
);

HB1xp67_ASAP7_75t_L g4572 ( 
.A(n_4485),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_4455),
.B(n_4354),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4487),
.B(n_4386),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4526),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_4498),
.B(n_4338),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_4519),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4503),
.Y(n_4578)
);

BUFx6f_ASAP7_75t_L g4579 ( 
.A(n_4517),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4523),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4456),
.B(n_4342),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4519),
.Y(n_4582)
);

AND2x2_ASAP7_75t_L g4583 ( 
.A(n_4489),
.B(n_4416),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4489),
.B(n_4408),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4458),
.B(n_4450),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4484),
.B(n_4396),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4450),
.B(n_4368),
.Y(n_4587)
);

BUFx6f_ASAP7_75t_L g4588 ( 
.A(n_4502),
.Y(n_4588)
);

OR2x2_ASAP7_75t_L g4589 ( 
.A(n_4461),
.B(n_4347),
.Y(n_4589)
);

INVx2_ASAP7_75t_L g4590 ( 
.A(n_4429),
.Y(n_4590)
);

AND2x2_ASAP7_75t_L g4591 ( 
.A(n_4454),
.B(n_4423),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4454),
.B(n_4347),
.Y(n_4592)
);

INVx2_ASAP7_75t_L g4593 ( 
.A(n_4433),
.Y(n_4593)
);

AO21x2_ASAP7_75t_L g4594 ( 
.A1(n_4464),
.A2(n_4373),
.B(n_4420),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4432),
.B(n_4318),
.Y(n_4595)
);

HB1xp67_ASAP7_75t_L g4596 ( 
.A(n_4481),
.Y(n_4596)
);

HB1xp67_ASAP7_75t_L g4597 ( 
.A(n_4462),
.Y(n_4597)
);

INVx2_ASAP7_75t_L g4598 ( 
.A(n_4488),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4510),
.Y(n_4599)
);

HB1xp67_ASAP7_75t_L g4600 ( 
.A(n_4436),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_L g4601 ( 
.A(n_4484),
.B(n_4318),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4488),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4443),
.B(n_4344),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_4490),
.Y(n_4604)
);

INVxp67_ASAP7_75t_SL g4605 ( 
.A(n_4504),
.Y(n_4605)
);

AND2x2_ASAP7_75t_L g4606 ( 
.A(n_4435),
.B(n_4415),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4566),
.B(n_4430),
.Y(n_4607)
);

OAI21xp5_ASAP7_75t_L g4608 ( 
.A1(n_4550),
.A2(n_4605),
.B(n_4595),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4566),
.B(n_4478),
.Y(n_4609)
);

NOR3xp33_ASAP7_75t_L g4610 ( 
.A(n_4544),
.B(n_4475),
.C(n_4404),
.Y(n_4610)
);

OAI21xp33_ASAP7_75t_SL g4611 ( 
.A1(n_4581),
.A2(n_4491),
.B(n_4474),
.Y(n_4611)
);

NAND2xp5_ASAP7_75t_L g4612 ( 
.A(n_4599),
.B(n_4476),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4581),
.B(n_4437),
.Y(n_4613)
);

OAI22xp5_ASAP7_75t_L g4614 ( 
.A1(n_4597),
.A2(n_4524),
.B1(n_4471),
.B2(n_4477),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_L g4615 ( 
.A(n_4599),
.B(n_4502),
.Y(n_4615)
);

AOI21xp5_ASAP7_75t_L g4616 ( 
.A1(n_4539),
.A2(n_4496),
.B(n_4439),
.Y(n_4616)
);

NOR2x1p5_ASAP7_75t_L g4617 ( 
.A(n_4545),
.B(n_4507),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_4572),
.B(n_4536),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_4583),
.B(n_4507),
.Y(n_4619)
);

OAI22xp33_ASAP7_75t_L g4620 ( 
.A1(n_4571),
.A2(n_4529),
.B1(n_4512),
.B2(n_4525),
.Y(n_4620)
);

AND2x2_ASAP7_75t_L g4621 ( 
.A(n_4596),
.B(n_4448),
.Y(n_4621)
);

OAI21xp33_ASAP7_75t_L g4622 ( 
.A1(n_4540),
.A2(n_4528),
.B(n_4513),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4537),
.B(n_4438),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4583),
.B(n_4495),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_L g4625 ( 
.A(n_4575),
.B(n_4447),
.Y(n_4625)
);

NAND3xp33_ASAP7_75t_L g4626 ( 
.A(n_4550),
.B(n_4554),
.C(n_4579),
.Y(n_4626)
);

OAI21xp5_ASAP7_75t_L g4627 ( 
.A1(n_4595),
.A2(n_4499),
.B(n_4451),
.Y(n_4627)
);

OAI21xp5_ASAP7_75t_SL g4628 ( 
.A1(n_4603),
.A2(n_4323),
.B(n_4427),
.Y(n_4628)
);

OAI21xp5_ASAP7_75t_L g4629 ( 
.A1(n_4571),
.A2(n_4403),
.B(n_4494),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4603),
.B(n_4442),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4588),
.B(n_4557),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4537),
.B(n_4522),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_4588),
.B(n_4449),
.Y(n_4633)
);

NAND3xp33_ASAP7_75t_L g4634 ( 
.A(n_4579),
.B(n_4501),
.C(n_4516),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_4575),
.B(n_4521),
.Y(n_4635)
);

OAI221xp5_ASAP7_75t_L g4636 ( 
.A1(n_4600),
.A2(n_4511),
.B1(n_4486),
.B2(n_4466),
.C(n_4460),
.Y(n_4636)
);

OAI21xp5_ASAP7_75t_SL g4637 ( 
.A1(n_4606),
.A2(n_4417),
.B(n_4459),
.Y(n_4637)
);

NAND3xp33_ASAP7_75t_L g4638 ( 
.A(n_4579),
.B(n_4446),
.C(n_276),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4580),
.B(n_276),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4580),
.B(n_278),
.Y(n_4640)
);

NAND3xp33_ASAP7_75t_L g4641 ( 
.A(n_4579),
.B(n_278),
.C(n_279),
.Y(n_4641)
);

OAI221xp5_ASAP7_75t_SL g4642 ( 
.A1(n_4544),
.A2(n_4585),
.B1(n_4587),
.B2(n_4549),
.C(n_4556),
.Y(n_4642)
);

NAND4xp25_ASAP7_75t_L g4643 ( 
.A(n_4545),
.B(n_279),
.C(n_282),
.D(n_283),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4594),
.B(n_285),
.Y(n_4644)
);

NAND3xp33_ASAP7_75t_L g4645 ( 
.A(n_4579),
.B(n_285),
.C(n_286),
.Y(n_4645)
);

AOI22xp33_ASAP7_75t_L g4646 ( 
.A1(n_4579),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_4646)
);

OAI21xp5_ASAP7_75t_SL g4647 ( 
.A1(n_4606),
.A2(n_290),
.B(n_291),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4594),
.B(n_4584),
.Y(n_4648)
);

AND2x2_ASAP7_75t_L g4649 ( 
.A(n_4557),
.B(n_291),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4594),
.B(n_292),
.Y(n_4650)
);

AND2x2_ASAP7_75t_SL g4651 ( 
.A(n_4544),
.B(n_292),
.Y(n_4651)
);

AOI211xp5_ASAP7_75t_L g4652 ( 
.A1(n_4549),
.A2(n_293),
.B(n_294),
.C(n_295),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4588),
.B(n_295),
.Y(n_4653)
);

NAND3xp33_ASAP7_75t_L g4654 ( 
.A(n_4587),
.B(n_296),
.C(n_297),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4644),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4650),
.Y(n_4656)
);

OAI21xp5_ASAP7_75t_L g4657 ( 
.A1(n_4626),
.A2(n_4574),
.B(n_4601),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4609),
.B(n_4545),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4648),
.Y(n_4659)
);

BUFx6f_ASAP7_75t_L g4660 ( 
.A(n_4653),
.Y(n_4660)
);

AND2x4_ASAP7_75t_SL g4661 ( 
.A(n_4607),
.B(n_4588),
.Y(n_4661)
);

AND2x2_ASAP7_75t_L g4662 ( 
.A(n_4621),
.B(n_4588),
.Y(n_4662)
);

NOR2xp33_ASAP7_75t_L g4663 ( 
.A(n_4613),
.B(n_4588),
.Y(n_4663)
);

BUFx3_ASAP7_75t_L g4664 ( 
.A(n_4649),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4651),
.Y(n_4665)
);

AOI221xp5_ASAP7_75t_L g4666 ( 
.A1(n_4642),
.A2(n_4608),
.B1(n_4628),
.B2(n_4611),
.C(n_4620),
.Y(n_4666)
);

AND2x2_ASAP7_75t_L g4667 ( 
.A(n_4613),
.B(n_4631),
.Y(n_4667)
);

AND2x4_ASAP7_75t_L g4668 ( 
.A(n_4617),
.B(n_4531),
.Y(n_4668)
);

AND2x4_ASAP7_75t_L g4669 ( 
.A(n_4631),
.B(n_4565),
.Y(n_4669)
);

AND2x4_ASAP7_75t_SL g4670 ( 
.A(n_4623),
.B(n_4553),
.Y(n_4670)
);

AND2x4_ASAP7_75t_L g4671 ( 
.A(n_4633),
.B(n_4565),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4630),
.B(n_4591),
.Y(n_4672)
);

AND3x2_ASAP7_75t_L g4673 ( 
.A(n_4652),
.B(n_4584),
.C(n_4563),
.Y(n_4673)
);

OR2x2_ASAP7_75t_L g4674 ( 
.A(n_4618),
.B(n_4551),
.Y(n_4674)
);

AND2x4_ASAP7_75t_L g4675 ( 
.A(n_4633),
.B(n_4565),
.Y(n_4675)
);

AND2x4_ASAP7_75t_L g4676 ( 
.A(n_4630),
.B(n_4565),
.Y(n_4676)
);

INVxp67_ASAP7_75t_SL g4677 ( 
.A(n_4632),
.Y(n_4677)
);

INVx3_ASAP7_75t_L g4678 ( 
.A(n_4651),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4653),
.B(n_4591),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4634),
.Y(n_4680)
);

AO21x2_ASAP7_75t_L g4681 ( 
.A1(n_4629),
.A2(n_4538),
.B(n_4535),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_4647),
.B(n_4594),
.Y(n_4682)
);

HB1xp67_ASAP7_75t_L g4683 ( 
.A(n_4612),
.Y(n_4683)
);

OAI33xp33_ASAP7_75t_L g4684 ( 
.A1(n_4614),
.A2(n_4541),
.A3(n_4555),
.B1(n_4560),
.B2(n_4556),
.B3(n_4559),
.Y(n_4684)
);

INVx1_ASAP7_75t_SL g4685 ( 
.A(n_4658),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4679),
.B(n_4610),
.Y(n_4686)
);

AND2x4_ASAP7_75t_L g4687 ( 
.A(n_4658),
.B(n_4619),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4679),
.Y(n_4688)
);

AND2x2_ASAP7_75t_L g4689 ( 
.A(n_4667),
.B(n_4615),
.Y(n_4689)
);

OR2x2_ASAP7_75t_L g4690 ( 
.A(n_4674),
.B(n_4555),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4660),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_4660),
.B(n_4610),
.Y(n_4692)
);

INVx1_ASAP7_75t_SL g4693 ( 
.A(n_4672),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_4681),
.Y(n_4694)
);

INVxp67_ASAP7_75t_L g4695 ( 
.A(n_4667),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4660),
.B(n_4622),
.Y(n_4696)
);

AND2x2_ASAP7_75t_L g4697 ( 
.A(n_4672),
.B(n_4662),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4681),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4660),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4660),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4664),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4664),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4674),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_L g4704 ( 
.A(n_4678),
.B(n_4569),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4662),
.B(n_4532),
.Y(n_4705)
);

AND2x2_ASAP7_75t_L g4706 ( 
.A(n_4661),
.B(n_4532),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4697),
.Y(n_4707)
);

AND2x2_ASAP7_75t_L g4708 ( 
.A(n_4697),
.B(n_4661),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4693),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4685),
.B(n_4678),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_SL g4711 ( 
.A(n_4690),
.B(n_4666),
.Y(n_4711)
);

OR2x2_ASAP7_75t_L g4712 ( 
.A(n_4690),
.B(n_4683),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4694),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4687),
.B(n_4676),
.Y(n_4714)
);

AND2x2_ASAP7_75t_L g4715 ( 
.A(n_4687),
.B(n_4676),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4688),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4694),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4698),
.Y(n_4718)
);

NAND2xp33_ASAP7_75t_R g4719 ( 
.A(n_4692),
.B(n_4678),
.Y(n_4719)
);

AND2x4_ASAP7_75t_L g4720 ( 
.A(n_4691),
.B(n_4676),
.Y(n_4720)
);

NOR3xp33_ASAP7_75t_L g4721 ( 
.A(n_4698),
.B(n_4684),
.C(n_4682),
.Y(n_4721)
);

NOR2xp33_ASAP7_75t_L g4722 ( 
.A(n_4712),
.B(n_4663),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4714),
.B(n_4687),
.Y(n_4723)
);

NAND2xp5_ASAP7_75t_L g4724 ( 
.A(n_4715),
.B(n_4689),
.Y(n_4724)
);

CKINVDCx20_ASAP7_75t_R g4725 ( 
.A(n_4708),
.Y(n_4725)
);

NAND2xp33_ASAP7_75t_SL g4726 ( 
.A(n_4707),
.B(n_4689),
.Y(n_4726)
);

INVxp67_ASAP7_75t_SL g4727 ( 
.A(n_4711),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4710),
.Y(n_4728)
);

OAI22xp33_ASAP7_75t_L g4729 ( 
.A1(n_4711),
.A2(n_4636),
.B1(n_4638),
.B2(n_4620),
.Y(n_4729)
);

AOI22xp5_ASAP7_75t_L g4730 ( 
.A1(n_4721),
.A2(n_4681),
.B1(n_4680),
.B2(n_4665),
.Y(n_4730)
);

AND2x2_ASAP7_75t_SL g4731 ( 
.A(n_4730),
.B(n_4721),
.Y(n_4731)
);

NAND3xp33_ASAP7_75t_L g4732 ( 
.A(n_4727),
.B(n_4719),
.C(n_4718),
.Y(n_4732)
);

INVx2_ASAP7_75t_L g4733 ( 
.A(n_4725),
.Y(n_4733)
);

AOI21xp33_ASAP7_75t_SL g4734 ( 
.A1(n_4722),
.A2(n_4724),
.B(n_4686),
.Y(n_4734)
);

AND2x2_ASAP7_75t_L g4735 ( 
.A(n_4723),
.B(n_4676),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4726),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4728),
.Y(n_4737)
);

OAI31xp33_ASAP7_75t_L g4738 ( 
.A1(n_4729),
.A2(n_4680),
.A3(n_4659),
.B(n_4656),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4727),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4727),
.Y(n_4740)
);

OR2x2_ASAP7_75t_L g4741 ( 
.A(n_4727),
.B(n_4695),
.Y(n_4741)
);

INVx2_ASAP7_75t_L g4742 ( 
.A(n_4725),
.Y(n_4742)
);

NOR2xp33_ASAP7_75t_L g4743 ( 
.A(n_4733),
.B(n_4665),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4742),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4741),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4739),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4740),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4732),
.Y(n_4748)
);

NOR2xp33_ASAP7_75t_L g4749 ( 
.A(n_4734),
.B(n_4670),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4735),
.B(n_4677),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4731),
.B(n_4699),
.Y(n_4751)
);

OR2x2_ASAP7_75t_L g4752 ( 
.A(n_4750),
.B(n_4701),
.Y(n_4752)
);

AOI221xp5_ASAP7_75t_L g4753 ( 
.A1(n_4748),
.A2(n_4732),
.B1(n_4659),
.B2(n_4738),
.C(n_4657),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4751),
.Y(n_4754)
);

INVx2_ASAP7_75t_L g4755 ( 
.A(n_4745),
.Y(n_4755)
);

NOR2xp33_ASAP7_75t_L g4756 ( 
.A(n_4744),
.B(n_4670),
.Y(n_4756)
);

NOR2x1_ASAP7_75t_L g4757 ( 
.A(n_4749),
.B(n_4736),
.Y(n_4757)
);

OAI322xp33_ASAP7_75t_L g4758 ( 
.A1(n_4743),
.A2(n_4731),
.A3(n_4719),
.B1(n_4703),
.B2(n_4696),
.C1(n_4700),
.C2(n_4704),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4746),
.B(n_4720),
.Y(n_4759)
);

OAI21xp5_ASAP7_75t_SL g4760 ( 
.A1(n_4753),
.A2(n_4738),
.B(n_4747),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4756),
.B(n_4720),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4755),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4759),
.Y(n_4763)
);

INVx2_ASAP7_75t_L g4764 ( 
.A(n_4752),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4758),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4757),
.B(n_4702),
.Y(n_4766)
);

XNOR2xp5_ASAP7_75t_L g4767 ( 
.A(n_4766),
.B(n_4709),
.Y(n_4767)
);

OR2x2_ASAP7_75t_L g4768 ( 
.A(n_4764),
.B(n_4705),
.Y(n_4768)
);

XOR2xp5_ASAP7_75t_L g4769 ( 
.A(n_4761),
.B(n_4754),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4762),
.B(n_4705),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4763),
.Y(n_4771)
);

AND2x2_ASAP7_75t_L g4772 ( 
.A(n_4765),
.B(n_4668),
.Y(n_4772)
);

NAND4xp25_ASAP7_75t_SL g4773 ( 
.A(n_4760),
.B(n_4716),
.C(n_4737),
.D(n_4706),
.Y(n_4773)
);

OAI31xp33_ASAP7_75t_L g4774 ( 
.A1(n_4760),
.A2(n_4655),
.A3(n_4656),
.B(n_4713),
.Y(n_4774)
);

AOI22xp5_ASAP7_75t_L g4775 ( 
.A1(n_4762),
.A2(n_4655),
.B1(n_4675),
.B2(n_4671),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4766),
.B(n_4706),
.Y(n_4776)
);

OAI22xp5_ASAP7_75t_L g4777 ( 
.A1(n_4764),
.A2(n_4675),
.B1(n_4671),
.B2(n_4669),
.Y(n_4777)
);

AOI222xp33_ASAP7_75t_L g4778 ( 
.A1(n_4760),
.A2(n_4717),
.B1(n_4713),
.B2(n_4675),
.C1(n_4671),
.C2(n_4535),
.Y(n_4778)
);

AND2x2_ASAP7_75t_L g4779 ( 
.A(n_4766),
.B(n_4668),
.Y(n_4779)
);

OAI21xp5_ASAP7_75t_SL g4780 ( 
.A1(n_4760),
.A2(n_4675),
.B(n_4671),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4768),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4769),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4767),
.Y(n_4783)
);

HB1xp67_ASAP7_75t_L g4784 ( 
.A(n_4779),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4776),
.Y(n_4785)
);

BUFx2_ASAP7_75t_L g4786 ( 
.A(n_4770),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4775),
.Y(n_4787)
);

INVxp33_ASAP7_75t_SL g4788 ( 
.A(n_4772),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4778),
.Y(n_4789)
);

BUFx6f_ASAP7_75t_L g4790 ( 
.A(n_4771),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4777),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4780),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4773),
.Y(n_4793)
);

INVx2_ASAP7_75t_L g4794 ( 
.A(n_4774),
.Y(n_4794)
);

INVx2_ASAP7_75t_L g4795 ( 
.A(n_4768),
.Y(n_4795)
);

INVx5_ASAP7_75t_SL g4796 ( 
.A(n_4769),
.Y(n_4796)
);

HB1xp67_ASAP7_75t_L g4797 ( 
.A(n_4779),
.Y(n_4797)
);

CKINVDCx20_ASAP7_75t_R g4798 ( 
.A(n_4769),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4768),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4768),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4778),
.B(n_4625),
.Y(n_4801)
);

INVxp67_ASAP7_75t_L g4802 ( 
.A(n_4779),
.Y(n_4802)
);

INVxp67_ASAP7_75t_L g4803 ( 
.A(n_4779),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4768),
.Y(n_4804)
);

INVx1_ASAP7_75t_SL g4805 ( 
.A(n_4779),
.Y(n_4805)
);

OAI211xp5_ASAP7_75t_L g4806 ( 
.A1(n_4802),
.A2(n_4717),
.B(n_4639),
.C(n_4640),
.Y(n_4806)
);

O2A1O1Ixp5_ASAP7_75t_L g4807 ( 
.A1(n_4795),
.A2(n_4669),
.B(n_4668),
.C(n_4535),
.Y(n_4807)
);

NOR2xp33_ASAP7_75t_L g4808 ( 
.A(n_4798),
.B(n_4788),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4784),
.Y(n_4809)
);

NAND4xp25_ASAP7_75t_SL g4810 ( 
.A(n_4792),
.B(n_4616),
.C(n_4624),
.D(n_4646),
.Y(n_4810)
);

AND2x2_ASAP7_75t_L g4811 ( 
.A(n_4797),
.B(n_4669),
.Y(n_4811)
);

AOI211x1_ASAP7_75t_SL g4812 ( 
.A1(n_4801),
.A2(n_4593),
.B(n_4590),
.C(n_4538),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4790),
.Y(n_4813)
);

OAI211xp5_ASAP7_75t_SL g4814 ( 
.A1(n_4803),
.A2(n_4646),
.B(n_4635),
.C(n_4637),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4790),
.Y(n_4815)
);

OAI22xp5_ASAP7_75t_L g4816 ( 
.A1(n_4781),
.A2(n_4800),
.B1(n_4804),
.B2(n_4799),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4796),
.Y(n_4817)
);

OAI21xp5_ASAP7_75t_L g4818 ( 
.A1(n_4789),
.A2(n_4669),
.B(n_4538),
.Y(n_4818)
);

INVx1_ASAP7_75t_SL g4819 ( 
.A(n_4805),
.Y(n_4819)
);

OAI22xp33_ASAP7_75t_L g4820 ( 
.A1(n_4790),
.A2(n_4560),
.B1(n_4593),
.B2(n_4590),
.Y(n_4820)
);

INVx2_ASAP7_75t_L g4821 ( 
.A(n_4796),
.Y(n_4821)
);

OAI22xp5_ASAP7_75t_L g4822 ( 
.A1(n_4786),
.A2(n_4564),
.B1(n_4562),
.B2(n_4569),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4782),
.Y(n_4823)
);

OAI22xp5_ASAP7_75t_L g4824 ( 
.A1(n_4785),
.A2(n_4564),
.B1(n_4562),
.B2(n_4563),
.Y(n_4824)
);

INVxp67_ASAP7_75t_L g4825 ( 
.A(n_4787),
.Y(n_4825)
);

AOI221xp5_ASAP7_75t_L g4826 ( 
.A1(n_4794),
.A2(n_4590),
.B1(n_4593),
.B2(n_4654),
.C(n_4641),
.Y(n_4826)
);

OAI22xp5_ASAP7_75t_L g4827 ( 
.A1(n_4783),
.A2(n_4791),
.B1(n_4793),
.B2(n_4561),
.Y(n_4827)
);

CKINVDCx20_ASAP7_75t_R g4828 ( 
.A(n_4798),
.Y(n_4828)
);

OAI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_4784),
.A2(n_4563),
.B(n_4561),
.Y(n_4829)
);

NAND4xp25_ASAP7_75t_L g4830 ( 
.A(n_4805),
.B(n_4561),
.C(n_4643),
.D(n_4533),
.Y(n_4830)
);

INVx1_ASAP7_75t_SL g4831 ( 
.A(n_4798),
.Y(n_4831)
);

NAND2xp5_ASAP7_75t_L g4832 ( 
.A(n_4796),
.B(n_4673),
.Y(n_4832)
);

OAI221xp5_ASAP7_75t_L g4833 ( 
.A1(n_4802),
.A2(n_4645),
.B1(n_4627),
.B2(n_4552),
.C(n_4533),
.Y(n_4833)
);

AOI22xp5_ASAP7_75t_L g4834 ( 
.A1(n_4828),
.A2(n_4570),
.B1(n_4552),
.B2(n_4576),
.Y(n_4834)
);

OAI221xp5_ASAP7_75t_L g4835 ( 
.A1(n_4831),
.A2(n_4533),
.B1(n_4552),
.B2(n_4585),
.C(n_4582),
.Y(n_4835)
);

OAI211xp5_ASAP7_75t_L g4836 ( 
.A1(n_4819),
.A2(n_4582),
.B(n_4577),
.C(n_4546),
.Y(n_4836)
);

AOI221xp5_ASAP7_75t_L g4837 ( 
.A1(n_4808),
.A2(n_4570),
.B1(n_4576),
.B2(n_4577),
.C(n_4582),
.Y(n_4837)
);

AOI211xp5_ASAP7_75t_L g4838 ( 
.A1(n_4816),
.A2(n_4577),
.B(n_4604),
.C(n_4602),
.Y(n_4838)
);

AOI221xp5_ASAP7_75t_L g4839 ( 
.A1(n_4817),
.A2(n_4821),
.B1(n_4809),
.B2(n_4818),
.C(n_4827),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4811),
.B(n_4604),
.Y(n_4840)
);

NAND4xp25_ASAP7_75t_L g4841 ( 
.A(n_4832),
.B(n_4604),
.C(n_4602),
.D(n_4598),
.Y(n_4841)
);

AOI221xp5_ASAP7_75t_SL g4842 ( 
.A1(n_4813),
.A2(n_4534),
.B1(n_4546),
.B2(n_4547),
.C(n_4559),
.Y(n_4842)
);

AOI211xp5_ASAP7_75t_L g4843 ( 
.A1(n_4815),
.A2(n_4823),
.B(n_4806),
.C(n_4822),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4807),
.Y(n_4844)
);

OAI211xp5_ASAP7_75t_SL g4845 ( 
.A1(n_4812),
.A2(n_4586),
.B(n_4589),
.C(n_4598),
.Y(n_4845)
);

NAND2xp5_ASAP7_75t_L g4846 ( 
.A(n_4829),
.B(n_4820),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4825),
.Y(n_4847)
);

OR2x2_ASAP7_75t_L g4848 ( 
.A(n_4830),
.B(n_4598),
.Y(n_4848)
);

AOI221x1_ASAP7_75t_L g4849 ( 
.A1(n_4814),
.A2(n_4824),
.B1(n_4810),
.B2(n_4833),
.C(n_4826),
.Y(n_4849)
);

NAND3xp33_ASAP7_75t_SL g4850 ( 
.A(n_4828),
.B(n_4602),
.C(n_4589),
.Y(n_4850)
);

AOI21xp5_ASAP7_75t_L g4851 ( 
.A1(n_4831),
.A2(n_4547),
.B(n_4534),
.Y(n_4851)
);

OAI222xp33_ASAP7_75t_L g4852 ( 
.A1(n_4831),
.A2(n_4558),
.B1(n_4592),
.B2(n_4548),
.C1(n_4543),
.C2(n_4567),
.Y(n_4852)
);

AOI211x1_ASAP7_75t_SL g4853 ( 
.A1(n_4818),
.A2(n_4567),
.B(n_4543),
.C(n_4548),
.Y(n_4853)
);

AOI221x1_ASAP7_75t_L g4854 ( 
.A1(n_4827),
.A2(n_4573),
.B1(n_4542),
.B2(n_4578),
.C(n_4592),
.Y(n_4854)
);

AOI322xp5_ASAP7_75t_L g4855 ( 
.A1(n_4828),
.A2(n_4567),
.A3(n_4578),
.B1(n_4573),
.B2(n_4542),
.C1(n_4558),
.C2(n_4568),
.Y(n_4855)
);

OAI211xp5_ASAP7_75t_L g4856 ( 
.A1(n_4831),
.A2(n_297),
.B(n_299),
.C(n_300),
.Y(n_4856)
);

NOR2x1p5_ASAP7_75t_L g4857 ( 
.A(n_4809),
.B(n_300),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_4828),
.B(n_4568),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4858),
.Y(n_4859)
);

A2O1A1Ixp33_ASAP7_75t_L g4860 ( 
.A1(n_4844),
.A2(n_4568),
.B(n_303),
.C(n_304),
.Y(n_4860)
);

AOI211xp5_ASAP7_75t_L g4861 ( 
.A1(n_4839),
.A2(n_301),
.B(n_303),
.C(n_306),
.Y(n_4861)
);

AOI221xp5_ASAP7_75t_L g4862 ( 
.A1(n_4835),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.C(n_310),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4840),
.Y(n_4863)
);

AND4x2_ASAP7_75t_L g4864 ( 
.A(n_4851),
.B(n_4837),
.C(n_4843),
.D(n_4849),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4853),
.Y(n_4865)
);

AOI222xp33_ASAP7_75t_L g4866 ( 
.A1(n_4850),
.A2(n_4847),
.B1(n_4852),
.B2(n_4845),
.C1(n_4836),
.C2(n_4846),
.Y(n_4866)
);

AO22x2_ASAP7_75t_L g4867 ( 
.A1(n_4856),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_4867)
);

AOI221xp5_ASAP7_75t_SL g4868 ( 
.A1(n_4841),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.C(n_315),
.Y(n_4868)
);

OAI22xp5_ASAP7_75t_L g4869 ( 
.A1(n_4834),
.A2(n_312),
.B1(n_313),
.B2(n_317),
.Y(n_4869)
);

AOI22xp5_ASAP7_75t_L g4870 ( 
.A1(n_4848),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_4870)
);

OAI221xp5_ASAP7_75t_L g4871 ( 
.A1(n_4842),
.A2(n_318),
.B1(n_319),
.B2(n_321),
.C(n_322),
.Y(n_4871)
);

NOR2x1_ASAP7_75t_L g4872 ( 
.A(n_4857),
.B(n_4854),
.Y(n_4872)
);

AOI222xp33_ASAP7_75t_L g4873 ( 
.A1(n_4838),
.A2(n_321),
.B1(n_322),
.B2(n_325),
.C1(n_326),
.C2(n_327),
.Y(n_4873)
);

NOR4xp25_ASAP7_75t_L g4874 ( 
.A(n_4855),
.B(n_326),
.C(n_328),
.D(n_329),
.Y(n_4874)
);

BUFx3_ASAP7_75t_L g4875 ( 
.A(n_4847),
.Y(n_4875)
);

OA22x2_ASAP7_75t_L g4876 ( 
.A1(n_4844),
.A2(n_328),
.B1(n_331),
.B2(n_332),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4872),
.Y(n_4877)
);

NOR2xp67_ASAP7_75t_L g4878 ( 
.A(n_4871),
.B(n_331),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4860),
.Y(n_4879)
);

AND2x2_ASAP7_75t_SL g4880 ( 
.A(n_4874),
.B(n_4863),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_SL g4881 ( 
.A(n_4866),
.B(n_333),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_4875),
.B(n_333),
.Y(n_4882)
);

INVxp67_ASAP7_75t_L g4883 ( 
.A(n_4865),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4867),
.Y(n_4884)
);

AOI22xp5_ASAP7_75t_L g4885 ( 
.A1(n_4859),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4876),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4864),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4867),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4870),
.Y(n_4889)
);

AOI22xp5_ASAP7_75t_L g4890 ( 
.A1(n_4868),
.A2(n_334),
.B1(n_336),
.B2(n_338),
.Y(n_4890)
);

AND2x2_ASAP7_75t_L g4891 ( 
.A(n_4873),
.B(n_338),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4877),
.Y(n_4892)
);

NAND4xp75_ASAP7_75t_L g4893 ( 
.A(n_4887),
.B(n_4862),
.C(n_4861),
.D(n_4869),
.Y(n_4893)
);

AND2x2_ASAP7_75t_SL g4894 ( 
.A(n_4880),
.B(n_339),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_SL g4895 ( 
.A(n_4884),
.B(n_340),
.Y(n_4895)
);

NAND2xp5_ASAP7_75t_L g4896 ( 
.A(n_4888),
.B(n_341),
.Y(n_4896)
);

NAND2x1p5_ASAP7_75t_L g4897 ( 
.A(n_4886),
.B(n_342),
.Y(n_4897)
);

INVx2_ASAP7_75t_L g4898 ( 
.A(n_4891),
.Y(n_4898)
);

BUFx6f_ASAP7_75t_L g4899 ( 
.A(n_4881),
.Y(n_4899)
);

NOR2x1p5_ASAP7_75t_L g4900 ( 
.A(n_4879),
.B(n_342),
.Y(n_4900)
);

AOI22xp33_ASAP7_75t_L g4901 ( 
.A1(n_4883),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_4901)
);

NOR2x1_ASAP7_75t_L g4902 ( 
.A(n_4882),
.B(n_344),
.Y(n_4902)
);

AOI22xp33_ASAP7_75t_L g4903 ( 
.A1(n_4889),
.A2(n_4878),
.B1(n_4890),
.B2(n_4885),
.Y(n_4903)
);

AND2x4_ASAP7_75t_L g4904 ( 
.A(n_4877),
.B(n_346),
.Y(n_4904)
);

HB1xp67_ASAP7_75t_L g4905 ( 
.A(n_4887),
.Y(n_4905)
);

NAND2xp33_ASAP7_75t_SL g4906 ( 
.A(n_4892),
.B(n_346),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_SL g4907 ( 
.A(n_4894),
.B(n_347),
.Y(n_4907)
);

NOR2xp33_ASAP7_75t_R g4908 ( 
.A(n_4896),
.B(n_4905),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4898),
.B(n_349),
.Y(n_4909)
);

NOR3xp33_ASAP7_75t_SL g4910 ( 
.A(n_4895),
.B(n_350),
.C(n_351),
.Y(n_4910)
);

NOR2xp33_ASAP7_75t_R g4911 ( 
.A(n_4899),
.B(n_351),
.Y(n_4911)
);

NOR2xp33_ASAP7_75t_R g4912 ( 
.A(n_4899),
.B(n_353),
.Y(n_4912)
);

NOR2xp33_ASAP7_75t_R g4913 ( 
.A(n_4904),
.B(n_4903),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_SL g4914 ( 
.A(n_4897),
.B(n_354),
.Y(n_4914)
);

NOR2xp33_ASAP7_75t_R g4915 ( 
.A(n_4901),
.B(n_355),
.Y(n_4915)
);

AOI221xp5_ASAP7_75t_L g4916 ( 
.A1(n_4906),
.A2(n_4900),
.B1(n_4902),
.B2(n_4893),
.C(n_358),
.Y(n_4916)
);

NOR2x1p5_ASAP7_75t_L g4917 ( 
.A(n_4909),
.B(n_355),
.Y(n_4917)
);

INVx2_ASAP7_75t_L g4918 ( 
.A(n_4907),
.Y(n_4918)
);

NAND3xp33_ASAP7_75t_L g4919 ( 
.A(n_4914),
.B(n_356),
.C(n_357),
.Y(n_4919)
);

OAI221xp5_ASAP7_75t_L g4920 ( 
.A1(n_4910),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.C(n_359),
.Y(n_4920)
);

CKINVDCx20_ASAP7_75t_R g4921 ( 
.A(n_4913),
.Y(n_4921)
);

NOR3xp33_ASAP7_75t_L g4922 ( 
.A(n_4908),
.B(n_361),
.C(n_362),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4921),
.B(n_4911),
.Y(n_4923)
);

NOR3xp33_ASAP7_75t_L g4924 ( 
.A(n_4916),
.B(n_4912),
.C(n_4915),
.Y(n_4924)
);

NAND3x1_ASAP7_75t_L g4925 ( 
.A(n_4922),
.B(n_361),
.C(n_362),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4923),
.Y(n_4926)
);

AOI22xp33_ASAP7_75t_L g4927 ( 
.A1(n_4924),
.A2(n_4918),
.B1(n_4917),
.B2(n_4919),
.Y(n_4927)
);

OAI22xp5_ASAP7_75t_SL g4928 ( 
.A1(n_4927),
.A2(n_4920),
.B1(n_4925),
.B2(n_365),
.Y(n_4928)
);

AOI22xp5_ASAP7_75t_L g4929 ( 
.A1(n_4926),
.A2(n_363),
.B1(n_364),
.B2(n_366),
.Y(n_4929)
);

INVx2_ASAP7_75t_L g4930 ( 
.A(n_4928),
.Y(n_4930)
);

OR3x1_ASAP7_75t_L g4931 ( 
.A(n_4929),
.B(n_363),
.C(n_367),
.Y(n_4931)
);

BUFx2_ASAP7_75t_SL g4932 ( 
.A(n_4929),
.Y(n_4932)
);

AOI31xp33_ASAP7_75t_L g4933 ( 
.A1(n_4930),
.A2(n_4932),
.A3(n_4931),
.B(n_369),
.Y(n_4933)
);

AOI31xp33_ASAP7_75t_L g4934 ( 
.A1(n_4930),
.A2(n_367),
.A3(n_368),
.B(n_371),
.Y(n_4934)
);

AOI22xp33_ASAP7_75t_L g4935 ( 
.A1(n_4930),
.A2(n_368),
.B1(n_374),
.B2(n_375),
.Y(n_4935)
);

AOI22xp33_ASAP7_75t_L g4936 ( 
.A1(n_4930),
.A2(n_374),
.B1(n_375),
.B2(n_376),
.Y(n_4936)
);

AOI22xp5_ASAP7_75t_L g4937 ( 
.A1(n_4935),
.A2(n_376),
.B1(n_377),
.B2(n_378),
.Y(n_4937)
);

AOI22xp5_ASAP7_75t_L g4938 ( 
.A1(n_4936),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4933),
.Y(n_4939)
);

INVx3_ASAP7_75t_L g4940 ( 
.A(n_4934),
.Y(n_4940)
);

AOI22xp5_ASAP7_75t_L g4941 ( 
.A1(n_4935),
.A2(n_379),
.B1(n_382),
.B2(n_383),
.Y(n_4941)
);

AO21x2_ASAP7_75t_L g4942 ( 
.A1(n_4939),
.A2(n_384),
.B(n_385),
.Y(n_4942)
);

NAND2x1p5_ASAP7_75t_L g4943 ( 
.A(n_4940),
.B(n_384),
.Y(n_4943)
);

INVx1_ASAP7_75t_SL g4944 ( 
.A(n_4941),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_L g4945 ( 
.A(n_4937),
.B(n_385),
.Y(n_4945)
);

AOI22xp33_ASAP7_75t_L g4946 ( 
.A1(n_4938),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4940),
.Y(n_4947)
);

NAND2xp5_ASAP7_75t_L g4948 ( 
.A(n_4939),
.B(n_387),
.Y(n_4948)
);

OAI221xp5_ASAP7_75t_SL g4949 ( 
.A1(n_4939),
.A2(n_390),
.B1(n_392),
.B2(n_393),
.C(n_394),
.Y(n_4949)
);

AND2x2_ASAP7_75t_L g4950 ( 
.A(n_4939),
.B(n_395),
.Y(n_4950)
);

AOI21xp5_ASAP7_75t_L g4951 ( 
.A1(n_4939),
.A2(n_395),
.B(n_396),
.Y(n_4951)
);

INVxp67_ASAP7_75t_SL g4952 ( 
.A(n_4939),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4952),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4947),
.Y(n_4954)
);

XNOR2x1_ASAP7_75t_L g4955 ( 
.A(n_4944),
.B(n_396),
.Y(n_4955)
);

AOI22xp33_ASAP7_75t_SL g4956 ( 
.A1(n_4943),
.A2(n_397),
.B1(n_398),
.B2(n_401),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4945),
.Y(n_4957)
);

AO21x2_ASAP7_75t_L g4958 ( 
.A1(n_4951),
.A2(n_397),
.B(n_401),
.Y(n_4958)
);

AOI22xp33_ASAP7_75t_SL g4959 ( 
.A1(n_4950),
.A2(n_402),
.B1(n_403),
.B2(n_404),
.Y(n_4959)
);

INVx2_ASAP7_75t_SL g4960 ( 
.A(n_4942),
.Y(n_4960)
);

AOI222xp33_ASAP7_75t_L g4961 ( 
.A1(n_4946),
.A2(n_403),
.B1(n_405),
.B2(n_406),
.C1(n_407),
.C2(n_409),
.Y(n_4961)
);

XOR2xp5_ASAP7_75t_L g4962 ( 
.A(n_4953),
.B(n_4954),
.Y(n_4962)
);

AOI21xp33_ASAP7_75t_SL g4963 ( 
.A1(n_4960),
.A2(n_4948),
.B(n_4949),
.Y(n_4963)
);

XNOR2xp5_ASAP7_75t_L g4964 ( 
.A(n_4957),
.B(n_4955),
.Y(n_4964)
);

INVxp67_ASAP7_75t_L g4965 ( 
.A(n_4958),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4956),
.Y(n_4966)
);

AOI322xp5_ASAP7_75t_L g4967 ( 
.A1(n_4965),
.A2(n_4959),
.A3(n_4961),
.B1(n_409),
.B2(n_410),
.C1(n_412),
.C2(n_414),
.Y(n_4967)
);

AOI22xp5_ASAP7_75t_L g4968 ( 
.A1(n_4962),
.A2(n_4964),
.B1(n_4966),
.B2(n_4963),
.Y(n_4968)
);

AOI322xp5_ASAP7_75t_L g4969 ( 
.A1(n_4965),
.A2(n_406),
.A3(n_407),
.B1(n_410),
.B2(n_415),
.C1(n_416),
.C2(n_417),
.Y(n_4969)
);

BUFx4_ASAP7_75t_R g4970 ( 
.A(n_4962),
.Y(n_4970)
);

OAI221xp5_ASAP7_75t_R g4971 ( 
.A1(n_4968),
.A2(n_415),
.B1(n_416),
.B2(n_418),
.C(n_420),
.Y(n_4971)
);

AOI221xp5_ASAP7_75t_L g4972 ( 
.A1(n_4970),
.A2(n_424),
.B1(n_425),
.B2(n_427),
.C(n_428),
.Y(n_4972)
);

AOI22xp33_ASAP7_75t_L g4973 ( 
.A1(n_4972),
.A2(n_4967),
.B1(n_4969),
.B2(n_447),
.Y(n_4973)
);

AOI211xp5_ASAP7_75t_L g4974 ( 
.A1(n_4973),
.A2(n_4971),
.B(n_445),
.C(n_448),
.Y(n_4974)
);


endmodule