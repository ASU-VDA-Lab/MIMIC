module real_jpeg_29799_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_4),
.B1(n_25),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_29),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_20),
.B1(n_23),
.B2(n_29),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_3),
.A2(n_20),
.B(n_22),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_3),
.A2(n_29),
.B1(n_45),
.B2(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_19),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_9),
.B(n_38),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_42),
.B(n_46),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_3),
.B(n_51),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_4),
.A2(n_7),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_4),
.A2(n_21),
.B(n_29),
.C(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_5),
.Y(n_105)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_6),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_7),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_7),
.A2(n_26),
.B1(n_45),
.B2(n_46),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_9),
.A2(n_20),
.B1(n_23),
.B2(n_52),
.Y(n_57)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_10),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_109),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_107),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_83),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_15),
.B(n_83),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_60),
.C(n_73),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_16),
.B(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_32),
.B1(n_58),
.B2(n_59),
.Y(n_16)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_17),
.B(n_33),
.C(n_49),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_24),
.B(n_27),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_19),
.A2(n_28),
.B1(n_30),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

INVx5_ASAP7_75t_SL g23 ( 
.A(n_20),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_20),
.A2(n_29),
.B(n_115),
.C(n_116),
.Y(n_114)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_29),
.A2(n_38),
.B(n_43),
.C(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_29),
.B(n_70),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_29),
.B(n_44),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_36),
.B(n_40),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_36),
.A2(n_40),
.B1(n_44),
.B2(n_99),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_45),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_67),
.Y(n_66)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_97),
.C(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_48),
.A2(n_49),
.B1(n_96),
.B2(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_54),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_53),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_60),
.A2(n_61),
.B1(n_73),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_71),
.B2(n_72),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_71),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_64),
.A2(n_72),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_64),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_64),
.B(n_153),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_64),
.B(n_130),
.C(n_142),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_67),
.B(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_66),
.B(n_67),
.Y(n_119)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_73),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.C(n_81),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_74),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_89),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_81),
.B1(n_82),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_77),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_104),
.B(n_106),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_96),
.A2(n_97),
.B1(n_137),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_97),
.B(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_101),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_163),
.B(n_168),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_133),
.B(n_162),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_121),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_112),
.B(n_121),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_120),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_127),
.B2(n_128),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_130),
.C(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_129),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_132),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_157),
.B(n_161),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_144),
.B(n_156),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_139),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_137),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_140),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_141),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_148),
.B(n_155),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.B(n_154),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.Y(n_168)
);


endmodule