module fake_jpeg_18202_n_114 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx4f_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_15),
.B1(n_17),
.B2(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_10),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_13),
.Y(n_40)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_23),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_12),
.B(n_9),
.Y(n_47)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_20),
.C(n_10),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_19),
.B1(n_30),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_12),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_46),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_22),
.B(n_10),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_43),
.C(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_53),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_38),
.B1(n_43),
.B2(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_27),
.B(n_20),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_22),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_32),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_36),
.C(n_16),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_36),
.B1(n_41),
.B2(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_63),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_11),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_70),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_72),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_59),
.C(n_1),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_16),
.B(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_75),
.Y(n_81)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_42),
.B(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_80),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_57),
.C(n_62),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_82),
.C(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_91),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_96),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_76),
.B(n_72),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_82),
.B1(n_77),
.B2(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_93),
.C(n_92),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.C(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_54),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_0),
.B(n_1),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_3),
.B(n_4),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_11),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_2),
.C2(n_7),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_106),
.B(n_3),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_2),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_107),
.B(n_104),
.CI(n_6),
.CON(n_110),
.SN(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_110),
.A2(n_6),
.B(n_8),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_112),
.B(n_110),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_111),
.Y(n_114)
);


endmodule