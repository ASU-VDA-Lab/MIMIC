module fake_jpeg_11284_n_544 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_544);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_544;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_19),
.B(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_67),
.B(n_72),
.Y(n_152)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_74),
.Y(n_177)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_15),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_76),
.B(n_95),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_78),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_32),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g184 ( 
.A(n_87),
.Y(n_184)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_88),
.Y(n_151)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_90),
.Y(n_192)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_19),
.B(n_0),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_99),
.B(n_112),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_18),
.Y(n_109)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_18),
.Y(n_110)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_43),
.B(n_12),
.Y(n_112)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_25),
.Y(n_114)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_35),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_1),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_37),
.Y(n_161)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_119),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_33),
.Y(n_120)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_42),
.Y(n_122)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_45),
.B1(n_56),
.B2(n_47),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_124),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_126),
.A2(n_3),
.B(n_5),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_35),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_127),
.B(n_129),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_50),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_131),
.B(n_140),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_34),
.B1(n_49),
.B2(n_51),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_137),
.A2(n_157),
.B1(n_176),
.B2(n_190),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_67),
.B(n_50),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_139),
.B(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_99),
.B(n_31),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_103),
.A2(n_34),
.B1(n_46),
.B2(n_37),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_144),
.B(n_98),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_104),
.A2(n_34),
.B1(n_51),
.B2(n_46),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_161),
.B(n_180),
.Y(n_264)
);

INVx6_ASAP7_75t_SL g165 ( 
.A(n_74),
.Y(n_165)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_109),
.A2(n_26),
.B1(n_37),
.B2(n_51),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_64),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_178),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_88),
.B(n_56),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_87),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_24),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_119),
.A2(n_46),
.B1(n_37),
.B2(n_53),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_110),
.A2(n_53),
.B1(n_47),
.B2(n_58),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_200),
.A2(n_157),
.B1(n_137),
.B2(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_201),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_173),
.A2(n_38),
.B1(n_58),
.B2(n_54),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_202),
.Y(n_269)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_203),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_175),
.A2(n_38),
.B1(n_54),
.B2(n_48),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_205),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_156),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_206),
.B(n_222),
.Y(n_272)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_208),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_152),
.B(n_31),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_210),
.B(n_219),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_211),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_200),
.A2(n_36),
.B(n_48),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_212),
.B(n_225),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_97),
.B1(n_90),
.B2(n_86),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_85),
.B1(n_83),
.B2(n_79),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_138),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_215),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_145),
.A2(n_20),
.B1(n_36),
.B2(n_30),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_218),
.A2(n_220),
.B1(n_231),
.B2(n_267),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_152),
.B(n_20),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_146),
.A2(n_30),
.B1(n_24),
.B2(n_23),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_135),
.B(n_23),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_223),
.B(n_226),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_167),
.B(n_3),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_224),
.B(n_158),
.C(n_159),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_176),
.A2(n_78),
.B1(n_77),
.B2(n_71),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_227),
.A2(n_240),
.B1(n_251),
.B2(n_257),
.Y(n_307)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_228),
.Y(n_291)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_161),
.A2(n_65),
.B1(n_7),
.B2(n_8),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_230),
.A2(n_143),
.B(n_187),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_167),
.B(n_7),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_232),
.B(n_234),
.Y(n_283)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_133),
.Y(n_233)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_233),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_199),
.B(n_8),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_196),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_236),
.B(n_248),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_141),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_237),
.B(n_243),
.Y(n_284)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_148),
.Y(n_238)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_190),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_199),
.B(n_9),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_255),
.Y(n_270)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_242),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_141),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_177),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_245),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_171),
.B(n_9),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_151),
.B(n_11),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_249),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_147),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_136),
.B(n_11),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_151),
.B(n_128),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_160),
.Y(n_250)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_168),
.B(n_150),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_181),
.Y(n_256)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_192),
.A2(n_183),
.B1(n_134),
.B2(n_166),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_154),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_259),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_125),
.B(n_130),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_155),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_266),
.Y(n_276)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_262),
.Y(n_311)
);

AOI22x1_ASAP7_75t_L g299 ( 
.A1(n_264),
.A2(n_230),
.B1(n_216),
.B2(n_227),
.Y(n_299)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_265),
.Y(n_312)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_132),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_153),
.A2(n_138),
.B1(n_194),
.B2(n_174),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_255),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_273),
.B(n_275),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_262),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_209),
.A2(n_142),
.B1(n_169),
.B2(n_158),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_279),
.A2(n_314),
.B1(n_246),
.B2(n_249),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_217),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_310),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_286),
.A2(n_235),
.B(n_237),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_293),
.B(n_297),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_224),
.B(n_159),
.C(n_169),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_295),
.B(n_300),
.C(n_316),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_210),
.B(n_174),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_194),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_305),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_299),
.A2(n_250),
.B(n_242),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_229),
.C(n_264),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_219),
.B(n_204),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_301),
.B(n_236),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_248),
.B(n_241),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_217),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_234),
.A2(n_231),
.B1(n_232),
.B2(n_221),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_201),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_279),
.A2(n_258),
.B1(n_235),
.B2(n_206),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_322),
.A2(n_341),
.B1(n_347),
.B2(n_360),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_323),
.B(n_346),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_276),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_327),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_300),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_329),
.C(n_289),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_276),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_271),
.Y(n_328)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_270),
.B(n_239),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_269),
.A2(n_226),
.B(n_208),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_330),
.A2(n_349),
.B(n_350),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_331),
.A2(n_352),
.B(n_355),
.Y(n_367)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_268),
.Y(n_332)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_332),
.Y(n_391)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_294),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_334),
.B(n_338),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_284),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_278),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_337),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_277),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_339),
.B(n_290),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_272),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_342),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_299),
.A2(n_304),
.B1(n_308),
.B2(n_307),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_345),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_303),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_278),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_240),
.B1(n_266),
.B2(n_260),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_298),
.B(n_265),
.Y(n_349)
);

NAND2x1_ASAP7_75t_L g350 ( 
.A(n_289),
.B(n_228),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_307),
.A2(n_238),
.B1(n_253),
.B2(n_233),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_351),
.B(n_354),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_269),
.A2(n_247),
.B1(n_203),
.B2(n_261),
.Y(n_352)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_356),
.B(n_358),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_270),
.A2(n_207),
.B1(n_215),
.B2(n_252),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_359),
.Y(n_392)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_282),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_285),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_274),
.A2(n_254),
.B1(n_256),
.B2(n_289),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_305),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_375),
.C(n_383),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_350),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_369),
.B(n_328),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_341),
.A2(n_286),
.B1(n_295),
.B2(n_293),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_370),
.A2(n_373),
.B1(n_388),
.B2(n_390),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_347),
.A2(n_274),
.B1(n_317),
.B2(n_319),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_320),
.C(n_319),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_344),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_379),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_336),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_355),
.A2(n_274),
.B(n_320),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_382),
.A2(n_389),
.B(n_367),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_353),
.B(n_292),
.C(n_287),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_325),
.B(n_292),
.C(n_287),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_333),
.C(n_356),
.Y(n_414)
);

NOR3xp33_ASAP7_75t_SL g387 ( 
.A(n_348),
.B(n_302),
.C(n_283),
.Y(n_387)
);

AOI21xp33_ASAP7_75t_L g401 ( 
.A1(n_387),
.A2(n_340),
.B(n_334),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_324),
.A2(n_288),
.B1(n_317),
.B2(n_309),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_360),
.A2(n_313),
.B(n_315),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_327),
.A2(n_288),
.B1(n_309),
.B2(n_315),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_291),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_337),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_348),
.B(n_291),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_394),
.B(n_349),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_378),
.Y(n_395)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_395),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_375),
.Y(n_427)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_397),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_378),
.A2(n_362),
.B(n_382),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_405),
.Y(n_437)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_377),
.Y(n_399)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_399),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_412),
.C(n_416),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_401),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_364),
.Y(n_402)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_379),
.A2(n_323),
.B1(n_338),
.B2(n_359),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_404),
.A2(n_410),
.B1(n_423),
.B2(n_372),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_362),
.A2(n_331),
.B(n_330),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_406),
.B(n_409),
.Y(n_431)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_407),
.Y(n_447)
);

AOI21xp33_ASAP7_75t_L g408 ( 
.A1(n_376),
.A2(n_350),
.B(n_352),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_408),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_364),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_373),
.A2(n_351),
.B1(n_357),
.B2(n_321),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_371),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_390),
.B1(n_388),
.B2(n_381),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_349),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_403),
.C(n_420),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_361),
.B(n_332),
.Y(n_416)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_417),
.B(n_367),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_371),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_418),
.Y(n_436)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_374),
.Y(n_419)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_358),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_365),
.C(n_394),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_374),
.Y(n_421)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_385),
.Y(n_422)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_422),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_368),
.A2(n_346),
.B1(n_354),
.B2(n_342),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_429),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_386),
.Y(n_429)
);

AOI32xp33_ASAP7_75t_L g430 ( 
.A1(n_405),
.A2(n_365),
.A3(n_387),
.B1(n_366),
.B2(n_392),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_430),
.A2(n_413),
.B1(n_417),
.B2(n_410),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_411),
.A2(n_368),
.B1(n_370),
.B2(n_392),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_434),
.A2(n_413),
.B1(n_397),
.B2(n_393),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_449),
.C(n_395),
.Y(n_464)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_419),
.Y(n_441)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_441),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_442),
.A2(n_409),
.B1(n_398),
.B2(n_402),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_SL g444 ( 
.A(n_415),
.B(n_369),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_414),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_423),
.A2(n_384),
.B1(n_387),
.B2(n_391),
.Y(n_446)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_446),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_436),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_459),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_412),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_452),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_416),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_453),
.A2(n_460),
.B1(n_470),
.B2(n_439),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_399),
.Y(n_458)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_458),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_436),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_429),
.B(n_400),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_462),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_396),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_463),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_465),
.C(n_471),
.Y(n_478)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_469),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_407),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_428),
.A2(n_421),
.B1(n_422),
.B2(n_391),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_438),
.B(n_303),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_447),
.C(n_440),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_476),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_451),
.B(n_427),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_477),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_457),
.A2(n_428),
.B1(n_425),
.B2(n_445),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_461),
.B(n_437),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_432),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_481),
.C(n_464),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_432),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_466),
.B(n_394),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_488),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_466),
.B(n_425),
.Y(n_488)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_489),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_450),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_490),
.B(n_453),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_491),
.B(n_500),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_483),
.A2(n_456),
.B1(n_455),
.B2(n_468),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_496),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_485),
.A2(n_455),
.B(n_469),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_495),
.A2(n_501),
.B(n_503),
.Y(n_507)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_487),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_480),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_467),
.C(n_441),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_499),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_473),
.B(n_435),
.C(n_454),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_435),
.C(n_448),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_478),
.A2(n_384),
.B(n_380),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_479),
.A2(n_389),
.B(n_380),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_488),
.C(n_477),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_509),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_508),
.B(n_511),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_479),
.C(n_481),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_482),
.C(n_484),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_502),
.A2(n_385),
.B1(n_343),
.B2(n_345),
.Y(n_512)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_512),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_306),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_514),
.Y(n_522)
);

INVx11_ASAP7_75t_L g514 ( 
.A(n_495),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_494),
.B(n_296),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_515),
.A2(n_296),
.B1(n_313),
.B2(n_280),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_516),
.B(n_501),
.C(n_503),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_518),
.B(n_523),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_493),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_521),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_514),
.A2(n_492),
.B(n_504),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_509),
.B(n_493),
.C(n_318),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_525),
.B(n_507),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_525),
.Y(n_526)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_526),
.Y(n_533)
);

XOR2x2_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_507),
.Y(n_528)
);

AOI21xp33_ASAP7_75t_L g534 ( 
.A1(n_528),
.A2(n_527),
.B(n_530),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_522),
.Y(n_529)
);

O2A1O1Ixp33_ASAP7_75t_SL g536 ( 
.A1(n_529),
.A2(n_510),
.B(n_505),
.C(n_521),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_511),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_531),
.B(n_532),
.Y(n_535)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_534),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_536),
.A2(n_524),
.B(n_318),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_533),
.B(n_527),
.C(n_528),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_538),
.A2(n_539),
.B(n_535),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_537),
.C(n_280),
.Y(n_541)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_541),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_311),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_311),
.Y(n_544)
);


endmodule