module fake_jpeg_27221_n_97 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_97);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_97;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_26),
.Y(n_29)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_1),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_23),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_13),
.B1(n_19),
.B2(n_18),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_24),
.B2(n_27),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_18),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_37),
.B(n_39),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_17),
.B1(n_15),
.B2(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_27),
.C(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_22),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_53),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_26),
.B1(n_28),
.B2(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_54),
.B1(n_30),
.B2(n_22),
.Y(n_63)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_5),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_7),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_21),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_57),
.B1(n_59),
.B2(n_21),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_74),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_52),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_51),
.C(n_56),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_68),
.C(n_14),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_10),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_1),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_10),
.C(n_17),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_79),
.A2(n_72),
.B(n_63),
.C(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NOR2xp67_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_74),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_78),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_1),
.B(n_2),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_16),
.C(n_14),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_2),
.C(n_80),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_2),
.B(n_14),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_94),
.Y(n_97)
);


endmodule