module real_aes_14927_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_92;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
wire n_237;
wire n_91;
OAI221xp5_ASAP7_75t_L g528 ( .A1(n_0), .A2(n_529), .B1(n_534), .B2(n_545), .C(n_550), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_0), .A2(n_26), .B1(n_616), .B2(n_618), .Y(n_615) );
OA21x2_ASAP7_75t_L g108 ( .A1(n_1), .A2(n_39), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g238 ( .A(n_1), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_2), .A2(n_20), .B1(n_563), .B2(n_564), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_2), .A2(n_63), .B1(n_586), .B2(n_589), .Y(n_585) );
AND2x2_ASAP7_75t_L g163 ( .A(n_3), .B(n_155), .Y(n_163) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_4), .A2(n_74), .B1(n_83), .B2(n_187), .C(n_213), .Y(n_263) );
BUFx3_ASAP7_75t_L g495 ( .A(n_5), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_6), .B(n_140), .Y(n_159) );
INVx3_ASAP7_75t_L g492 ( .A(n_7), .Y(n_492) );
INVx2_ASAP7_75t_L g502 ( .A(n_8), .Y(n_502) );
INVx1_ASAP7_75t_L g606 ( .A(n_8), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_9), .B(n_113), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_10), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g88 ( .A(n_11), .Y(n_88) );
BUFx3_ASAP7_75t_L g115 ( .A(n_11), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_12), .B(n_125), .Y(n_170) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_13), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_14), .Y(n_224) );
BUFx10_ASAP7_75t_L g654 ( .A(n_15), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_16), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_17), .B(n_131), .Y(n_221) );
OAI21xp33_ASAP7_75t_L g332 ( .A1(n_17), .A2(n_51), .B(n_333), .Y(n_332) );
O2A1O1Ixp5_ASAP7_75t_L g264 ( .A1(n_18), .A2(n_157), .B(n_192), .C(n_265), .Y(n_264) );
OAI222xp33_ASAP7_75t_L g551 ( .A1(n_19), .A2(n_70), .B1(n_552), .B2(n_557), .C1(n_565), .C2(n_568), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_19), .Y(n_610) );
AOI221x1_ASAP7_75t_L g620 ( .A1(n_20), .A2(n_49), .B1(n_621), .B2(n_622), .C(n_624), .Y(n_620) );
AND2x2_ASAP7_75t_L g510 ( .A(n_21), .B(n_27), .Y(n_510) );
AND2x2_ASAP7_75t_L g517 ( .A(n_21), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g548 ( .A(n_21), .Y(n_548) );
INVx1_ASAP7_75t_L g93 ( .A(n_22), .Y(n_93) );
INVx2_ASAP7_75t_L g508 ( .A(n_23), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_24), .B(n_118), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_25), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g561 ( .A(n_26), .Y(n_561) );
INVx2_ASAP7_75t_L g518 ( .A(n_27), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_27), .B(n_548), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_28), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_29), .B(n_125), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_30), .A2(n_45), .B1(n_542), .B2(n_543), .Y(n_541) );
OAI211xp5_ASAP7_75t_L g575 ( .A1(n_30), .A2(n_576), .B(n_584), .C(n_614), .Y(n_575) );
AND2x4_ASAP7_75t_L g92 ( .A(n_31), .B(n_93), .Y(n_92) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_31), .Y(n_644) );
NAND2x1_ASAP7_75t_L g154 ( .A(n_32), .B(n_155), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_33), .Y(n_231) );
INVx1_ASAP7_75t_L g149 ( .A(n_34), .Y(n_149) );
INVx1_ASAP7_75t_L g500 ( .A(n_35), .Y(n_500) );
INVx1_ASAP7_75t_L g583 ( .A(n_35), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_36), .Y(n_249) );
AND2x2_ASAP7_75t_L g162 ( .A(n_37), .B(n_123), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_38), .B(n_117), .Y(n_206) );
INVx1_ASAP7_75t_L g239 ( .A(n_39), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_40), .B(n_140), .Y(n_258) );
INVx1_ASAP7_75t_L g109 ( .A(n_41), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_42), .B(n_123), .Y(n_169) );
OAI222xp33_ASAP7_75t_L g513 ( .A1(n_43), .A2(n_49), .B1(n_71), .B2(n_514), .C1(n_523), .C2(n_524), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_43), .A2(n_71), .B1(n_591), .B2(n_592), .C(n_596), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_44), .B(n_131), .Y(n_217) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_45), .A2(n_604), .B(n_607), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_46), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_47), .B(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_48), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g688 ( .A(n_48), .Y(n_688) );
AND2x2_ASAP7_75t_L g167 ( .A(n_50), .B(n_140), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_51), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_52), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_53), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_54), .B(n_117), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_55), .Y(n_266) );
NOR2xp67_ASAP7_75t_L g486 ( .A(n_56), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_57), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_58), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_59), .B(n_132), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_60), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g537 ( .A(n_61), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_61), .A2(n_70), .B1(n_629), .B2(n_631), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_62), .Y(n_233) );
INVx1_ASAP7_75t_L g560 ( .A(n_63), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_64), .B(n_186), .Y(n_214) );
INVx1_ASAP7_75t_L g671 ( .A(n_65), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_66), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_666) );
INVx2_ASAP7_75t_L g669 ( .A(n_66), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_67), .B(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_67), .Y(n_675) );
INVx1_ASAP7_75t_L g84 ( .A(n_68), .Y(n_84) );
BUFx3_ASAP7_75t_L g128 ( .A(n_68), .Y(n_128) );
INVx1_ASAP7_75t_L g158 ( .A(n_68), .Y(n_158) );
XNOR2xp5_ASAP7_75t_L g483 ( .A(n_69), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g507 ( .A(n_72), .Y(n_507) );
AND2x2_ASAP7_75t_L g527 ( .A(n_72), .B(n_508), .Y(n_527) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_72), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_73), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_73), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_75), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g494 ( .A(n_76), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_482), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_89), .Y(n_80) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_81), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_85), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_82), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_SL g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g234 ( .A(n_83), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_83), .A2(n_245), .B1(n_247), .B2(n_250), .Y(n_244) );
BUFx3_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g120 ( .A(n_84), .Y(n_120) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx2_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
INVx1_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
INVx2_ASAP7_75t_L g192 ( .A(n_87), .Y(n_192) );
INVx2_ASAP7_75t_L g230 ( .A(n_87), .Y(n_230) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx2_ASAP7_75t_L g188 ( .A(n_88), .Y(n_188) );
BUFx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
BUFx6f_ASAP7_75t_SL g129 ( .A(n_92), .Y(n_129) );
INVx3_ASAP7_75t_L g175 ( .A(n_92), .Y(n_175) );
INVx2_ASAP7_75t_L g216 ( .A(n_92), .Y(n_216) );
INVx1_ASAP7_75t_L g236 ( .A(n_92), .Y(n_236) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_93), .Y(n_642) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NOR2x1_ASAP7_75t_L g96 ( .A(n_97), .B(n_408), .Y(n_96) );
NAND4xp25_ASAP7_75t_L g97 ( .A(n_98), .B(n_316), .C(n_357), .D(n_390), .Y(n_97) );
NOR2xp33_ASAP7_75t_L g98 ( .A(n_99), .B(n_291), .Y(n_98) );
OAI222xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_198), .B1(n_259), .B2(n_274), .C1(n_279), .C2(n_286), .Y(n_99) );
NOR2xp67_ASAP7_75t_SL g100 ( .A(n_101), .B(n_176), .Y(n_100) );
AND2x2_ASAP7_75t_L g391 ( .A(n_101), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_134), .Y(n_101) );
AND2x2_ASAP7_75t_L g325 ( .A(n_102), .B(n_179), .Y(n_325) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_102), .Y(n_342) );
INVx1_ASAP7_75t_L g363 ( .A(n_102), .Y(n_363) );
INVx1_ASAP7_75t_L g412 ( .A(n_102), .Y(n_412) );
AND2x2_ASAP7_75t_L g452 ( .A(n_102), .B(n_383), .Y(n_452) );
INVx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g196 ( .A(n_103), .B(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g355 ( .A(n_103), .B(n_136), .Y(n_355) );
AND2x2_ASAP7_75t_L g426 ( .A(n_103), .B(n_278), .Y(n_426) );
BUFx3_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g313 ( .A(n_104), .Y(n_313) );
OAI21x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_110), .B(n_130), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g333 ( .A(n_107), .Y(n_333) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g133 ( .A(n_108), .Y(n_133) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_108), .Y(n_140) );
INVx1_ASAP7_75t_L g240 ( .A(n_109), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_121), .B(n_129), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_119), .Y(n_111) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g232 ( .A(n_114), .Y(n_232) );
INVx1_ASAP7_75t_L g246 ( .A(n_114), .Y(n_246) );
INVx2_ASAP7_75t_L g254 ( .A(n_114), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_114), .B(n_266), .Y(n_265) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g118 ( .A(n_115), .Y(n_118) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_115), .Y(n_126) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
INVx1_ASAP7_75t_L g184 ( .A(n_118), .Y(n_184) );
INVx2_ASAP7_75t_L g226 ( .A(n_118), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_119), .A2(n_183), .B(n_185), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_119), .A2(n_211), .B(n_214), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_119), .A2(n_252), .B(n_255), .Y(n_251) );
BUFx10_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_124), .B(n_127), .Y(n_121) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx3_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
INVx3_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g144 ( .A(n_128), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_128), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g228 ( .A(n_128), .Y(n_228) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_129), .A2(n_142), .B(n_151), .Y(n_141) );
INVx1_ASAP7_75t_L g194 ( .A(n_129), .Y(n_194) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_132), .B(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g324 ( .A(n_134), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g343 ( .A(n_134), .B(n_312), .Y(n_343) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g416 ( .A(n_135), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_160), .Y(n_135) );
INVx2_ASAP7_75t_L g197 ( .A(n_136), .Y(n_197) );
AND2x4_ASAP7_75t_SL g290 ( .A(n_136), .B(n_195), .Y(n_290) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_136), .Y(n_301) );
INVx1_ASAP7_75t_L g315 ( .A(n_136), .Y(n_315) );
INVxp67_ASAP7_75t_L g384 ( .A(n_136), .Y(n_384) );
INVx1_ASAP7_75t_L g401 ( .A(n_136), .Y(n_401) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_141), .B(n_159), .Y(n_137) );
INVx1_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVxp33_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_140), .Y(n_203) );
INVx1_ASAP7_75t_L g270 ( .A(n_140), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B(n_147), .Y(n_142) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
AOI21x1_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_154), .B(n_156), .Y(n_151) );
INVx1_ASAP7_75t_L g208 ( .A(n_153), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_156), .A2(n_190), .B(n_191), .Y(n_189) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g209 ( .A(n_157), .Y(n_209) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g165 ( .A(n_158), .Y(n_165) );
INVx2_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
INVx1_ASAP7_75t_L g278 ( .A(n_160), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_160), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g370 ( .A(n_160), .B(n_277), .Y(n_370) );
OR2x2_ASAP7_75t_L g405 ( .A(n_160), .B(n_179), .Y(n_405) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_166), .B(n_172), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_164), .Y(n_161) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g171 ( .A(n_165), .Y(n_171) );
NOR2xp67_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
AOI21xp33_ASAP7_75t_L g172 ( .A1(n_167), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_171), .Y(n_168) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR3xp33_ASAP7_75t_L g262 ( .A(n_175), .B(n_263), .C(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_196), .Y(n_177) );
AND2x2_ASAP7_75t_L g352 ( .A(n_178), .B(n_353), .Y(n_352) );
BUFx3_ASAP7_75t_L g373 ( .A(n_178), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_178), .B(n_363), .Y(n_454) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_195), .Y(n_178) );
INVx3_ASAP7_75t_L g277 ( .A(n_179), .Y(n_277) );
INVx1_ASAP7_75t_L g288 ( .A(n_179), .Y(n_288) );
AND2x2_ASAP7_75t_L g383 ( .A(n_179), .B(n_384), .Y(n_383) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_179), .Y(n_389) );
INVx1_ASAP7_75t_L g450 ( .A(n_179), .Y(n_450) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_189), .B(n_193), .Y(n_181) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g213 ( .A(n_188), .Y(n_213) );
BUFx2_ASAP7_75t_L g341 ( .A(n_195), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_196), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g435 ( .A(n_196), .Y(n_435) );
AND2x2_ASAP7_75t_L g480 ( .A(n_196), .B(n_450), .Y(n_480) );
AND2x2_ASAP7_75t_L g423 ( .A(n_197), .B(n_313), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_199), .B(n_218), .Y(n_198) );
INVx2_ASAP7_75t_L g294 ( .A(n_199), .Y(n_294) );
AND2x2_ASAP7_75t_L g356 ( .A(n_199), .B(n_304), .Y(n_356) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g339 ( .A(n_200), .B(n_285), .Y(n_339) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g345 ( .A(n_201), .B(n_261), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .B(n_217), .Y(n_201) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_202), .A2(n_243), .B(n_258), .Y(n_242) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_202), .A2(n_243), .B(n_258), .Y(n_283) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_202), .A2(n_204), .B(n_217), .Y(n_308) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OAI21x1_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_210), .B(n_215), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_209), .Y(n_205) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_SL g257 ( .A(n_216), .Y(n_257) );
AND2x2_ASAP7_75t_L g402 ( .A(n_218), .B(n_345), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_218), .B(n_294), .Y(n_413) );
AND2x2_ASAP7_75t_L g418 ( .A(n_218), .B(n_312), .Y(n_418) );
AND2x2_ASAP7_75t_L g432 ( .A(n_218), .B(n_339), .Y(n_432) );
AND2x2_ASAP7_75t_L g462 ( .A(n_218), .B(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_241), .Y(n_218) );
INVx1_ASAP7_75t_L g446 ( .A(n_219), .Y(n_446) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g273 ( .A(n_220), .Y(n_273) );
INVx2_ASAP7_75t_L g296 ( .A(n_220), .Y(n_296) );
AND2x2_ASAP7_75t_L g304 ( .A(n_220), .B(n_242), .Y(n_304) );
AND2x2_ASAP7_75t_L g444 ( .A(n_220), .B(n_282), .Y(n_444) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_222), .B(n_332), .C(n_334), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .C(n_235), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_227), .C(n_228), .Y(n_223) );
INVx2_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
OAI221xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B1(n_232), .B2(n_233), .C(n_234), .Y(n_229) );
INVx2_ASAP7_75t_L g256 ( .A(n_230), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g336 ( .A(n_237), .Y(n_336) );
AOI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_240), .Y(n_237) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_238), .A2(n_239), .B(n_240), .Y(n_267) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x4_ASAP7_75t_L g295 ( .A(n_242), .B(n_296), .Y(n_295) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_251), .B(n_257), .Y(n_243) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_248), .A2(n_646), .B1(n_665), .B2(n_678), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_248), .A2(n_665), .B1(n_680), .B2(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_271), .Y(n_259) );
AND2x2_ASAP7_75t_L g297 ( .A(n_260), .B(n_281), .Y(n_297) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g285 ( .A(n_261), .Y(n_285) );
AND2x2_ASAP7_75t_L g306 ( .A(n_261), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g420 ( .A(n_261), .Y(n_420) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_267), .B(n_268), .Y(n_261) );
NAND2xp33_ASAP7_75t_L g334 ( .A(n_262), .B(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_R g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_272), .Y(n_359) );
AND2x2_ASAP7_75t_L g433 ( .A(n_272), .B(n_306), .Y(n_433) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g284 ( .A(n_273), .B(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g298 ( .A(n_275), .B(n_299), .Y(n_298) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_284), .Y(n_279) );
AND2x2_ASAP7_75t_L g305 ( .A(n_280), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g338 ( .A(n_281), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g441 ( .A(n_281), .Y(n_441) );
BUFx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx3_ASAP7_75t_L g322 ( .A(n_283), .Y(n_322) );
AND2x4_ASAP7_75t_L g463 ( .A(n_285), .B(n_379), .Y(n_463) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g392 ( .A(n_287), .Y(n_392) );
AOI32xp33_ASAP7_75t_L g417 ( .A1(n_287), .A2(n_418), .A3(n_419), .B1(n_421), .B2(n_422), .Y(n_417) );
AND2x4_ASAP7_75t_L g459 ( .A(n_287), .B(n_416), .Y(n_459) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g400 ( .A(n_288), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g366 ( .A(n_289), .Y(n_366) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g319 ( .A(n_290), .B(n_312), .Y(n_319) );
AND2x2_ASAP7_75t_L g350 ( .A(n_290), .B(n_311), .Y(n_350) );
AND2x2_ASAP7_75t_L g388 ( .A(n_290), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_302), .Y(n_291) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_297), .B(n_298), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g303 ( .A(n_294), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g475 ( .A(n_294), .B(n_407), .Y(n_475) );
AND2x2_ASAP7_75t_L g348 ( .A(n_295), .B(n_345), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_295), .A2(n_325), .B1(n_352), .B2(n_356), .Y(n_351) );
AND2x2_ASAP7_75t_L g421 ( .A(n_295), .B(n_306), .Y(n_421) );
AND2x2_ASAP7_75t_L g429 ( .A(n_295), .B(n_339), .Y(n_429) );
AND2x4_ASAP7_75t_SL g481 ( .A(n_295), .B(n_463), .Y(n_481) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVxp67_ASAP7_75t_L g369 ( .A(n_301), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B(n_309), .Y(n_302) );
AND2x2_ASAP7_75t_L g375 ( .A(n_304), .B(n_345), .Y(n_375) );
INVx1_ASAP7_75t_L g393 ( .A(n_304), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_306), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g379 ( .A(n_307), .Y(n_379) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_L g329 ( .A(n_308), .Y(n_329) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g477 ( .A(n_312), .B(n_370), .Y(n_477) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g411 ( .A(n_314), .B(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_346), .Y(n_316) );
OAI221xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .B1(n_323), .B2(n_326), .C(n_337), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g344 ( .A(n_321), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g381 ( .A(n_322), .Y(n_381) );
OR2x2_ASAP7_75t_L g407 ( .A(n_322), .B(n_331), .Y(n_407) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g394 ( .A(n_328), .Y(n_394) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g386 ( .A(n_329), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g380 ( .A(n_331), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g387 ( .A(n_331), .Y(n_387) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B1(n_343), .B2(n_344), .Y(n_337) );
AND2x2_ASAP7_75t_L g358 ( .A(n_338), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g397 ( .A(n_341), .Y(n_397) );
AND2x2_ASAP7_75t_L g422 ( .A(n_341), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g398 ( .A(n_342), .Y(n_398) );
AND2x2_ASAP7_75t_L g445 ( .A(n_345), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_345), .B(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g472 ( .A(n_345), .B(n_444), .Y(n_472) );
OAI21xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_349), .B(n_351), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_350), .B(n_392), .Y(n_439) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g449 ( .A(n_355), .B(n_450), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B(n_371), .Y(n_357) );
NAND3xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_364), .C(n_367), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g403 ( .A(n_362), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B1(n_376), .B2(n_382), .C(n_385), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_377), .B(n_415), .Y(n_414) );
NOR2x1p5_ASAP7_75t_SL g377 ( .A(n_378), .B(n_380), .Y(n_377) );
AND2x2_ASAP7_75t_L g443 ( .A(n_378), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_378), .B(n_418), .Y(n_457) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_386), .A2(n_465), .B(n_468), .Y(n_464) );
AOI322xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .A3(n_394), .B1(n_395), .B2(n_402), .C1(n_403), .C2(n_406), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_399), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g427 ( .A(n_399), .Y(n_427) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_405), .Y(n_436) );
INVx2_ASAP7_75t_L g469 ( .A(n_405), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_405), .B(n_423), .Y(n_474) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_407), .B(n_454), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_437), .C(n_455), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_424), .Y(n_409) );
OAI211xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B(n_414), .C(n_417), .Y(n_410) );
INVx2_ASAP7_75t_L g479 ( .A(n_411), .Y(n_479) );
BUFx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI221x1_ASAP7_75t_L g442 ( .A1(n_422), .A2(n_443), .B1(n_445), .B2(n_447), .C(n_453), .Y(n_442) );
AND2x2_ASAP7_75t_L g468 ( .A(n_423), .B(n_469), .Y(n_468) );
OAI21xp33_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_428), .B(n_430), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_433), .B2(n_434), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_433), .B(n_441), .Y(n_440) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B(n_442), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI21xp33_ASAP7_75t_SL g456 ( .A1(n_440), .A2(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g467 ( .A(n_446), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_449), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NOR3xp33_ASAP7_75t_SL g455 ( .A(n_456), .B(n_460), .C(n_470), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_461), .B(n_464), .Y(n_460) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .B1(n_475), .B2(n_476), .C(n_478), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B(n_481), .Y(n_478) );
OAI221xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_636), .B2(n_645), .C(n_684), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_484), .A2(n_685), .B1(n_687), .B2(n_689), .Y(n_684) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_486), .B(n_511), .Y(n_485) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_503), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_496), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g509 ( .A(n_492), .B(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g516 ( .A(n_492), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g549 ( .A(n_492), .Y(n_549) );
AND2x4_ASAP7_75t_SL g556 ( .A(n_492), .B(n_510), .Y(n_556) );
INVx2_ASAP7_75t_L g635 ( .A(n_492), .Y(n_635) );
INVx2_ASAP7_75t_L g578 ( .A(n_493), .Y(n_578) );
OR2x2_ASAP7_75t_L g629 ( .A(n_493), .B(n_630), .Y(n_629) );
OR2x6_ASAP7_75t_SL g631 ( .A(n_493), .B(n_632), .Y(n_631) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g598 ( .A(n_494), .Y(n_598) );
BUFx2_ASAP7_75t_L g627 ( .A(n_494), .Y(n_627) );
OR2x2_ASAP7_75t_L g597 ( .A(n_495), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g602 ( .A(n_495), .B(n_598), .Y(n_602) );
AND2x4_ASAP7_75t_L g626 ( .A(n_495), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g619 ( .A(n_498), .Y(n_619) );
BUFx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx12f_ASAP7_75t_L g591 ( .A(n_499), .Y(n_591) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
AND2x4_ASAP7_75t_L g605 ( .A(n_500), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g613 ( .A(n_500), .Y(n_613) );
AND2x4_ASAP7_75t_L g595 ( .A(n_501), .B(n_582), .Y(n_595) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g581 ( .A(n_502), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g588 ( .A(n_502), .B(n_583), .Y(n_588) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_509), .Y(n_504) );
OR2x6_ASAP7_75t_L g523 ( .A(n_505), .B(n_515), .Y(n_523) );
INVx3_ASAP7_75t_L g536 ( .A(n_505), .Y(n_536) );
INVx2_ASAP7_75t_SL g559 ( .A(n_505), .Y(n_559) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
INVx2_ASAP7_75t_L g521 ( .A(n_507), .Y(n_521) );
AND2x4_ASAP7_75t_L g532 ( .A(n_507), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g522 ( .A(n_508), .Y(n_522) );
INVx2_ASAP7_75t_L g533 ( .A(n_508), .Y(n_533) );
OR2x6_ASAP7_75t_L g550 ( .A(n_509), .B(n_519), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_574), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_528), .C(n_551), .Y(n_512) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
OR2x2_ASAP7_75t_L g524 ( .A(n_515), .B(n_525), .Y(n_524) );
OR2x6_ASAP7_75t_L g529 ( .A(n_515), .B(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g567 ( .A(n_518), .B(n_548), .Y(n_567) );
INVx3_ASAP7_75t_L g539 ( .A(n_519), .Y(n_539) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2x1p5_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
BUFx3_ASAP7_75t_L g555 ( .A(n_522), .Y(n_555) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx12f_ASAP7_75t_SL g542 ( .A(n_526), .Y(n_542) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g563 ( .A(n_527), .Y(n_563) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx5_ASAP7_75t_L g544 ( .A(n_532), .Y(n_544) );
OAI221xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_537), .B1(n_538), .B2(n_540), .C(n_541), .Y(n_534) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_538), .A2(n_558), .B1(n_560), .B2(n_561), .C(n_562), .Y(n_557) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_540), .A2(n_594), .B1(n_608), .B2(n_610), .C(n_611), .Y(n_607) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g564 ( .A(n_544), .Y(n_564) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x6_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
OR2x2_ASAP7_75t_L g565 ( .A(n_549), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x4_ASAP7_75t_L g569 ( .A(n_556), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI21xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_628), .B(n_633), .Y(n_574) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx5_ASAP7_75t_L g589 ( .A(n_580), .Y(n_589) );
BUFx3_ASAP7_75t_L g617 ( .A(n_580), .Y(n_617) );
INVx3_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_590), .B1(n_599), .B2(n_603), .Y(n_584) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx5_ASAP7_75t_L g621 ( .A(n_587), .Y(n_621) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx5_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g632 ( .A(n_595), .Y(n_632) );
BUFx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_597), .Y(n_656) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g664 ( .A(n_602), .Y(n_664) );
CKINVDCx8_ASAP7_75t_R g604 ( .A(n_605), .Y(n_604) );
INVx8_ASAP7_75t_L g630 ( .A(n_605), .Y(n_630) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_606), .Y(n_609) );
INVx1_ASAP7_75t_L g655 ( .A(n_606), .Y(n_655) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_620), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx4_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
BUFx6f_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_638), .Y(n_637) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_643), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AO21x2_ASAP7_75t_L g691 ( .A1(n_641), .A2(n_692), .B(n_693), .Y(n_691) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g650 ( .A(n_642), .Y(n_650) );
AND2x2_ASAP7_75t_L g693 ( .A(n_643), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_644), .B(n_650), .Y(n_649) );
BUFx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx5_ASAP7_75t_L g686 ( .A(n_647), .Y(n_686) );
AND2x6_ASAP7_75t_L g647 ( .A(n_648), .B(n_657), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVxp67_ASAP7_75t_L g682 ( .A(n_649), .Y(n_682) );
INVx1_ASAP7_75t_L g694 ( .A(n_650), .Y(n_694) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_652), .B(n_661), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .C(n_656), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
CKINVDCx11_ASAP7_75t_R g659 ( .A(n_654), .Y(n_659) );
AND2x4_ASAP7_75t_L g662 ( .A(n_655), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
XOR2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_670), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B1(n_673), .B2(n_677), .Y(n_670) );
INVx2_ASAP7_75t_L g677 ( .A(n_671), .Y(n_677) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx4f_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx4_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_691), .Y(n_690) );
endmodule