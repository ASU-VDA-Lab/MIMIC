module fake_jpeg_27803_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_53),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_31),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_34),
.B(n_21),
.C(n_30),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_31),
.B1(n_16),
.B2(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_57),
.B1(n_45),
.B2(n_21),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_31),
.B1(n_18),
.B2(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_23),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_67),
.B(n_72),
.Y(n_126)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_23),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_73),
.A2(n_89),
.B(n_93),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_35),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_101),
.B(n_35),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_81),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_79),
.A2(n_98),
.B1(n_100),
.B2(n_28),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_24),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_82),
.B(n_84),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_37),
.B1(n_41),
.B2(n_43),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_37),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_85),
.Y(n_138)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_61),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_93),
.Y(n_132)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_38),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_97),
.Y(n_133)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_26),
.B1(n_20),
.B2(n_41),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_26),
.B1(n_20),
.B2(n_41),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_30),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_102),
.B(n_104),
.CI(n_107),
.CON(n_127),
.SN(n_127)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_46),
.B(n_15),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_47),
.B(n_11),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_53),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_109),
.B1(n_43),
.B2(n_44),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_61),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_17),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_116),
.C(n_117),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_113),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_0),
.B(n_1),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_0),
.B(n_1),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_43),
.B1(n_38),
.B2(n_40),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_88),
.B1(n_87),
.B2(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_35),
.C(n_40),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_40),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_121),
.B(n_39),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_39),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_102),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_67),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_71),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_142),
.B(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_144),
.B(n_147),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_164),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_94),
.B1(n_97),
.B2(n_75),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_154),
.B1(n_160),
.B2(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_152),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_166),
.B1(n_129),
.B2(n_111),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_167),
.B(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_106),
.B1(n_92),
.B2(n_95),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_74),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_118),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_161),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_101),
.B1(n_69),
.B2(n_85),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_66),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_87),
.B1(n_109),
.B2(n_68),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_163),
.A2(n_111),
.B1(n_138),
.B2(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_96),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_130),
.B(n_120),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_103),
.B(n_2),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_86),
.B1(n_105),
.B2(n_35),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_32),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_186),
.B1(n_152),
.B2(n_149),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_127),
.B(n_132),
.C(n_114),
.D(n_113),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_174),
.B(n_185),
.CI(n_27),
.CON(n_219),
.SN(n_219)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_169),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_175),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_178),
.B(n_180),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_116),
.Y(n_178)
);

OA21x2_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_127),
.B(n_131),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_181),
.B(n_10),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_146),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_184),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_127),
.B(n_115),
.C(n_30),
.D(n_139),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_203),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_134),
.C(n_119),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_32),
.C(n_28),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_138),
.B1(n_135),
.B2(n_77),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_192),
.B1(n_197),
.B2(n_22),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_167),
.A2(n_19),
.B(n_25),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_193),
.B(n_196),
.Y(n_205)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_163),
.B1(n_150),
.B2(n_154),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_25),
.B(n_19),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_142),
.B(n_19),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_156),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_118),
.B(n_25),
.C(n_22),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_32),
.B1(n_28),
.B2(n_27),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_0),
.B(n_2),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_145),
.B(n_32),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_4),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_12),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_144),
.B1(n_147),
.B2(n_161),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_204),
.A2(n_208),
.B1(n_209),
.B2(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_212),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_194),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_158),
.B1(n_157),
.B2(n_159),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_211),
.C(n_222),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_44),
.C(n_22),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_28),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_44),
.Y(n_218)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_230),
.Y(n_236)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_224),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_27),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_199),
.C(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_225),
.A2(n_201),
.B1(n_196),
.B2(n_178),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_3),
.Y(n_227)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_27),
.C(n_5),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_231),
.C(n_177),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_229),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_10),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_210),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_8),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_196),
.B1(n_219),
.B2(n_227),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_250),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_245),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_200),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_178),
.B1(n_203),
.B2(n_185),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_253),
.B1(n_205),
.B2(n_193),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_214),
.B1(n_218),
.B2(n_204),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_248),
.B(n_219),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_198),
.Y(n_249)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_208),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_180),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_246),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_183),
.B1(n_174),
.B2(n_196),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_211),
.C(n_215),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_266),
.C(n_275),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_261),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_218),
.B(n_191),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_264),
.A2(n_270),
.B(n_237),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_268),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_227),
.C(n_228),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_230),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_272),
.Y(n_277)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_262),
.B1(n_264),
.B2(n_263),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_11),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_236),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_244),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_8),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_286),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_249),
.B(n_255),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_290),
.B1(n_266),
.B2(n_258),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_252),
.B(n_240),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_288),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_236),
.B1(n_248),
.B2(n_245),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_238),
.B(n_5),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_257),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_258),
.C(n_256),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_298),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_295),
.B(n_303),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_300),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_6),
.C(n_7),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_7),
.Y(n_300)
);

A2O1A1Ixp33_ASAP7_75t_SL g301 ( 
.A1(n_279),
.A2(n_283),
.B(n_281),
.C(n_276),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_278),
.B(n_286),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_7),
.C(n_8),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_276),
.B1(n_289),
.B2(n_282),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_307),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_291),
.B(n_284),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_296),
.B(n_301),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_311),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_285),
.B1(n_12),
.B2(n_13),
.Y(n_311)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_310),
.Y(n_315)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_300),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_318),
.A2(n_319),
.B(n_306),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_297),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_322),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_325),
.C(n_316),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_321),
.A2(n_316),
.B(n_314),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_323),
.C(n_301),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_307),
.C(n_12),
.Y(n_328)
);

AOI221xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_4),
.B1(n_13),
.B2(n_14),
.C(n_108),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_14),
.Y(n_330)
);


endmodule