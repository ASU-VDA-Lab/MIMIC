module real_jpeg_2545_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_0),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_0),
.A2(n_35),
.B1(n_37),
.B2(n_141),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_0),
.A2(n_69),
.B1(n_71),
.B2(n_141),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_0),
.A2(n_58),
.B1(n_64),
.B2(n_141),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_2),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_2),
.A2(n_35),
.B1(n_37),
.B2(n_175),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_2),
.A2(n_69),
.B1(n_71),
.B2(n_175),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_2),
.A2(n_58),
.B1(n_64),
.B2(n_175),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_6),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_85),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_6),
.A2(n_69),
.B1(n_71),
.B2(n_85),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g211 ( 
.A1(n_6),
.A2(n_58),
.B1(n_64),
.B2(n_85),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_7),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_7),
.A2(n_35),
.B1(n_37),
.B2(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_68),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_7),
.A2(n_58),
.B1(n_64),
.B2(n_68),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_8),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_35),
.B1(n_37),
.B2(n_83),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_8),
.A2(n_69),
.B1(n_71),
.B2(n_83),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_8),
.A2(n_58),
.B1(n_64),
.B2(n_83),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_9),
.A2(n_40),
.B1(n_58),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_9),
.A2(n_40),
.B1(n_69),
.B2(n_71),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_9),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_10),
.A2(n_43),
.B1(n_69),
.B2(n_71),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_10),
.A2(n_35),
.B1(n_37),
.B2(n_43),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_10),
.A2(n_43),
.B1(n_58),
.B2(n_64),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_11),
.A2(n_35),
.B1(n_37),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_91),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_11),
.A2(n_69),
.B1(n_71),
.B2(n_91),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_11),
.A2(n_58),
.B1(n_64),
.B2(n_91),
.Y(n_187)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_16),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_16),
.A2(n_35),
.B1(n_37),
.B2(n_194),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_16),
.A2(n_69),
.B1(n_71),
.B2(n_194),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_16),
.A2(n_58),
.B1(n_64),
.B2(n_194),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_18),
.B(n_29),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_18),
.B(n_38),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_18),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_18),
.A2(n_29),
.B(n_184),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_18),
.B(n_94),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g252 ( 
.A1(n_18),
.A2(n_37),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_18),
.B(n_58),
.C(n_74),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_18),
.A2(n_69),
.B1(n_71),
.B2(n_220),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_18),
.B(n_61),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_18),
.B(n_78),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_46),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_41),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_38),
.B(n_39),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_27),
.A2(n_38),
.B1(n_140),
.B2(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_27),
.A2(n_38),
.B1(n_42),
.B2(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_34),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g183 ( 
.A1(n_30),
.A2(n_33),
.A3(n_37),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_32),
.B(n_35),
.Y(n_185)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_34),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_34),
.A2(n_81),
.B1(n_84),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_34),
.A2(n_81),
.B1(n_82),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_34),
.A2(n_81),
.B1(n_104),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_34),
.A2(n_81),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_34),
.A2(n_81),
.B1(n_193),
.B2(n_231),
.Y(n_230)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_35),
.A2(n_37),
.B1(n_95),
.B2(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_35),
.B(n_220),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_37),
.A2(n_69),
.A3(n_95),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_41),
.B(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_45),
.B(n_329),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_325),
.B(n_327),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_313),
.B(n_324),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_155),
.B(n_310),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_142),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_115),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_51),
.B(n_115),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_86),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_52),
.B(n_101),
.C(n_113),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_79),
.B(n_80),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_53),
.A2(n_54),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.Y(n_54)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_55),
.A2(n_79),
.B1(n_80),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_55),
.A2(n_65),
.B1(n_66),
.B2(n_79),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_62),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_56),
.A2(n_60),
.B1(n_129),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_56),
.A2(n_60),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_56),
.A2(n_60),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_57),
.A2(n_61),
.B1(n_63),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_57),
.A2(n_61),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_57),
.A2(n_61),
.B1(n_187),
.B2(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_57),
.A2(n_61),
.B1(n_224),
.B2(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_57),
.A2(n_61),
.B1(n_220),
.B2(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_57),
.A2(n_61),
.B1(n_273),
.B2(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_58),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_64),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_58),
.B(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_72),
.B1(n_78),
.B2(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_69),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AO22x2_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_71),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_69),
.B(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_71),
.B(n_96),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_77),
.B1(n_78),
.B2(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_78),
.B(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_72),
.A2(n_78),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_72),
.A2(n_78),
.B1(n_216),
.B2(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_72),
.A2(n_78),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_72),
.A2(n_78),
.B1(n_243),
.B2(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_76),
.A2(n_133),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_76),
.A2(n_168),
.B1(n_215),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_101),
.B1(n_113),
.B2(n_114),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_88),
.B(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_99),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B1(n_94),
.B2(n_98),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_93),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_94),
.B1(n_98),
.B2(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_92),
.A2(n_94),
.B1(n_136),
.B2(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_92),
.A2(n_94),
.B(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_93),
.A2(n_111),
.B1(n_137),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_93),
.A2(n_137),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_93),
.A2(n_137),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_93),
.A2(n_137),
.B1(n_190),
.B2(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_93),
.A2(n_137),
.B1(n_205),
.B2(n_252),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_103),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_107),
.C(n_109),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_103),
.B(n_146),
.C(n_153),
.Y(n_314)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_112),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_107),
.B(n_149),
.C(n_151),
.Y(n_323)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_123),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_134),
.C(n_138),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_125),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_126),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_196)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_138),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_142),
.A2(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_154),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_143),
.B(n_154),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_153),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_150),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_152),
.Y(n_320)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_176),
.B(n_309),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_157),
.B(n_159),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_164),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.C(n_173),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_166),
.B(n_169),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_173),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_199),
.B(n_308),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_197),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_178),
.B(n_197),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_196),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_179),
.B(n_196),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_181),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.C(n_192),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_182),
.B(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_186),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_189),
.B(n_192),
.Y(n_299)
);

AOI31xp33_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_293),
.A3(n_302),
.B(n_305),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_238),
.B(n_292),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_226),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_202),
.B(n_226),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_213),
.C(n_217),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_203),
.B(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_208),
.C(n_212),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_213),
.B(n_217),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_226),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_226),
.B(n_303),
.Y(n_306)
);

FAx1_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.CI(n_229),
.CON(n_226),
.SN(n_226)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_230),
.B(n_233),
.C(n_237),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_287),
.B(n_291),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_256),
.B(n_286),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_245),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_251),
.C(n_254),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_267),
.B(n_285),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_265),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_279),
.B(n_284),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_274),
.B(n_278),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_297),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_315),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_323),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_319),
.B1(n_321),
.B2(n_322),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_321),
.C(n_323),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_326),
.Y(n_329)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule