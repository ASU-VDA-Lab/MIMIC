module real_jpeg_24705_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_1),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_1),
.A2(n_60),
.B(n_65),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_1),
.B(n_90),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_1),
.A2(n_110),
.B1(n_201),
.B2(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_1),
.A2(n_26),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_1),
.B(n_50),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_69),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_2),
.A2(n_34),
.B1(n_69),
.B2(n_128),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_5),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_174),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_174),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_5),
.A2(n_33),
.B1(n_38),
.B2(n_174),
.Y(n_282)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_32),
.B1(n_39),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_52),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_7),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_7),
.A2(n_52),
.B1(n_64),
.B2(n_65),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_8),
.A2(n_31),
.B1(n_38),
.B2(n_41),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_41),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_8),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_41),
.B1(n_64),
.B2(n_65),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_9),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_9),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_9),
.A2(n_35),
.B1(n_64),
.B2(n_65),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_33),
.B1(n_38),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_11),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_154),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_154),
.Y(n_278)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_13),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_183),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_183),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_13),
.A2(n_38),
.B1(n_45),
.B2(n_183),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_15),
.Y(n_116)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_15),
.Y(n_149)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_15),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_91),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_19),
.B(n_91),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_85),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_47),
.B1(n_83),
.B2(n_84),
.Y(n_20)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_54),
.C(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_21),
.A2(n_83),
.B1(n_93),
.B2(n_95),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_30),
.B(n_36),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_22),
.B(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_22),
.A2(n_43),
.B1(n_153),
.B2(n_294),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_23),
.A2(n_24),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g263 ( 
.A1(n_23),
.A2(n_27),
.A3(n_39),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_24),
.B(n_26),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_26),
.A2(n_27),
.B1(n_75),
.B2(n_76),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_26),
.A2(n_58),
.A3(n_75),
.B1(n_217),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_27),
.B(n_171),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_34),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_34),
.B(n_171),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_37),
.B(n_50),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_38),
.A2(n_171),
.B(n_264),
.Y(n_281)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_42),
.A2(n_50),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_42),
.A2(n_50),
.B1(n_282),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_43),
.A2(n_126),
.B(n_129),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_43),
.A2(n_153),
.B(n_155),
.Y(n_152)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_50),
.B(n_127),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_70),
.B1(n_71),
.B2(n_82),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_82),
.B1(n_86),
.B2(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_67),
.B(n_68),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_55),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_55),
.A2(n_67),
.B1(n_173),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_55),
.A2(n_67),
.B1(n_182),
.B2(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_55),
.A2(n_68),
.B(n_123),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_58),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_57),
.B(n_76),
.Y(n_226)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_58),
.A2(n_62),
.B(n_171),
.C(n_176),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_63),
.B(n_102),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_63),
.A2(n_120),
.B1(n_121),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_63),
.A2(n_120),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_63),
.B(n_171),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_63),
.A2(n_100),
.B(n_151),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_64),
.B(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_73),
.A2(n_79),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_74),
.A2(n_78),
.B(n_105),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_74),
.A2(n_215),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_77),
.A2(n_89),
.B(n_218),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_87),
.B1(n_90),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_79),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_79),
.A2(n_90),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_79),
.A2(n_90),
.B1(n_241),
.B2(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_106),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_92),
.A2(n_96),
.B1(n_97),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_98),
.B(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_99),
.A2(n_120),
.B(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_124),
.B(n_125),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_108),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_124),
.B1(n_125),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_109),
.A2(n_119),
.B1(n_124),
.B2(n_327),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_114),
.B(n_117),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_110),
.A2(n_147),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_110),
.A2(n_114),
.B1(n_191),
.B2(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_110),
.A2(n_117),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_110),
.A2(n_228),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_111),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_111),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_266)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_114),
.Y(n_268)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_116),
.Y(n_248)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_118),
.B(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_119),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_122),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_160),
.B(n_342),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_157),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_134),
.B(n_157),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.C(n_141),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_135),
.A2(n_139),
.B1(n_140),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_135),
.Y(n_331)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_141),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_152),
.C(n_156),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_142),
.A2(n_143),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_144),
.B(n_150),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_145),
.A2(n_247),
.B(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_146),
.B(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_171),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_152),
.B(n_156),
.Y(n_324)
);

AOI311xp33_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_320),
.A3(n_332),
.B(n_336),
.C(n_337),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_284),
.C(n_315),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_258),
.B(n_283),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_234),
.B(n_257),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_210),
.B(n_233),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_187),
.B(n_209),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_177),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_167),
.B(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_175),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_169),
.B1(n_175),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_185),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_184),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_184),
.C(n_185),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_197),
.B(n_208),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_195),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_202),
.B(n_207),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_224),
.B1(n_231),
.B2(n_232),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_213)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_223),
.C(n_231),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_227),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_236),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_250),
.B2(n_251),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_253),
.C(n_255),
.Y(n_259)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_244),
.C(n_245),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_252),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_253),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_259),
.B(n_260),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_275),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_261)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_274),
.C(n_275),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_266),
.B1(n_270),
.B2(n_271),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_270),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_266),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_280),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_279),
.C(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI21xp33_ASAP7_75t_L g338 ( 
.A1(n_285),
.A2(n_339),
.B(n_340),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_300),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_286),
.B(n_300),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_295),
.C(n_296),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_287),
.A2(n_288),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_291),
.C(n_292),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_295),
.B(n_296),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_299),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_300)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_310),
.B2(n_311),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_311),
.C(n_314),
.Y(n_334)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_309),
.Y(n_303)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_308),
.C(n_309),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_310),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_317),
.Y(n_339)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_321),
.A2(n_333),
.B(n_338),
.C(n_341),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_329),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_329),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.C(n_328),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_323),
.B(n_326),
.CI(n_328),
.CON(n_335),
.SN(n_335)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_334),
.B(n_335),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_335),
.Y(n_344)
);


endmodule