module fake_jpeg_22765_n_75 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_38;
wire n_74;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_69;
wire n_40;
wire n_71;
wire n_35;
wire n_48;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_32;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_0),
.Y(n_52)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_40),
.B1(n_41),
.B2(n_37),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_51),
.C(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_2),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_49),
.B1(n_48),
.B2(n_46),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_61),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_54),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_59),
.B(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_36),
.B1(n_5),
.B2(n_6),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_34),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_3),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_64),
.C(n_9),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_4),
.C(n_8),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_62),
.B1(n_67),
.B2(n_13),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_11),
.C(n_12),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_14),
.B(n_15),
.Y(n_71)
);

AOI322xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_21),
.C1(n_22),
.C2(n_24),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_31),
.Y(n_74)
);

FAx1_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_25),
.CI(n_26),
.CON(n_75),
.SN(n_75)
);


endmodule