module fake_netlist_1_6945_n_28 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_28);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx3_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_2), .Y(n_11) );
INVx2_ASAP7_75t_SL g12 ( .A(n_6), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_4), .B(n_1), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_7), .B(n_4), .Y(n_15) );
AOI21x1_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_8), .B(n_9), .Y(n_16) );
NAND3xp33_ASAP7_75t_SL g17 ( .A(n_11), .B(n_1), .C(n_2), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_14), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
OAI22xp5_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_13), .B1(n_12), .B2(n_10), .Y(n_20) );
INVx5_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_17), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
AOI221x1_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_20), .B1(n_10), .B2(n_22), .C(n_15), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
BUFx12f_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OAI22xp5_ASAP7_75t_SL g27 ( .A1(n_26), .A2(n_3), .B1(n_5), .B2(n_21), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_26), .B1(n_25), .B2(n_21), .Y(n_28) );
endmodule