module real_jpeg_21591_n_16 (n_338, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_338;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_0),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_0),
.A2(n_24),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_0),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_0),
.A2(n_9),
.B1(n_24),
.B2(n_44),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_22),
.B1(n_25),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_1),
.A2(n_41),
.B1(n_48),
.B2(n_53),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_1),
.A2(n_9),
.B1(n_44),
.B2(n_53),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_53),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_26),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_2),
.A2(n_9),
.B(n_14),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_2),
.A2(n_41),
.B1(n_48),
.B2(n_119),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_2),
.A2(n_93),
.B1(n_98),
.B2(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_2),
.B(n_73),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_2),
.B(n_29),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_2),
.A2(n_29),
.B(n_206),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_3),
.A2(n_22),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_9),
.B1(n_44),
.B2(n_55),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_3),
.A2(n_41),
.B1(n_48),
.B2(n_55),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_55),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_4),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_4),
.A2(n_22),
.B1(n_25),
.B2(n_114),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_4),
.A2(n_9),
.B1(n_44),
.B2(n_114),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_4),
.A2(n_41),
.B1(n_48),
.B2(n_114),
.Y(n_194)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_6),
.A2(n_22),
.B1(n_25),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_6),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_121),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_6),
.A2(n_41),
.B1(n_48),
.B2(n_121),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_6),
.A2(n_9),
.B1(n_44),
.B2(n_121),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_7),
.B(n_44),
.Y(n_94)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_8),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_9),
.B1(n_44),
.B2(n_116),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_8),
.A2(n_41),
.B1(n_48),
.B2(n_116),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_8),
.A2(n_22),
.B1(n_25),
.B2(n_116),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_9),
.A2(n_14),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_9),
.A2(n_11),
.B1(n_32),
.B2(n_44),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_11),
.A2(n_22),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_11),
.A2(n_32),
.B1(n_41),
.B2(n_48),
.Y(n_103)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_41),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_15),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_81),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_79),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_35),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_20),
.A2(n_51),
.B(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_21),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_26),
.B(n_28),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_28),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g118 ( 
.A(n_22),
.B(n_119),
.CON(n_118),
.SN(n_118)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_26),
.B(n_31),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_26),
.A2(n_33),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_27),
.A2(n_34),
.B1(n_118),
.B2(n_125),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_27),
.A2(n_41),
.A3(n_63),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_28),
.B(n_29),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_29),
.A2(n_61),
.B(n_62),
.C(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_29),
.B(n_62),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_30),
.A2(n_52),
.B(n_56),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_33),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_71),
.C(n_75),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_37),
.A2(n_38),
.B1(n_332),
.B2(n_334),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_49),
.C(n_57),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_39),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_39),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_39),
.A2(n_57),
.B1(n_58),
.B2(n_312),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_43),
.B(n_46),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_40),
.A2(n_46),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_40),
.A2(n_43),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_40),
.A2(n_43),
.B1(n_174),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_40),
.A2(n_43),
.B1(n_194),
.B2(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_40),
.A2(n_213),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_40),
.A2(n_43),
.B1(n_101),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_40),
.A2(n_109),
.B(n_246),
.Y(n_280)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_43),
.B(n_119),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_44),
.B(n_183),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_45),
.A2(n_48),
.B(n_119),
.C(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_47),
.B(n_110),
.Y(n_228)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_48),
.B(n_62),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_49),
.A2(n_50),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_51),
.A2(n_56),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_51),
.A2(n_56),
.B1(n_132),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_51),
.A2(n_78),
.B(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_60),
.A2(n_66),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_61),
.A2(n_67),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_61),
.A2(n_67),
.B1(n_152),
.B2(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_61),
.B(n_70),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_61),
.A2(n_65),
.B(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_61),
.A2(n_67),
.B1(n_271),
.B2(n_292),
.Y(n_291)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_66),
.A2(n_73),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_66),
.A2(n_74),
.B(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_66),
.A2(n_257),
.B(n_315),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_71),
.A2(n_72),
.B1(n_75),
.B2(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_75),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_329),
.B(n_335),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_305),
.A3(n_324),
.B1(n_327),
.B2(n_328),
.C(n_338),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_284),
.B(n_304),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_262),
.B(n_283),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_154),
.B(n_237),
.C(n_261),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_137),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_87),
.B(n_137),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_122),
.B2(n_136),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_106),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_90),
.B(n_106),
.C(n_136),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_100),
.B2(n_105),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_91),
.B(n_105),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_93),
.A2(n_146),
.B1(n_163),
.B2(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_93),
.A2(n_166),
.B(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_93),
.A2(n_146),
.B(n_279),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_94),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_94),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_94),
.A2(n_97),
.B(n_198),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_98),
.B(n_119),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_99),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_102),
.B(n_228),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_117),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_115),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_123),
.B(n_129),
.C(n_134),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_126),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_138),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.C(n_150),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_144),
.A2(n_145),
.B1(n_149),
.B2(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_147),
.B(n_196),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_150),
.B(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_236),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_231),
.B(n_235),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_218),
.B(n_230),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_200),
.B(n_217),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_186),
.B(n_199),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_175),
.B(n_185),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_171),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_180),
.B(n_184),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_178),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_187),
.B(n_188),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_201)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_198),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_202),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_208),
.B1(n_215),
.B2(n_216),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_211),
.B1(n_212),
.B2(n_214),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_209),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_220),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_227),
.C(n_229),
.Y(n_232)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2x2_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_232),
.B(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_239),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_259),
.B2(n_260),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_248),
.C(n_260),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_258),
.Y(n_248)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_256),
.C(n_258),
.Y(n_282)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_264),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_282),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_275),
.B2(n_276),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_276),
.C(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_272),
.C(n_274),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_270),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_278),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_277),
.A2(n_295),
.B(n_299),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_280),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_280),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_285),
.B(n_286),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_302),
.B2(n_303),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_294),
.C(n_303),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B(n_293),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_292),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_307),
.C(n_316),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g326 ( 
.A(n_293),
.B(n_307),
.CI(n_316),
.CON(n_326),
.SN(n_326)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_299),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_302),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_317),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_317),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_309),
.B1(n_319),
.B2(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_312),
.C(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_322),
.C(n_323),
.Y(n_330)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_326),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_332),
.Y(n_334)
);


endmodule