module fake_jpeg_22715_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_17),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_44),
.B(n_45),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_22),
.B1(n_16),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_20),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_22),
.B1(n_16),
.B2(n_21),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_28),
.B1(n_29),
.B2(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_20),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_28),
.B1(n_32),
.B2(n_24),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_62),
.Y(n_109)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_61),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_63),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_37),
.B1(n_18),
.B2(n_29),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_70),
.B1(n_75),
.B2(n_82),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_28),
.B1(n_24),
.B2(n_32),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_32),
.B1(n_24),
.B2(n_15),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_71),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_37),
.B1(n_41),
.B2(n_34),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_15),
.B1(n_21),
.B2(n_18),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_73),
.B(n_51),
.C(n_23),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_39),
.A3(n_36),
.B1(n_29),
.B2(n_15),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_79),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_41),
.B1(n_34),
.B2(n_25),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_35),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_39),
.B1(n_20),
.B2(n_36),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_83),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_39),
.B(n_55),
.C(n_35),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_96),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_39),
.B1(n_51),
.B2(n_55),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_110),
.B1(n_61),
.B2(n_86),
.Y(n_128)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_111),
.Y(n_142)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_66),
.C(n_67),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_39),
.C(n_17),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_55),
.B1(n_39),
.B2(n_26),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_26),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_40),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_59),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_118),
.B(n_119),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_72),
.B1(n_70),
.B2(n_75),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_134),
.B1(n_105),
.B2(n_99),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_123),
.A2(n_91),
.B(n_103),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_132),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_95),
.B1(n_102),
.B2(n_104),
.Y(n_151)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_135),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_131),
.C(n_136),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_40),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_40),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_113),
.A2(n_74),
.B1(n_76),
.B2(n_69),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_137),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_61),
.B1(n_27),
.B2(n_30),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_140),
.B1(n_145),
.B2(n_100),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_141),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_27),
.B1(n_30),
.B2(n_58),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_112),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_93),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_100),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_144),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_89),
.A2(n_60),
.B1(n_31),
.B2(n_23),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_146),
.A2(n_151),
.B1(n_154),
.B2(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_148),
.B(n_150),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_149),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_114),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_152),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_95),
.B1(n_116),
.B2(n_107),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_166),
.C(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_156),
.B(n_158),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_0),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_157),
.A2(n_170),
.B(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_160),
.Y(n_188)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_19),
.B1(n_23),
.B2(n_104),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_163),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_97),
.B1(n_104),
.B2(n_98),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_164),
.A2(n_133),
.B1(n_92),
.B2(n_23),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_165),
.B(n_167),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_97),
.C(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_169),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_103),
.B(n_91),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_9),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_122),
.A2(n_93),
.B1(n_90),
.B2(n_96),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_120),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_143),
.B(n_118),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_190),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_185),
.C(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_130),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_121),
.C(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

AO22x1_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_128),
.B1(n_138),
.B2(n_135),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_93),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_195),
.C(n_177),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_92),
.C(n_31),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_153),
.B(n_163),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_19),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_146),
.A2(n_164),
.B1(n_154),
.B2(n_168),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_9),
.C(n_14),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_151),
.A2(n_19),
.B1(n_13),
.B2(n_12),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_1),
.B(n_2),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_13),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_216),
.C(n_224),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_158),
.C(n_156),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_204),
.A2(n_151),
.B1(n_175),
.B2(n_173),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_218),
.A2(n_189),
.B1(n_181),
.B2(n_195),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_150),
.B1(n_151),
.B2(n_148),
.Y(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_157),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_149),
.C(n_160),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_161),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_152),
.C(n_161),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_198),
.C(n_191),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_188),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_206),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_209),
.Y(n_236)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_179),
.B1(n_200),
.B2(n_196),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_238),
.B1(n_252),
.B2(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_208),
.B(n_197),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_196),
.B1(n_192),
.B2(n_203),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_202),
.B1(n_192),
.B2(n_183),
.Y(n_241)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_208),
.C(n_184),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_250),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_216),
.C(n_224),
.Y(n_255)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_247),
.A2(n_249),
.B1(n_210),
.B2(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_190),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_211),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_194),
.B1(n_186),
.B2(n_205),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_12),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_13),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_258),
.B1(n_267),
.B2(n_249),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_3),
.C(n_4),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_256),
.B(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_243),
.B(n_215),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_242),
.A2(n_213),
.B1(n_225),
.B2(n_214),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_4),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_213),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_266),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_222),
.C(n_214),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_264),
.C(n_10),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_223),
.C(n_221),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_269),
.A2(n_252),
.B1(n_239),
.B2(n_240),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_SL g271 ( 
.A1(n_259),
.A2(n_237),
.B(n_238),
.C(n_234),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_272),
.B(n_282),
.Y(n_288)
);

XNOR2x1_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_245),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_263),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_261),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_247),
.B1(n_240),
.B2(n_248),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_244),
.B1(n_253),
.B2(n_5),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_262),
.B1(n_270),
.B2(n_269),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_10),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_10),
.C(n_11),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_4),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_286),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_291),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_272),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_266),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_11),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_292),
.B(n_4),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_293),
.B(n_6),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_295),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_300),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_281),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_276),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_271),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_301),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_310),
.Y(n_313)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_271),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_271),
.B(n_294),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_307),
.B(n_308),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_309),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_313),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_306),
.B(n_305),
.C(n_295),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_315),
.B(n_296),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_6),
.B(n_7),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_7),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_7),
.B(n_305),
.Y(n_320)
);


endmodule