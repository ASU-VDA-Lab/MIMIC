module fake_jpeg_2630_n_66 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_66);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_66;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_19),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_20),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_28),
.B1(n_26),
.B2(n_24),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_24),
.B(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_39),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_37),
.B1(n_25),
.B2(n_33),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_21),
.Y(n_46)
);

NOR4xp25_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_24),
.C(n_21),
.D(n_35),
.Y(n_48)
);

OAI322xp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_51),
.A3(n_0),
.B1(n_1),
.B2(n_3),
.C1(n_4),
.C2(n_6),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_52),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_25),
.C(n_20),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_46),
.B1(n_33),
.B2(n_2),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_56),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_51),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_12),
.C(n_3),
.Y(n_60)
);

OAI211xp5_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_15),
.B(n_14),
.C(n_13),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_57),
.B(n_53),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_58),
.C(n_4),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_62),
.B(n_1),
.C(n_6),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_63),
.A2(n_7),
.B(n_8),
.Y(n_64)
);

AOI222xp33_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_53),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_11),
.Y(n_66)
);


endmodule