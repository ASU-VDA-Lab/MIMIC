module fake_jpeg_31356_n_441 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_441);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_45),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_47),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_19),
.B(n_8),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_41),
.Y(n_111)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_63),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_72),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_76),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_78),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_21),
.B(n_18),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_34),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_85),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_56),
.B(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_92),
.B(n_108),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_39),
.B1(n_37),
.B2(n_43),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_95),
.A2(n_42),
.B1(n_57),
.B2(n_22),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_49),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_117),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_45),
.A2(n_29),
.B1(n_40),
.B2(n_28),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_42),
.B1(n_27),
.B2(n_28),
.Y(n_170)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_48),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_54),
.B(n_33),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_26),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_49),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_123),
.B(n_128),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_48),
.B(n_29),
.Y(n_128)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_74),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_143),
.Y(n_195)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_89),
.B(n_69),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_74),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_23),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_148),
.Y(n_186)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_23),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_100),
.A2(n_88),
.B1(n_80),
.B2(n_75),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_152),
.B1(n_133),
.B2(n_95),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_162),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_62),
.B1(n_66),
.B2(n_83),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_170),
.B1(n_171),
.B2(n_93),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_112),
.B1(n_98),
.B2(n_104),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_153),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_71),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_164),
.B(n_126),
.Y(n_196)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_93),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_118),
.Y(n_169)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_176),
.B(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_107),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_194),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_153),
.A2(n_132),
.B1(n_129),
.B2(n_40),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_152),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_129),
.B1(n_28),
.B2(n_27),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_143),
.B1(n_145),
.B2(n_153),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_138),
.B(n_103),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_198),
.Y(n_225)
);

NOR2x1p5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_164),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_201),
.A2(n_205),
.B(n_130),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_209),
.B1(n_215),
.B2(n_226),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_212),
.Y(n_229)
);

HAxp5_ASAP7_75t_SL g205 ( 
.A(n_194),
.B(n_138),
.CON(n_205),
.SN(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_140),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_210),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_211),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_161),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_214),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_183),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_143),
.B1(n_171),
.B2(n_135),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_139),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_199),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_164),
.B(n_116),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_145),
.B(n_164),
.Y(n_240)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_166),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_178),
.B1(n_197),
.B2(n_116),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_169),
.B1(n_144),
.B2(n_167),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_213),
.Y(n_227)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_195),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_248),
.C(n_222),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_195),
.B1(n_196),
.B2(n_182),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_234),
.A2(n_249),
.B1(n_96),
.B2(n_177),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_214),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_237),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_211),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_217),
.A2(n_182),
.B1(n_181),
.B2(n_199),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_226),
.B1(n_202),
.B2(n_201),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_246),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_240),
.A2(n_177),
.B(n_193),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_215),
.B(n_217),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_218),
.B(n_212),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_247),
.A2(n_240),
.B(n_238),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_174),
.C(n_187),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_187),
.B1(n_174),
.B2(n_200),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_208),
.B1(n_219),
.B2(n_225),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_232),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_252),
.B(n_269),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_254),
.A2(n_250),
.B1(n_158),
.B2(n_141),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_275),
.Y(n_286)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_201),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_274),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_257),
.A2(n_261),
.B(n_271),
.Y(n_307)
);

AND2x6_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_201),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_258),
.B(n_280),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_40),
.Y(n_310)
);

NOR4xp25_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_218),
.C(n_210),
.D(n_216),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_244),
.Y(n_288)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_206),
.Y(n_267)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_241),
.A2(n_223),
.B(n_203),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_172),
.Y(n_270)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_200),
.C(n_172),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_147),
.C(n_114),
.Y(n_299)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_230),
.A2(n_219),
.B1(n_208),
.B2(n_224),
.Y(n_274)
);

OA22x2_ASAP7_75t_L g275 ( 
.A1(n_230),
.A2(n_224),
.B1(n_159),
.B2(n_160),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_242),
.B1(n_235),
.B2(n_227),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_231),
.B(n_193),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_281),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_229),
.B(n_26),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_278),
.B(n_279),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_229),
.B(n_33),
.Y(n_279)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_115),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_285),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_284),
.A2(n_297),
.B1(n_273),
.B2(n_266),
.Y(n_326)
);

NOR4xp25_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_242),
.C(n_248),
.D(n_237),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_233),
.B1(n_243),
.B2(n_239),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_287),
.A2(n_290),
.B1(n_297),
.B2(n_291),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_299),
.C(n_300),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_233),
.B1(n_243),
.B2(n_250),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_253),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_305),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_264),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_303),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_121),
.C(n_165),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_270),
.B(n_27),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_264),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_268),
.B(n_60),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_306),
.B(n_269),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_313),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_272),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_286),
.A2(n_263),
.B1(n_260),
.B2(n_276),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_290),
.Y(n_337)
);

OAI22x1_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_261),
.B1(n_275),
.B2(n_280),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_286),
.A2(n_275),
.B1(n_255),
.B2(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_319),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_267),
.C(n_277),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_309),
.C(n_292),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_258),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_315),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_283),
.A2(n_259),
.B(n_271),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_323),
.B(n_325),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_259),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_330),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_283),
.A2(n_275),
.B(n_281),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_326),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_265),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_302),
.Y(n_343)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_295),
.Y(n_328)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_328),
.Y(n_345)
);

A2O1A1Ixp33_ASAP7_75t_SL g329 ( 
.A1(n_307),
.A2(n_178),
.B(n_133),
.C(n_90),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_329),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_154),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_284),
.A2(n_168),
.B1(n_155),
.B2(n_22),
.Y(n_331)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_334),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_291),
.A2(n_163),
.B(n_142),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_335),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_337),
.A2(n_317),
.B1(n_334),
.B2(n_329),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_320),
.A2(n_298),
.B1(n_286),
.B2(n_308),
.Y(n_338)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_350),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_332),
.A2(n_298),
.B1(n_304),
.B2(n_287),
.Y(n_344)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_304),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_354),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_314),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_335),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_349),
.B(n_346),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_301),
.C(n_293),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_329),
.C(n_90),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_301),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_318),
.A2(n_86),
.B1(n_126),
.B2(n_122),
.Y(n_355)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_154),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_358),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_321),
.B(n_122),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_312),
.Y(n_360)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_339),
.B(n_323),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_364),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_316),
.Y(n_365)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_325),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_366),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_311),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_368),
.B(n_370),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_329),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_374),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_16),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_373),
.A2(n_375),
.B(n_376),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_354),
.C(n_350),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_352),
.A2(n_15),
.B(n_18),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_352),
.A2(n_133),
.B1(n_101),
.B2(n_51),
.Y(n_377)
);

INVx11_ASAP7_75t_L g387 ( 
.A(n_377),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_71),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_341),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_359),
.A2(n_342),
.B1(n_340),
.B2(n_348),
.Y(n_379)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_379),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_101),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_385),
.B(n_369),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_392),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_358),
.C(n_343),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_32),
.C(n_101),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_371),
.A2(n_356),
.B(n_14),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_391),
.A2(n_14),
.B(n_17),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_369),
.B(n_12),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_363),
.C(n_367),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_394),
.B(n_395),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_365),
.C(n_372),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_396),
.B(n_401),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_383),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_399),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_382),
.A2(n_360),
.B(n_361),
.Y(n_398)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_398),
.A2(n_379),
.B(n_387),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_362),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_376),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_404),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_388),
.A2(n_378),
.B(n_60),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_405),
.B(n_392),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_385),
.C(n_386),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_410),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_398),
.A2(n_388),
.B(n_401),
.Y(n_412)
);

AOI322xp5_ASAP7_75t_L g419 ( 
.A1(n_412),
.A2(n_413),
.A3(n_403),
.B1(n_32),
.B2(n_6),
.C1(n_15),
.C2(n_16),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_400),
.A2(n_390),
.B1(n_387),
.B2(n_389),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_416),
.Y(n_423)
);

AOI21xp33_ASAP7_75t_L g415 ( 
.A1(n_405),
.A2(n_8),
.B(n_11),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g418 ( 
.A(n_415),
.Y(n_418)
);

NOR3xp33_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_22),
.C(n_8),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_419),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_5),
.Y(n_420)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_420),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_411),
.A2(n_87),
.B1(n_6),
.B2(n_12),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_2),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_16),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_424),
.B(n_425),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_12),
.Y(n_425)
);

AOI322xp5_ASAP7_75t_L g426 ( 
.A1(n_410),
.A2(n_416),
.A3(n_32),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_1),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_426),
.A2(n_0),
.B(n_2),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_423),
.A2(n_32),
.B(n_1),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_428),
.B(n_431),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_432),
.B(n_418),
.Y(n_435)
);

AOI322xp5_ASAP7_75t_L g433 ( 
.A1(n_427),
.A2(n_3),
.A3(n_4),
.B1(n_418),
.B2(n_422),
.C1(n_429),
.C2(n_430),
.Y(n_433)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_433),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_435),
.B(n_434),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_437),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_438),
.B(n_436),
.C(n_3),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_439),
.A2(n_3),
.B(n_4),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_4),
.Y(n_441)
);


endmodule