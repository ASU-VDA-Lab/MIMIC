module fake_jpeg_30950_n_498 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_498);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_498;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_54),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_61),
.Y(n_108)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_67),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_13),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_0),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_13),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_68),
.B(n_70),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_31),
.B(n_11),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_72),
.B(n_82),
.Y(n_139)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_40),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_34),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_83),
.B(n_90),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_33),
.B(n_10),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_43),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_50),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_103),
.B(n_109),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_65),
.B(n_50),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_46),
.B(n_45),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_114),
.B(n_132),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_126),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_55),
.Y(n_126)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_33),
.Y(n_132)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_66),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_52),
.Y(n_162)
);

INVx6_ASAP7_75t_SL g144 ( 
.A(n_52),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_144),
.Y(n_196)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_53),
.Y(n_149)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_57),
.Y(n_153)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_58),
.Y(n_154)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_60),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_159),
.B(n_177),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_160),
.B(n_171),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_162),
.B(n_167),
.Y(n_225)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_166),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_37),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_37),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_168),
.B(n_173),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_123),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_170),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_108),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_174),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_45),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_83),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_102),
.A2(n_19),
.B1(n_78),
.B2(n_79),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_188),
.B1(n_91),
.B2(n_154),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_105),
.A2(n_80),
.B1(n_81),
.B2(n_99),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_176),
.A2(n_142),
.B1(n_127),
.B2(n_106),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_76),
.C(n_69),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_111),
.B(n_46),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_195),
.Y(n_236)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_118),
.A2(n_62),
.B1(n_56),
.B2(n_94),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_197),
.B1(n_148),
.B2(n_138),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_112),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_198),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_124),
.A2(n_19),
.B1(n_32),
.B2(n_42),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_123),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_49),
.C(n_30),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_17),
.C(n_86),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_140),
.B(n_32),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_156),
.A2(n_30),
.B1(n_29),
.B2(n_16),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_112),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_118),
.B(n_42),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_44),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_152),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_200),
.B(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_152),
.B(n_25),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_100),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_136),
.B(n_86),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_203),
.Y(n_239)
);

BUFx2_ASAP7_75t_R g204 ( 
.A(n_115),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_204),
.A2(n_153),
.B1(n_125),
.B2(n_17),
.Y(n_220)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_104),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_209),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_29),
.B(n_16),
.C(n_17),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_211),
.B(n_238),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_215),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_137),
.B1(n_133),
.B2(n_151),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_137),
.B1(n_133),
.B2(n_147),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_208),
.A2(n_177),
.B1(n_199),
.B2(n_194),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_176),
.A2(n_155),
.B1(n_148),
.B2(n_147),
.Y(n_216)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_221),
.Y(n_273)
);

AO21x2_ASAP7_75t_SL g281 ( 
.A1(n_223),
.A2(n_182),
.B(n_158),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_159),
.A2(n_44),
.B1(n_25),
.B2(n_24),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_241),
.B(n_244),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_74),
.B(n_106),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_159),
.A2(n_1),
.B(n_4),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_129),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_247),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_186),
.A2(n_141),
.B1(n_138),
.B2(n_129),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_157),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_251),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_207),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_253),
.B(n_261),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_204),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_268),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_256),
.Y(n_323)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_258),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_196),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_189),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_262),
.B(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_263),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_170),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_230),
.B(n_197),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_276),
.Y(n_297)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_164),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_161),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_269),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_235),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_270),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_242),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_272),
.Y(n_295)
);

NOR3xp33_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_206),
.C(n_161),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_274),
.Y(n_298)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_232),
.A2(n_47),
.B(n_190),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_278),
.A2(n_226),
.B(n_219),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_163),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_280),
.A2(n_285),
.B(n_238),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g313 ( 
.A1(n_281),
.A2(n_287),
.B(n_237),
.C(n_192),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_178),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_282),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_185),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_288),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_250),
.Y(n_284)
);

INVx8_ASAP7_75t_L g317 ( 
.A(n_284),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g285 ( 
.A(n_241),
.B(n_169),
.Y(n_285)
);

INVx3_ASAP7_75t_SL g286 ( 
.A(n_246),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_286),
.Y(n_304)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_236),
.B(n_169),
.Y(n_288)
);

XOR2x1_ASAP7_75t_SL g289 ( 
.A(n_271),
.B(n_211),
.Y(n_289)
);

XNOR2x1_ASAP7_75t_SL g326 ( 
.A(n_289),
.B(n_255),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_260),
.A2(n_244),
.B(n_240),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_291),
.A2(n_318),
.B(n_324),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_221),
.B1(n_245),
.B2(n_247),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_292),
.A2(n_303),
.B1(n_316),
.B2(n_265),
.Y(n_338)
);

AND2x2_ASAP7_75t_SL g299 ( 
.A(n_260),
.B(n_212),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_299),
.Y(n_352)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_302),
.A2(n_310),
.B(n_313),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_273),
.A2(n_223),
.B1(n_220),
.B2(n_122),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_259),
.B(n_223),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_308),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_259),
.B(n_223),
.Y(n_308)
);

AO22x1_ASAP7_75t_SL g309 ( 
.A1(n_281),
.A2(n_248),
.B1(n_218),
.B2(n_227),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_277),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_285),
.A2(n_233),
.B(n_205),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_266),
.A2(n_122),
.B1(n_128),
.B2(n_141),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_312),
.A2(n_315),
.B1(n_286),
.B2(n_272),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_281),
.A2(n_128),
.B1(n_181),
.B2(n_183),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_279),
.A2(n_277),
.B1(n_271),
.B2(n_288),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_278),
.A2(n_233),
.B(n_237),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_283),
.B(n_227),
.C(n_226),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_257),
.C(n_258),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_256),
.Y(n_325)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_328),
.Y(n_361)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_329),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_290),
.B(n_270),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_330),
.B(n_336),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_341),
.C(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_332),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_333),
.A2(n_338),
.B1(n_353),
.B2(n_312),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_335),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_315),
.A2(n_280),
.B1(n_281),
.B2(n_268),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_319),
.B(n_252),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_306),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_356),
.Y(n_372)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_299),
.B(n_263),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_276),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_323),
.Y(n_343)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_291),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_267),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_346),
.Y(n_384)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_349),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_297),
.A2(n_265),
.B1(n_254),
.B2(n_252),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_351),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_254),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_303),
.A2(n_286),
.B1(n_179),
.B2(n_181),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_289),
.A2(n_287),
.B(n_231),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_354),
.A2(n_318),
.B(n_324),
.Y(n_380)
);

INVx3_ASAP7_75t_SL g355 ( 
.A(n_317),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_293),
.Y(n_356)
);

AND2x6_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_320),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_360),
.A2(n_380),
.B(n_370),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_351),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_369),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_368),
.A2(n_334),
.B1(n_337),
.B2(n_309),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_340),
.B(n_314),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_302),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_348),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_322),
.Y(n_375)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_375),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_294),
.Y(n_376)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_321),
.Y(n_377)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_338),
.A2(n_298),
.B1(n_295),
.B2(n_292),
.Y(n_378)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_349),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_381),
.B(n_385),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_353),
.A2(n_295),
.B1(n_310),
.B2(n_308),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_373),
.A2(n_352),
.B1(n_343),
.B2(n_365),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_387),
.A2(n_399),
.B1(n_406),
.B2(n_383),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_357),
.A2(n_347),
.B1(n_354),
.B2(n_344),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_388),
.A2(n_392),
.B1(n_382),
.B2(n_374),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_393),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_371),
.B(n_348),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_391),
.B(n_396),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_357),
.A2(n_347),
.B1(n_344),
.B2(n_335),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_372),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_350),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_400),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_398),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_367),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_366),
.B(n_342),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_361),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_341),
.C(n_307),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_382),
.C(n_358),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_309),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_410),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_379),
.Y(n_404)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_404),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_363),
.B(n_304),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_405),
.B(n_363),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_368),
.A2(n_313),
.B1(n_304),
.B2(n_311),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_380),
.A2(n_313),
.B(n_329),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_408),
.A2(n_313),
.B(n_383),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_359),
.B(n_300),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_359),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_412),
.B(n_415),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_375),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_418),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_360),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_420),
.A2(n_399),
.B1(n_358),
.B2(n_362),
.Y(n_444)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_404),
.Y(n_421)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_421),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_426),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_429),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_374),
.C(n_365),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_428),
.C(n_410),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_361),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_409),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_431),
.B(n_439),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_413),
.Y(n_432)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_432),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_392),
.C(n_407),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_433),
.B(n_436),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_206),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_388),
.C(n_403),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_389),
.C(n_398),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_437),
.B(n_182),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_430),
.A2(n_425),
.B(n_424),
.Y(n_439)
);

BUFx12_ASAP7_75t_L g440 ( 
.A(n_411),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_242),
.Y(n_455)
);

OAI21xp33_ASAP7_75t_L g442 ( 
.A1(n_411),
.A2(n_386),
.B(n_406),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_444),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_412),
.C(n_426),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_450),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_441),
.B(n_415),
.C(n_427),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_446),
.A2(n_362),
.B1(n_427),
.B2(n_158),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_455),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_275),
.C(n_231),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_456),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_438),
.Y(n_454)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_454),
.Y(n_466)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_219),
.C(n_179),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_460),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_47),
.C(n_183),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_10),
.C(n_11),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_462),
.B(n_432),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_453),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_463),
.B(n_455),
.Y(n_478)
);

XNOR2x1_ASAP7_75t_SL g464 ( 
.A(n_448),
.B(n_440),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_464),
.A2(n_4),
.B(n_6),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_470),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_459),
.B(n_434),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_454),
.A2(n_443),
.B1(n_446),
.B2(n_442),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_7),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_461),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_474),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_461),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_476),
.B(n_477),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_473),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_478),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_469),
.A2(n_440),
.B(n_5),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_480),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_467),
.C(n_471),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_483),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_466),
.C(n_471),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_486),
.A2(n_478),
.B(n_475),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_490),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_485),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_487),
.B(n_7),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_484),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_492),
.B(n_484),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_494),
.A2(n_493),
.B(n_488),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_495),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_496),
.B(n_7),
.Y(n_497)
);

XOR2x2_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_7),
.Y(n_498)
);


endmodule