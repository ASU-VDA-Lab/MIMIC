module fake_jpeg_4974_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_SL g11 ( 
.A(n_0),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_21),
.B(n_28),
.C(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_21),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_53),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_32),
.B(n_26),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_54),
.B(n_24),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_12),
.B1(n_14),
.B2(n_22),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_49),
.B1(n_4),
.B2(n_6),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_12),
.B1(n_14),
.B2(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_32),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_55),
.B(n_51),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_60),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_54),
.C(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_79),
.B(n_81),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_69),
.C(n_70),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_60),
.B1(n_48),
.B2(n_44),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_65),
.B1(n_71),
.B2(n_69),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_57),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_80),
.B1(n_63),
.B2(n_53),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_85),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_74),
.C(n_84),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_91),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_80),
.B1(n_76),
.B2(n_81),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_90),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_63),
.B1(n_68),
.B2(n_75),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

XOR2x2_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_86),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_4),
.B(n_6),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_90),
.A3(n_93),
.B1(n_85),
.B2(n_87),
.C1(n_47),
.C2(n_9),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_99),
.B(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_96),
.Y(n_101)
);

AOI21x1_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_97),
.B(n_7),
.Y(n_103)
);

OAI321xp33_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_102),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C(n_2),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);


endmodule