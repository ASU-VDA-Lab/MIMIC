module fake_jpeg_5870_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_8),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_51),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_35),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_17),
.B(n_26),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_57),
.B1(n_30),
.B2(n_29),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_58),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_18),
.B1(n_21),
.B2(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_18),
.B1(n_21),
.B2(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_37),
.B1(n_29),
.B2(n_25),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_34),
.A2(n_21),
.B1(n_26),
.B2(n_31),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_42),
.B1(n_34),
.B2(n_41),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_39),
.B1(n_42),
.B2(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_40),
.Y(n_94)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_67),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_36),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_34),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_75),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_78),
.B1(n_82),
.B2(n_84),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_76),
.B1(n_85),
.B2(n_62),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_74),
.Y(n_116)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_34),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_42),
.B1(n_39),
.B2(n_31),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_91),
.B1(n_22),
.B2(n_9),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_39),
.B1(n_41),
.B2(n_35),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_86),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_33),
.B1(n_26),
.B2(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_40),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_41),
.B1(n_37),
.B2(n_36),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_30),
.B1(n_16),
.B2(n_19),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_45),
.B(n_36),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_25),
.B1(n_19),
.B2(n_16),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_53),
.B1(n_47),
.B2(n_48),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_98),
.B1(n_74),
.B2(n_68),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_47),
.B1(n_48),
.B2(n_62),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_117),
.Y(n_127)
);

OAI22x1_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_32),
.B1(n_27),
.B2(n_20),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_111),
.B1(n_112),
.B2(n_68),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_36),
.Y(n_103)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_106),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_25),
.B(n_22),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_109),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_63),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_22),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_75),
.C(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_69),
.B(n_22),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_12),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_70),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_72),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_123),
.B(n_128),
.Y(n_183)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_131),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_125),
.A2(n_151),
.B(n_102),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_121),
.C(n_108),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_87),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_93),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_148),
.B1(n_152),
.B2(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_24),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_139),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_141),
.B1(n_98),
.B2(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_108),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_146),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_86),
.B1(n_64),
.B2(n_20),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_113),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_100),
.A2(n_20),
.B1(n_27),
.B2(n_32),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_0),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_27),
.B1(n_32),
.B2(n_38),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_13),
.B(n_15),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_110),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_172),
.B(n_176),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_3),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_98),
.B(n_107),
.C(n_117),
.D(n_95),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_10),
.C(n_12),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_161),
.B1(n_167),
.B2(n_65),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_98),
.B1(n_106),
.B2(n_96),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_168),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_96),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_173),
.C(n_108),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_171),
.B1(n_175),
.B2(n_180),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_114),
.B1(n_27),
.B2(n_32),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_134),
.B(n_13),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_177),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_114),
.B1(n_73),
.B2(n_38),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_81),
.B(n_67),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_178),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_38),
.B1(n_73),
.B2(n_65),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_127),
.A2(n_0),
.B(n_1),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_127),
.B(n_11),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_127),
.B(n_146),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_136),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_105),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_135),
.B1(n_140),
.B2(n_149),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_126),
.A2(n_46),
.B(n_38),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_182),
.A2(n_184),
.B(n_2),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_132),
.A2(n_128),
.B(n_135),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_187),
.C(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_201),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_148),
.C(n_124),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_189),
.B(n_202),
.Y(n_233)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_191),
.Y(n_229)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_153),
.B1(n_170),
.B2(n_183),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_136),
.C(n_105),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_46),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_207),
.B1(n_174),
.B2(n_176),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_46),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_204),
.C(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_158),
.B(n_46),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_0),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_14),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_206),
.B(n_167),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_168),
.A2(n_165),
.B1(n_162),
.B2(n_171),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_9),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_4),
.B(n_5),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_210),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_186),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_187),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_227),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_221),
.C(n_228),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_224),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_153),
.C(n_182),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_192),
.Y(n_247)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_160),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_192),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_188),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_193),
.B1(n_191),
.B2(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_205),
.B(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_239),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_211),
.B(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_211),
.B(n_159),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_246),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_170),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_178),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_233),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_204),
.C(n_188),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_215),
.C(n_216),
.Y(n_252)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_251),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_184),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_215),
.C(n_221),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_255),
.B(n_248),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_228),
.C(n_233),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_219),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_259),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_197),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_190),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_220),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_265),
.A2(n_240),
.B(n_236),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_262),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_261),
.B(n_250),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_246),
.B(n_239),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_249),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_273),
.A2(n_274),
.B(n_276),
.Y(n_285)
);

A2O1A1O1Ixp25_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_237),
.B(n_244),
.C(n_251),
.D(n_243),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_259),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_237),
.B(n_243),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_284),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_253),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_286),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_234),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_256),
.B(n_202),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_252),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_266),
.B(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_293),
.C(n_7),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_242),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_292),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_281),
.B(n_242),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_285),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C1(n_10),
.C2(n_13),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_242),
.C(n_3),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_283),
.B(n_280),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_294),
.A2(n_296),
.B(n_287),
.Y(n_299)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_295),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_287),
.C(n_297),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_SL g301 ( 
.A1(n_300),
.A2(n_291),
.A3(n_298),
.B1(n_3),
.B2(n_14),
.C1(n_10),
.C2(n_7),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_14),
.Y(n_302)
);


endmodule