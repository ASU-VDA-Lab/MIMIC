module fake_jpeg_14027_n_484 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_484);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_484;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_9),
.B(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_64),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_33),
.A2(n_17),
.B(n_16),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_62),
.A2(n_56),
.B(n_41),
.C(n_25),
.Y(n_154)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_63),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_30),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_106),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_37),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g178 ( 
.A(n_72),
.Y(n_178)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_73),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_74),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_82),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_78),
.Y(n_193)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_81),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_18),
.B(n_17),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx2_ASAP7_75t_SL g148 ( 
.A(n_83),
.Y(n_148)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

BUFx2_ASAP7_75t_SL g192 ( 
.A(n_84),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_87),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_19),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_16),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_90),
.B(n_117),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_95),
.Y(n_149)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

INVx2_ASAP7_75t_R g95 ( 
.A(n_43),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_98),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_28),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_101),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_105),
.B(n_115),
.Y(n_184)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_108),
.Y(n_151)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_46),
.B(n_15),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_110),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_51),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_112),
.Y(n_183)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_10),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_118),
.Y(n_134)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_114),
.B(n_116),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_43),
.B(n_1),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_99),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_124),
.B(n_178),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_34),
.B1(n_29),
.B2(n_26),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_125),
.A2(n_157),
.B1(n_160),
.B2(n_170),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_63),
.A2(n_55),
.B1(n_26),
.B2(n_34),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_135),
.A2(n_139),
.B1(n_143),
.B2(n_145),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_55),
.B1(n_47),
.B2(n_26),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_136),
.B(n_162),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_81),
.A2(n_55),
.B1(n_103),
.B2(n_58),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_58),
.A2(n_32),
.B1(n_40),
.B2(n_45),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_83),
.A2(n_32),
.B1(n_40),
.B2(n_45),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_73),
.A2(n_52),
.B1(n_50),
.B2(n_44),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_146),
.A2(n_147),
.B1(n_171),
.B2(n_174),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_57),
.A2(n_52),
.B1(n_50),
.B2(n_44),
.Y(n_147)
);

OR2x2_ASAP7_75t_SL g235 ( 
.A(n_154),
.B(n_187),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_83),
.A2(n_40),
.B1(n_41),
.B2(n_56),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_155),
.A2(n_173),
.B1(n_188),
.B2(n_191),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_97),
.A2(n_25),
.B1(n_40),
.B2(n_22),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_102),
.A2(n_38),
.B1(n_36),
.B2(n_3),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_92),
.A2(n_38),
.B1(n_36),
.B2(n_3),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_59),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_164),
.A2(n_190),
.B1(n_136),
.B2(n_162),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_80),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_60),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_95),
.B(n_4),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_177),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_85),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_65),
.A2(n_6),
.B1(n_9),
.B2(n_74),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_86),
.B(n_93),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_107),
.A2(n_78),
.B1(n_75),
.B2(n_77),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_182),
.A2(n_170),
.B1(n_151),
.B2(n_193),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_104),
.A2(n_115),
.B1(n_105),
.B2(n_114),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_185),
.A2(n_164),
.B1(n_168),
.B2(n_137),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_120),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_85),
.A2(n_99),
.B1(n_66),
.B2(n_69),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_79),
.A2(n_106),
.B1(n_70),
.B2(n_67),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_119),
.A2(n_61),
.B1(n_64),
.B2(n_55),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_71),
.B(n_62),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_190),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_195),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_123),
.B(n_138),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_196),
.B(n_199),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_134),
.B(n_194),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_197),
.B(n_246),
.Y(n_265)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_177),
.A3(n_172),
.B1(n_163),
.B2(n_149),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_198),
.B(n_203),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_169),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_132),
.A2(n_175),
.B(n_183),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_200),
.B(n_204),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_202),
.A2(n_251),
.B1(n_168),
.B2(n_159),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_176),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_205),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_126),
.B(n_127),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_206),
.B(n_227),
.Y(n_290)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_131),
.Y(n_207)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_210),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_211),
.B(n_229),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_212),
.Y(n_282)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_215),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_221),
.Y(n_262)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_218),
.Y(n_298)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_129),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_220),
.Y(n_303)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_121),
.Y(n_221)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_222),
.Y(n_272)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_223),
.B(n_226),
.Y(n_307)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_129),
.Y(n_224)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_126),
.B(n_127),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_122),
.B(n_153),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_228),
.B(n_241),
.Y(n_293)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_141),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_230),
.A2(n_207),
.B1(n_205),
.B2(n_231),
.Y(n_301)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_231),
.Y(n_287)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_140),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_232),
.B(n_233),
.Y(n_305)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_159),
.B(n_225),
.Y(n_261)
);

NOR2x1_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_243),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_182),
.A2(n_190),
.B1(n_158),
.B2(n_133),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_236),
.A2(n_239),
.B1(n_247),
.B2(n_250),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_141),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_184),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_235),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_133),
.A2(n_158),
.B1(n_184),
.B2(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_142),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_122),
.B(n_153),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_122),
.B(n_153),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_242),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_151),
.Y(n_243)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_128),
.Y(n_245)
);

BUFx8_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_120),
.B(n_189),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_144),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_151),
.B(n_120),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_161),
.Y(n_250)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_128),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_137),
.A2(n_148),
.B(n_133),
.C(n_158),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_161),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_179),
.B(n_152),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_179),
.B(n_152),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_193),
.B(n_166),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_258),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_166),
.B(n_144),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_260),
.A2(n_296),
.B1(n_269),
.B2(n_280),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_261),
.B(n_265),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_208),
.A2(n_236),
.B1(n_217),
.B2(n_201),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_263),
.A2(n_301),
.B1(n_304),
.B2(n_282),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_264),
.A2(n_270),
.B(n_275),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_202),
.A2(n_208),
.B1(n_213),
.B2(n_246),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_268),
.A2(n_276),
.B1(n_280),
.B2(n_294),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_217),
.B(n_239),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_216),
.A2(n_244),
.B1(n_201),
.B2(n_238),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_252),
.B1(n_198),
.B2(n_197),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_220),
.A2(n_224),
.B1(n_229),
.B2(n_247),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_212),
.B(n_253),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_286),
.B(n_298),
.C(n_291),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_218),
.A2(n_219),
.B(n_209),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_291),
.A2(n_262),
.B(n_307),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g292 ( 
.A(n_221),
.B(n_226),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_286),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_237),
.A2(n_232),
.B1(n_223),
.B2(n_222),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_305),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_309),
.B(n_326),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_313),
.Y(n_349)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_288),
.Y(n_311)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_311),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_312),
.A2(n_333),
.B(n_334),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_265),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_275),
.A2(n_260),
.B1(n_270),
.B2(n_274),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_315),
.B1(n_323),
.B2(n_328),
.Y(n_345)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_284),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_317),
.B(n_319),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_324),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_259),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_259),
.B(n_297),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_320),
.B(n_321),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_273),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_293),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_331),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_271),
.A2(n_263),
.B1(n_264),
.B2(n_297),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_271),
.A2(n_262),
.B1(n_279),
.B2(n_292),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_306),
.B(n_281),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_327),
.A2(n_344),
.B(n_287),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_279),
.A2(n_262),
.B1(n_277),
.B2(n_266),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_302),
.B(n_277),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_298),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_307),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_332),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_304),
.A2(n_266),
.B1(n_294),
.B2(n_283),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

INVx3_ASAP7_75t_SL g348 ( 
.A(n_335),
.Y(n_348)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_267),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_339),
.A2(n_343),
.B1(n_299),
.B2(n_300),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_307),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_340),
.Y(n_356)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_341),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_272),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_342),
.Y(n_367)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_272),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_346),
.A2(n_344),
.B(n_342),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_287),
.C(n_303),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_360),
.C(n_371),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_325),
.A2(n_299),
.B(n_300),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_359),
.A2(n_369),
.B(n_326),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_299),
.C(n_300),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_366),
.A2(n_372),
.B1(n_374),
.B2(n_334),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_325),
.A2(n_333),
.B(n_327),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_323),
.B(n_320),
.C(n_319),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_314),
.B1(n_324),
.B2(n_317),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_332),
.A2(n_340),
.B1(n_318),
.B2(n_309),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_364),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_382),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_322),
.C(n_331),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_390),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_377),
.A2(n_380),
.B(n_356),
.Y(n_400)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_347),
.Y(n_378)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_381),
.A2(n_385),
.B1(n_387),
.B2(n_391),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_367),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_329),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_386),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_308),
.Y(n_384)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_372),
.A2(n_321),
.B1(n_311),
.B2(n_336),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_364),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_372),
.A2(n_337),
.B1(n_316),
.B2(n_341),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_338),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_388),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_343),
.C(n_330),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_345),
.A2(n_335),
.B1(n_341),
.B2(n_374),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_374),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_392),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_357),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_354),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_355),
.B(n_356),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_394),
.A2(n_398),
.B1(n_353),
.B2(n_365),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_370),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_397),
.Y(n_407)
);

INVx8_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_396),
.Y(n_406)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_392),
.A2(n_345),
.B1(n_361),
.B2(n_349),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_399),
.A2(n_412),
.B1(n_363),
.B2(n_387),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_377),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_403),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_381),
.A2(n_363),
.B1(n_349),
.B2(n_368),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_405),
.A2(n_413),
.B1(n_384),
.B2(n_354),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_357),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_410),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_393),
.B(n_371),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_380),
.A2(n_345),
.B1(n_359),
.B2(n_366),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_391),
.A2(n_363),
.B1(n_368),
.B2(n_370),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_375),
.A2(n_395),
.B1(n_383),
.B2(n_366),
.Y(n_414)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_414),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_419),
.B(n_389),
.C(n_390),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_389),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_426),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_411),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_424),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_408),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_430),
.B1(n_417),
.B2(n_415),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_389),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_394),
.Y(n_427)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_427),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_390),
.C(n_376),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_433),
.C(n_404),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_402),
.A2(n_385),
.B1(n_363),
.B2(n_388),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_431),
.A2(n_401),
.B1(n_418),
.B2(n_378),
.Y(n_449)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_435),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_360),
.C(n_362),
.Y(n_433)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_407),
.A2(n_382),
.B(n_360),
.C(n_397),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_416),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_436),
.B(n_415),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_448),
.C(n_429),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_405),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_440),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_425),
.A2(n_412),
.B1(n_417),
.B2(n_399),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_442),
.A2(n_434),
.B1(n_424),
.B2(n_423),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_444),
.B(n_422),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_400),
.B(n_413),
.Y(n_445)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_445),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_446),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_402),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_449),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_451),
.B(n_443),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_452),
.B(n_458),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_456),
.A2(n_438),
.B1(n_433),
.B2(n_440),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_435),
.Y(n_457)
);

OAI21x1_ASAP7_75t_SL g461 ( 
.A1(n_457),
.A2(n_459),
.B(n_439),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_444),
.B(n_430),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_401),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_350),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_448),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_462),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_461),
.A2(n_463),
.B1(n_465),
.B2(n_466),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_454),
.A2(n_406),
.B1(n_379),
.B2(n_358),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_450),
.C(n_428),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_455),
.A2(n_406),
.B1(n_358),
.B2(n_396),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_443),
.C(n_437),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_468),
.B(n_473),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_467),
.B(n_451),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_470),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_462),
.B(n_457),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_465),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_475),
.B(n_476),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_472),
.A2(n_450),
.B(n_463),
.Y(n_476)
);

XOR2x1_ASAP7_75t_SL g478 ( 
.A(n_474),
.B(n_468),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_478),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_477),
.A2(n_396),
.B1(n_373),
.B2(n_351),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_480),
.A2(n_351),
.B(n_352),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_481),
.B(n_479),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_483),
.A2(n_482),
.B(n_428),
.Y(n_484)
);


endmodule