module fake_ariane_20_n_14705 (n_913, n_1681, n_2163, n_1486, n_1507, n_1938, n_589, n_2484, n_1174, n_2346, n_1469, n_691, n_1353, n_1355, n_2131, n_2500, n_2509, n_423, n_1383, n_2182, n_603, n_373, n_2135, n_2334, n_1250, n_2030, n_1169, n_789, n_850, n_1916, n_610, n_245, n_1713, n_96, n_319, n_49, n_1436, n_2407, n_690, n_416, n_1109, n_1430, n_2537, n_525, n_187, n_2002, n_1463, n_2243, n_1238, n_2011, n_1515, n_817, n_1837, n_924, n_781, n_2013, n_1566, n_189, n_717, n_72, n_2006, n_952, n_864, n_2446, n_1096, n_1379, n_2436, n_57, n_2376, n_2367, n_1706, n_2207, n_2461, n_117, n_524, n_1214, n_634, n_1839, n_1246, n_1138, n_214, n_2042, n_2123, n_1853, n_764, n_1503, n_2238, n_2529, n_2374, n_462, n_1196, n_1181, n_32, n_1999, n_410, n_2380, n_1187, n_1131, n_1225, n_737, n_137, n_1298, n_1745, n_1366, n_232, n_52, n_2084, n_568, n_2278, n_1088, n_77, n_1424, n_766, n_1835, n_1457, n_377, n_2482, n_1682, n_1836, n_520, n_870, n_2547, n_1453, n_279, n_945, n_958, n_2554, n_2248, n_813, n_419, n_1985, n_2288, n_146, n_270, n_338, n_995, n_285, n_1909, n_2156, n_1184, n_1961, n_202, n_1535, n_500, n_665, n_754, n_903, n_871, n_2323, n_1073, n_239, n_402, n_1979, n_1277, n_2107, n_1746, n_54, n_829, n_1761, n_1062, n_339, n_738, n_1690, n_2221, n_672, n_740, n_1283, n_167, n_2317, n_1974, n_1736, n_1018, n_2342, n_2200, n_69, n_259, n_2442, n_953, n_1364, n_2390, n_143, n_1888, n_1224, n_2109, n_1425, n_625, n_557, n_2322, n_1107, n_1688, n_989, n_242, n_645, n_1944, n_331, n_559, n_2233, n_2370, n_267, n_495, n_1988, n_350, n_381, n_795, n_721, n_1084, n_1718, n_1276, n_1936, n_2149, n_2277, n_200, n_1428, n_1284, n_1241, n_821, n_561, n_770, n_1514, n_2539, n_1528, n_507, n_486, n_901, n_569, n_2078, n_1145, n_971, n_2359, n_2201, n_787, n_1650, n_31, n_1519, n_1195, n_2049, n_1522, n_518, n_1207, n_222, n_786, n_1404, n_868, n_2232, n_1847, n_2458, n_1542, n_1314, n_1512, n_2227, n_2301, n_1539, n_884, n_1851, n_2162, n_1415, n_1034, n_1652, n_2192, n_1676, n_1085, n_277, n_1636, n_432, n_293, n_823, n_1900, n_620, n_93, n_1074, n_859, n_1765, n_108, n_1889, n_587, n_1977, n_693, n_863, n_303, n_1254, n_929, n_2433, n_206, n_352, n_899, n_1703, n_2332, n_2391, n_611, n_1295, n_2060, n_1850, n_238, n_365, n_2004, n_1013, n_1495, n_1637, n_136, n_334, n_2427, n_192, n_661, n_2098, n_1751, n_300, n_533, n_1917, n_2456, n_104, n_1924, n_438, n_1560, n_1654, n_2341, n_1548, n_16, n_1811, n_2045, n_440, n_273, n_1396, n_1230, n_612, n_333, n_1840, n_376, n_512, n_1597, n_1771, n_1544, n_579, n_844, n_1012, n_1267, n_2061, n_2094, n_2512, n_1354, n_1790, n_149, n_1213, n_2382, n_237, n_2043, n_780, n_2349, n_1918, n_1021, n_1443, n_491, n_1465, n_1949, n_1595, n_1142, n_1140, n_705, n_570, n_260, n_942, n_1437, n_7, n_2077, n_1378, n_461, n_1121, n_1416, n_209, n_490, n_1461, n_17, n_1391, n_1947, n_225, n_1599, n_1876, n_1006, n_1830, n_575, n_546, n_503, n_2527, n_1112, n_700, n_1159, n_772, n_1216, n_1245, n_1669, n_1675, n_2466, n_676, n_42, n_2038, n_2263, n_2116, n_2271, n_2145, n_2326, n_1838, n_1594, n_680, n_1935, n_287, n_1716, n_302, n_1872, n_380, n_1585, n_2281, n_1432, n_94, n_2245, n_4, n_249, n_1108, n_355, n_212, n_65, n_123, n_444, n_851, n_1590, n_1351, n_2216, n_1274, n_257, n_2426, n_652, n_1819, n_475, n_135, n_947, n_2134, n_930, n_1260, n_1179, n_468, n_102, n_182, n_696, n_1442, n_482, n_798, n_577, n_1833, n_407, n_1691, n_27, n_916, n_1386, n_912, n_1884, n_460, n_1555, n_1842, n_2499, n_2549, n_366, n_762, n_1253, n_1468, n_1661, n_555, n_804, n_1656, n_1382, n_966, n_992, n_955, n_1182, n_794, n_78, n_2166, n_1692, n_1562, n_514, n_418, n_2185, n_2398, n_1376, n_513, n_288, n_179, n_1292, n_1178, n_1972, n_2015, n_1435, n_1750, n_1026, n_1506, n_1610, n_2202, n_2072, n_306, n_2415, n_92, n_203, n_436, n_150, n_324, n_2087, n_669, n_931, n_1491, n_619, n_337, n_437, n_111, n_21, n_274, n_967, n_1083, n_2161, n_1418, n_746, n_1357, n_292, n_1079, n_1787, n_2462, n_1389, n_2155, n_615, n_1139, n_76, n_2439, n_517, n_1312, n_1717, n_0, n_1812, n_824, n_428, n_159, n_2172, n_892, n_1880, n_959, n_30, n_2365, n_2257, n_1399, n_1101, n_1567, n_1343, n_563, n_2219, n_1855, n_2100, n_2333, n_144, n_990, n_1623, n_1903, n_867, n_2147, n_2435, n_1226, n_2224, n_944, n_749, n_1932, n_1780, n_1970, n_1920, n_2083, n_815, n_542, n_2167, n_2293, n_1340, n_470, n_1240, n_1087, n_2400, n_632, n_477, n_650, n_2388, n_425, n_2273, n_1433, n_1911, n_1825, n_1908, n_1155, n_1071, n_712, n_976, n_909, n_1392, n_767, n_1832, n_1841, n_1680, n_2066, n_2302, n_964, n_1627, n_2220, n_382, n_489, n_2294, n_80, n_2274, n_251, n_974, n_506, n_1731, n_799, n_1147, n_2378, n_397, n_2467, n_471, n_351, n_965, n_1914, n_155, n_2253, n_934, n_2213, n_1447, n_2363, n_1220, n_356, n_2019, n_698, n_2130, n_1674, n_2021, n_2025, n_2160, n_1992, n_124, n_307, n_1209, n_1020, n_1563, n_646, n_2507, n_2142, n_1633, n_34, n_404, n_172, n_1913, n_2069, n_2495, n_1058, n_2328, n_347, n_2434, n_1042, n_183, n_1234, n_2311, n_479, n_1578, n_2261, n_1455, n_2287, n_299, n_836, n_2223, n_1279, n_2473, n_2144, n_2511, n_564, n_133, n_66, n_205, n_1029, n_1247, n_760, n_522, n_2438, n_1568, n_20, n_1483, n_1363, n_367, n_1111, n_970, n_1689, n_2535, n_713, n_1255, n_1646, n_598, n_345, n_2262, n_1237, n_927, n_261, n_1095, n_1728, n_2335, n_370, n_706, n_2120, n_286, n_1401, n_1419, n_1531, n_776, n_424, n_2041, n_2113, n_1933, n_1651, n_85, n_130, n_1387, n_466, n_1263, n_346, n_1817, n_2404, n_2168, n_348, n_552, n_2312, n_670, n_1826, n_379, n_138, n_162, n_264, n_2483, n_441, n_1951, n_2490, n_1032, n_1217, n_1496, n_637, n_1592, n_73, n_327, n_1259, n_1177, n_1231, n_2132, n_980, n_1618, n_1869, n_1743, n_905, n_207, n_720, n_926, n_41, n_1943, n_2296, n_194, n_1802, n_2178, n_2112, n_1163, n_186, n_1795, n_1384, n_2237, n_145, n_2146, n_1868, n_59, n_1501, n_2241, n_2373, n_1173, n_2350, n_1068, n_1198, n_2531, n_1570, n_2099, n_487, n_1518, n_1456, n_90, n_1879, n_1886, n_1648, n_2187, n_1413, n_2481, n_2129, n_855, n_2327, n_158, n_808, n_1365, n_2476, n_553, n_2059, n_2437, n_1439, n_814, n_578, n_2074, n_1665, n_1287, n_405, n_1611, n_2122, n_120, n_2399, n_320, n_1414, n_1134, n_2067, n_1484, n_1901, n_647, n_2055, n_2027, n_1423, n_2117, n_481, n_600, n_1053, n_1609, n_1939, n_2308, n_2242, n_1906, n_529, n_1899, n_2195, n_502, n_2194, n_218, n_1467, n_247, n_1828, n_2159, n_1798, n_1304, n_1608, n_1744, n_2267, n_1105, n_547, n_439, n_604, n_677, n_478, n_703, n_1349, n_1709, n_1061, n_2102, n_326, n_681, n_227, n_874, n_2286, n_2023, n_1278, n_707, n_11, n_129, n_126, n_983, n_590, n_699, n_727, n_301, n_1726, n_2075, n_2523, n_1945, n_545, n_1015, n_2418, n_1377, n_1162, n_536, n_1614, n_2031, n_2496, n_2118, n_325, n_1740, n_1602, n_688, n_636, n_427, n_1098, n_1490, n_2338, n_442, n_777, n_1553, n_1080, n_920, n_1760, n_1086, n_1092, n_2225, n_986, n_1104, n_1963, n_729, n_887, n_2057, n_2218, n_1122, n_1205, n_1408, n_163, n_1693, n_2125, n_1132, n_390, n_1156, n_501, n_2184, n_314, n_1823, n_1120, n_1202, n_627, n_2254, n_1188, n_1498, n_1371, n_2033, n_233, n_957, n_388, n_1402, n_1242, n_1607, n_1489, n_1218, n_2217, n_221, n_321, n_86, n_2226, n_1586, n_861, n_1543, n_1431, n_877, n_1119, n_1863, n_1763, n_1666, n_1500, n_616, n_2214, n_1055, n_1395, n_1346, n_2256, n_1189, n_1089, n_281, n_1859, n_262, n_1502, n_1523, n_2190, n_1478, n_1883, n_2516, n_1969, n_735, n_297, n_1005, n_527, n_2379, n_46, n_84, n_1294, n_1667, n_845, n_888, n_2300, n_1649, n_2452, n_1677, n_2470, n_1927, n_1297, n_178, n_551, n_417, n_1708, n_70, n_343, n_1222, n_2284, n_1844, n_2283, n_582, n_2526, n_1957, n_1953, n_755, n_1097, n_1219, n_1711, n_710, n_1919, n_534, n_1791, n_2508, n_2124, n_1894, n_1460, n_1239, n_278, n_2266, n_2449, n_560, n_890, n_842, n_148, n_1898, n_451, n_745, n_1741, n_1572, n_1907, n_1793, n_61, n_742, n_1081, n_1373, n_1975, n_1388, n_1266, n_1540, n_1719, n_2119, n_769, n_1797, n_2366, n_2493, n_13, n_1753, n_1990, n_1372, n_476, n_832, n_55, n_535, n_744, n_1895, n_2474, n_982, n_1800, n_915, n_215, n_1075, n_2008, n_454, n_298, n_1331, n_1890, n_1529, n_1227, n_2127, n_655, n_1734, n_1860, n_403, n_2460, n_1007, n_1580, n_1319, n_657, n_837, n_812, n_2448, n_2211, n_2292, n_2480, n_606, n_951, n_862, n_1700, n_659, n_1332, n_2306, n_509, n_1854, n_666, n_1747, n_2071, n_2424, n_430, n_1206, n_1729, n_722, n_1508, n_2414, n_2082, n_1532, n_1171, n_1030, n_785, n_2389, n_1309, n_999, n_2280, n_1766, n_1338, n_1342, n_456, n_1867, n_852, n_1394, n_704, n_1060, n_1044, n_1714, n_521, n_2140, n_873, n_1301, n_1748, n_2157, n_1966, n_1243, n_2171, n_2468, n_1400, n_342, n_2035, n_1466, n_1513, n_1527, n_358, n_1783, n_608, n_2494, n_1538, n_2457, n_2128, n_1037, n_1329, n_317, n_1993, n_1545, n_134, n_1257, n_1480, n_1954, n_1668, n_1878, n_2540, n_1605, n_1078, n_266, n_2486, n_1897, n_157, n_2520, n_2137, n_1161, n_2489, n_811, n_624, n_791, n_876, n_618, n_1191, n_2492, n_736, n_1025, n_1215, n_241, n_1449, n_2337, n_2265, n_687, n_797, n_2026, n_1786, n_480, n_1327, n_1475, n_211, n_642, n_1804, n_2106, n_97, n_408, n_1406, n_595, n_1405, n_602, n_2272, n_1757, n_592, n_1499, n_854, n_1318, n_2091, n_393, n_1632, n_1769, n_474, n_1929, n_1950, n_2264, n_805, n_2032, n_2090, n_295, n_1658, n_190, n_2249, n_1072, n_695, n_1526, n_1305, n_64, n_180, n_730, n_386, n_1596, n_2348, n_1281, n_516, n_2364, n_1997, n_1137, n_1873, n_1258, n_197, n_640, n_463, n_1476, n_1524, n_1733, n_1856, n_2016, n_943, n_1118, n_678, n_651, n_1874, n_1293, n_961, n_469, n_1046, n_1807, n_726, n_1123, n_1657, n_878, n_1784, n_771, n_1321, n_752, n_2307, n_71, n_1488, n_985, n_421, n_1330, n_906, n_1180, n_1697, n_2295, n_283, n_806, n_1984, n_1350, n_1556, n_649, n_1561, n_2412, n_374, n_1352, n_2405, n_1824, n_643, n_1492, n_226, n_2383, n_1441, n_1822, n_682, n_36, n_1616, n_2416, n_819, n_2386, n_1971, n_586, n_1324, n_1429, n_2064, n_2353, n_2528, n_1778, n_1776, n_686, n_605, n_1154, n_584, n_1557, n_1759, n_1829, n_2325, n_1130, n_1450, n_349, n_756, n_2022, n_1016, n_2298, n_1149, n_1505, n_2408, n_2320, n_979, n_2329, n_1642, n_2417, n_2, n_2525, n_1815, n_897, n_2546, n_949, n_2454, n_1493, n_515, n_807, n_891, n_885, n_1659, n_2354, n_198, n_1864, n_1887, n_1208, n_1987, n_396, n_2368, n_802, n_23, n_1151, n_554, n_960, n_2352, n_2502, n_1256, n_87, n_714, n_2170, n_790, n_2244, n_2143, n_2393, n_354, n_140, n_725, n_2377, n_1577, n_151, n_1448, n_2198, n_28, n_1009, n_230, n_1133, n_154, n_883, n_142, n_473, n_1852, n_801, n_1286, n_818, n_1685, n_779, n_2410, n_2314, n_2477, n_2279, n_594, n_2222, n_1995, n_1877, n_1397, n_35, n_1052, n_272, n_1333, n_1306, n_1849, n_2076, n_2133, n_2203, n_833, n_1426, n_2250, n_2497, n_2247, n_2230, n_879, n_1117, n_38, n_422, n_1269, n_1303, n_1547, n_1438, n_1541, n_597, n_75, n_2001, n_1047, n_95, n_2506, n_1472, n_2413, n_1593, n_1050, n_566, n_2158, n_2285, n_152, n_169, n_106, n_1201, n_1288, n_173, n_858, n_1185, n_2475, n_2173, n_335, n_1035, n_1143, n_344, n_2070, n_2136, n_426, n_433, n_398, n_62, n_210, n_1090, n_2403, n_1367, n_2044, n_166, n_253, n_928, n_1153, n_271, n_465, n_825, n_1103, n_732, n_1565, n_1192, n_128, n_224, n_82, n_894, n_1380, n_1624, n_1801, n_420, n_1291, n_562, n_2020, n_748, n_2310, n_510, n_1045, n_256, n_1160, n_1882, n_1976, n_1023, n_1881, n_988, n_330, n_914, n_400, n_689, n_1116, n_282, n_328, n_368, n_1958, n_467, n_1511, n_2177, n_1422, n_1965, n_644, n_1197, n_276, n_497, n_1165, n_1641, n_168, n_81, n_538, n_1517, n_2036, n_576, n_843, n_511, n_455, n_429, n_588, n_638, n_2003, n_2533, n_2210, n_1307, n_1128, n_2053, n_1671, n_1417, n_1048, n_2343, n_775, n_667, n_2419, n_1049, n_2330, n_14, n_869, n_141, n_846, n_1398, n_1921, n_2450, n_2411, n_1356, n_1341, n_2234, n_2309, n_1504, n_1955, n_2110, n_2431, n_1773, n_1440, n_1370, n_1603, n_305, n_312, n_56, n_60, n_728, n_413, n_2401, n_715, n_889, n_1066, n_1549, n_2331, n_935, n_2478, n_685, n_911, n_361, n_89, n_623, n_1712, n_1403, n_1065, n_453, n_1534, n_1948, n_74, n_810, n_19, n_40, n_1290, n_181, n_1959, n_617, n_2396, n_543, n_1362, n_1559, n_2121, n_236, n_601, n_683, n_565, n_628, n_1300, n_1960, n_2068, n_743, n_1194, n_1647, n_1546, n_1420, n_2553, n_907, n_1454, n_660, n_464, n_2459, n_962, n_941, n_1210, n_847, n_747, n_1622, n_1135, n_918, n_1968, n_107, n_1885, n_639, n_452, n_673, n_2196, n_1038, n_2371, n_1978, n_414, n_571, n_1521, n_1694, n_1940, n_6, n_284, n_593, n_1695, n_1164, n_37, n_58, n_2313, n_609, n_1193, n_1345, n_613, n_1022, n_1336, n_1033, n_1774, n_409, n_171, n_519, n_384, n_1166, n_1056, n_2007, n_526, n_1994, n_1767, n_1040, n_674, n_1158, n_316, n_125, n_1973, n_1444, n_1803, n_820, n_1749, n_43, n_872, n_1653, n_254, n_2303, n_1157, n_1584, n_234, n_848, n_1664, n_280, n_629, n_1739, n_161, n_1814, n_532, n_2154, n_2441, n_2236, n_1789, n_763, n_1986, n_2174, n_99, n_540, n_216, n_692, n_5, n_2054, n_1857, n_2315, n_984, n_1687, n_2073, n_223, n_2150, n_1552, n_750, n_834, n_1612, n_2498, n_800, n_2046, n_1816, n_1910, n_1756, n_1606, n_2189, n_395, n_621, n_1587, n_213, n_2093, n_2340, n_2018, n_1772, n_67, n_2444, n_1014, n_724, n_2204, n_1427, n_1481, n_2040, n_493, n_1311, n_2199, n_1956, n_1589, n_114, n_2151, n_1100, n_585, n_875, n_1617, n_2455, n_827, n_2231, n_697, n_622, n_1626, n_1962, n_1335, n_1715, n_296, n_2305, n_880, n_793, n_2114, n_1175, n_2289, n_132, n_2530, n_2299, n_751, n_1027, n_1070, n_2406, n_1621, n_739, n_1485, n_1028, n_1221, n_530, n_1785, n_792, n_1262, n_1942, n_2180, n_580, n_1579, n_494, n_2181, n_434, n_2014, n_975, n_229, n_394, n_923, n_1645, n_1124, n_1381, n_1494, n_932, n_1893, n_1183, n_1326, n_2276, n_1805, n_2282, n_981, n_2141, n_1110, n_1758, n_2503, n_2270, n_243, n_2443, n_1407, n_185, n_2465, n_1204, n_1554, n_994, n_2428, n_1360, n_973, n_268, n_972, n_2251, n_164, n_184, n_856, n_1248, n_1176, n_1564, n_2010, n_1054, n_508, n_118, n_121, n_1679, n_2126, n_1952, n_2425, n_2394, n_1858, n_353, n_1678, n_1482, n_1361, n_2356, n_1601, n_1057, n_191, n_2487, n_1834, n_978, n_1011, n_1520, n_2534, n_2488, n_1509, n_828, n_322, n_1411, n_1359, n_558, n_1721, n_116, n_39, n_653, n_1445, n_1317, n_2050, n_2197, n_783, n_2550, n_556, n_1127, n_170, n_1536, n_1471, n_2385, n_160, n_119, n_2387, n_1008, n_332, n_581, n_294, n_1024, n_830, n_176, n_2291, n_1980, n_2518, n_987, n_936, n_2510, n_1620, n_2501, n_2542, n_1385, n_1525, n_1998, n_2165, n_541, n_499, n_1775, n_788, n_12, n_908, n_1036, n_2169, n_341, n_1270, n_109, n_1167, n_1272, n_549, n_591, n_969, n_2028, n_919, n_1663, n_50, n_2092, n_2175, n_1625, n_2086, n_1926, n_2402, n_318, n_1458, n_103, n_244, n_679, n_1630, n_220, n_663, n_1720, n_2409, n_443, n_2176, n_1412, n_1738, n_1550, n_528, n_1358, n_1200, n_387, n_406, n_826, n_139, n_2453, n_2344, n_1922, n_1735, n_1788, n_391, n_940, n_2392, n_1537, n_2138, n_2065, n_2543, n_2321, n_1077, n_607, n_956, n_445, n_1930, n_765, n_1809, n_1843, n_1904, n_122, n_2000, n_1268, n_385, n_2395, n_917, n_1271, n_372, n_2096, n_2440, n_2186, n_15, n_1530, n_2215, n_631, n_399, n_1170, n_2258, n_1261, n_2471, n_702, n_857, n_898, n_363, n_968, n_1067, n_1235, n_1323, n_2375, n_1462, n_1937, n_2012, n_1064, n_633, n_900, n_1446, n_1282, n_1701, n_1093, n_1551, n_2039, n_1755, n_1285, n_193, n_733, n_761, n_2212, n_731, n_336, n_1813, n_315, n_2268, n_311, n_1452, n_1573, n_8, n_668, n_758, n_2252, n_2111, n_2420, n_1996, n_1106, n_2009, n_47, n_153, n_18, n_648, n_784, n_269, n_816, n_1322, n_1473, n_835, n_446, n_1076, n_2024, n_1348, n_753, n_2445, n_1770, n_701, n_1003, n_2469, n_1125, n_2103, n_2358, n_1710, n_1865, n_2522, n_2463, n_309, n_1344, n_115, n_2355, n_1390, n_401, n_485, n_1792, n_504, n_2062, n_483, n_435, n_1141, n_1629, n_291, n_1640, n_822, n_1094, n_840, n_1459, n_2153, n_2324, n_1510, n_2505, n_2139, n_1099, n_839, n_79, n_1754, n_3, n_759, n_567, n_2397, n_91, n_2521, n_240, n_369, n_1727, n_2235, n_44, n_1991, n_1575, n_1848, n_1892, n_1172, n_614, n_1212, n_831, n_778, n_48, n_1619, n_2351, n_188, n_2260, n_323, n_550, n_1315, n_1660, n_1902, n_997, n_635, n_2206, n_2541, n_694, n_1643, n_1320, n_1113, n_2347, n_248, n_1152, n_2447, n_2034, n_1845, n_2538, n_1934, n_2101, n_921, n_2362, n_1615, n_1236, n_228, n_2104, n_1265, n_1576, n_2105, n_1470, n_671, n_1533, n_1806, n_2372, n_2552, n_1, n_1409, n_1148, n_1588, n_1684, n_1673, n_2422, n_1334, n_654, n_2290, n_2088, n_1275, n_488, n_904, n_505, n_88, n_2005, n_2048, n_1696, n_498, n_1875, n_1059, n_684, n_2429, n_2108, n_1039, n_2246, n_539, n_1150, n_977, n_449, n_2339, n_392, n_1628, n_1289, n_1831, n_2532, n_2191, n_1497, n_1866, n_2472, n_2056, n_459, n_1136, n_2515, n_1782, n_458, n_1190, n_1600, n_1144, n_383, n_838, n_1558, n_1941, n_1316, n_175, n_2519, n_950, n_1017, n_711, n_734, n_1915, n_2360, n_723, n_1393, n_2240, n_658, n_630, n_1369, n_53, n_362, n_310, n_1781, n_709, n_2544, n_24, n_809, n_2085, n_2432, n_1686, n_1964, n_235, n_881, n_1019, n_1477, n_1777, n_2188, n_1982, n_2097, n_662, n_641, n_2430, n_2504, n_910, n_290, n_741, n_939, n_1410, n_2297, n_371, n_199, n_217, n_1114, n_1325, n_1742, n_708, n_308, n_1223, n_2545, n_201, n_1768, n_2513, n_2193, n_2369, n_572, n_1199, n_865, n_10, n_1273, n_1983, n_1041, n_2451, n_2115, n_993, n_1862, n_948, n_2017, n_922, n_1004, n_1810, n_448, n_1347, n_860, n_1043, n_255, n_450, n_1923, n_1764, n_896, n_1737, n_1479, n_1613, n_902, n_1031, n_1723, n_1638, n_853, n_716, n_1571, n_1698, n_196, n_1337, n_774, n_1946, n_2148, n_933, n_1779, n_596, n_954, n_2051, n_1168, n_1821, n_219, n_1310, n_231, n_656, n_492, n_574, n_252, n_664, n_1591, n_1229, n_1683, n_2548, n_68, n_1896, n_2164, n_1732, n_415, n_2381, n_1967, n_2384, n_2179, n_63, n_1280, n_544, n_1516, n_1186, n_1705, n_599, n_768, n_1091, n_2052, n_2485, n_537, n_1063, n_25, n_991, n_2183, n_2205, n_83, n_2275, n_389, n_1724, n_1670, n_1707, n_1799, n_2080, n_2058, n_1126, n_2357, n_2029, n_195, n_1846, n_1912, n_938, n_1891, n_1328, n_895, n_110, n_304, n_1639, n_583, n_2209, n_2421, n_1302, n_1000, n_313, n_626, n_378, n_1581, n_1928, n_98, n_946, n_757, n_2047, n_375, n_113, n_1655, n_1818, n_33, n_1146, n_1634, n_1203, n_998, n_1699, n_1598, n_2269, n_472, n_937, n_1474, n_2081, n_2536, n_2524, n_265, n_1583, n_1604, n_208, n_1631, n_1702, n_156, n_174, n_275, n_100, n_1794, n_1375, n_147, n_204, n_1232, n_996, n_1211, n_1368, n_963, n_1264, n_51, n_1082, n_1725, n_496, n_2318, n_1827, n_866, n_26, n_246, n_925, n_1752, n_1313, n_1001, n_1722, n_2361, n_1115, n_2229, n_1339, n_1002, n_1644, n_105, n_1051, n_2551, n_719, n_131, n_263, n_1102, n_360, n_2255, n_1129, n_1252, n_2239, n_250, n_1464, n_1296, n_773, n_2316, n_165, n_2464, n_1010, n_882, n_2304, n_1249, n_101, n_803, n_1871, n_2514, n_329, n_718, n_1434, n_340, n_1905, n_1569, n_289, n_9, n_112, n_45, n_548, n_2336, n_523, n_1662, n_457, n_1299, n_1870, n_177, n_2063, n_1925, n_782, n_364, n_258, n_431, n_2491, n_1861, n_2079, n_1228, n_2319, n_2152, n_2517, n_1931, n_1244, n_1796, n_411, n_484, n_2259, n_849, n_2095, n_22, n_1820, n_29, n_357, n_412, n_1251, n_1989, n_447, n_1421, n_2208, n_2423, n_1762, n_1233, n_1808, n_1574, n_1672, n_2228, n_1635, n_1704, n_893, n_1582, n_841, n_2479, n_886, n_1069, n_1981, n_2037, n_359, n_1308, n_573, n_796, n_127, n_531, n_2345, n_1730, n_1374, n_1451, n_2089, n_1487, n_675, n_14705);

input n_913;
input n_1681;
input n_2163;
input n_1486;
input n_1507;
input n_1938;
input n_589;
input n_2484;
input n_1174;
input n_2346;
input n_1469;
input n_691;
input n_1353;
input n_1355;
input n_2131;
input n_2500;
input n_2509;
input n_423;
input n_1383;
input n_2182;
input n_603;
input n_373;
input n_2135;
input n_2334;
input n_1250;
input n_2030;
input n_1169;
input n_789;
input n_850;
input n_1916;
input n_610;
input n_245;
input n_1713;
input n_96;
input n_319;
input n_49;
input n_1436;
input n_2407;
input n_690;
input n_416;
input n_1109;
input n_1430;
input n_2537;
input n_525;
input n_187;
input n_2002;
input n_1463;
input n_2243;
input n_1238;
input n_2011;
input n_1515;
input n_817;
input n_1837;
input n_924;
input n_781;
input n_2013;
input n_1566;
input n_189;
input n_717;
input n_72;
input n_2006;
input n_952;
input n_864;
input n_2446;
input n_1096;
input n_1379;
input n_2436;
input n_57;
input n_2376;
input n_2367;
input n_1706;
input n_2207;
input n_2461;
input n_117;
input n_524;
input n_1214;
input n_634;
input n_1839;
input n_1246;
input n_1138;
input n_214;
input n_2042;
input n_2123;
input n_1853;
input n_764;
input n_1503;
input n_2238;
input n_2529;
input n_2374;
input n_462;
input n_1196;
input n_1181;
input n_32;
input n_1999;
input n_410;
input n_2380;
input n_1187;
input n_1131;
input n_1225;
input n_737;
input n_137;
input n_1298;
input n_1745;
input n_1366;
input n_232;
input n_52;
input n_2084;
input n_568;
input n_2278;
input n_1088;
input n_77;
input n_1424;
input n_766;
input n_1835;
input n_1457;
input n_377;
input n_2482;
input n_1682;
input n_1836;
input n_520;
input n_870;
input n_2547;
input n_1453;
input n_279;
input n_945;
input n_958;
input n_2554;
input n_2248;
input n_813;
input n_419;
input n_1985;
input n_2288;
input n_146;
input n_270;
input n_338;
input n_995;
input n_285;
input n_1909;
input n_2156;
input n_1184;
input n_1961;
input n_202;
input n_1535;
input n_500;
input n_665;
input n_754;
input n_903;
input n_871;
input n_2323;
input n_1073;
input n_239;
input n_402;
input n_1979;
input n_1277;
input n_2107;
input n_1746;
input n_54;
input n_829;
input n_1761;
input n_1062;
input n_339;
input n_738;
input n_1690;
input n_2221;
input n_672;
input n_740;
input n_1283;
input n_167;
input n_2317;
input n_1974;
input n_1736;
input n_1018;
input n_2342;
input n_2200;
input n_69;
input n_259;
input n_2442;
input n_953;
input n_1364;
input n_2390;
input n_143;
input n_1888;
input n_1224;
input n_2109;
input n_1425;
input n_625;
input n_557;
input n_2322;
input n_1107;
input n_1688;
input n_989;
input n_242;
input n_645;
input n_1944;
input n_331;
input n_559;
input n_2233;
input n_2370;
input n_267;
input n_495;
input n_1988;
input n_350;
input n_381;
input n_795;
input n_721;
input n_1084;
input n_1718;
input n_1276;
input n_1936;
input n_2149;
input n_2277;
input n_200;
input n_1428;
input n_1284;
input n_1241;
input n_821;
input n_561;
input n_770;
input n_1514;
input n_2539;
input n_1528;
input n_507;
input n_486;
input n_901;
input n_569;
input n_2078;
input n_1145;
input n_971;
input n_2359;
input n_2201;
input n_787;
input n_1650;
input n_31;
input n_1519;
input n_1195;
input n_2049;
input n_1522;
input n_518;
input n_1207;
input n_222;
input n_786;
input n_1404;
input n_868;
input n_2232;
input n_1847;
input n_2458;
input n_1542;
input n_1314;
input n_1512;
input n_2227;
input n_2301;
input n_1539;
input n_884;
input n_1851;
input n_2162;
input n_1415;
input n_1034;
input n_1652;
input n_2192;
input n_1676;
input n_1085;
input n_277;
input n_1636;
input n_432;
input n_293;
input n_823;
input n_1900;
input n_620;
input n_93;
input n_1074;
input n_859;
input n_1765;
input n_108;
input n_1889;
input n_587;
input n_1977;
input n_693;
input n_863;
input n_303;
input n_1254;
input n_929;
input n_2433;
input n_206;
input n_352;
input n_899;
input n_1703;
input n_2332;
input n_2391;
input n_611;
input n_1295;
input n_2060;
input n_1850;
input n_238;
input n_365;
input n_2004;
input n_1013;
input n_1495;
input n_1637;
input n_136;
input n_334;
input n_2427;
input n_192;
input n_661;
input n_2098;
input n_1751;
input n_300;
input n_533;
input n_1917;
input n_2456;
input n_104;
input n_1924;
input n_438;
input n_1560;
input n_1654;
input n_2341;
input n_1548;
input n_16;
input n_1811;
input n_2045;
input n_440;
input n_273;
input n_1396;
input n_1230;
input n_612;
input n_333;
input n_1840;
input n_376;
input n_512;
input n_1597;
input n_1771;
input n_1544;
input n_579;
input n_844;
input n_1012;
input n_1267;
input n_2061;
input n_2094;
input n_2512;
input n_1354;
input n_1790;
input n_149;
input n_1213;
input n_2382;
input n_237;
input n_2043;
input n_780;
input n_2349;
input n_1918;
input n_1021;
input n_1443;
input n_491;
input n_1465;
input n_1949;
input n_1595;
input n_1142;
input n_1140;
input n_705;
input n_570;
input n_260;
input n_942;
input n_1437;
input n_7;
input n_2077;
input n_1378;
input n_461;
input n_1121;
input n_1416;
input n_209;
input n_490;
input n_1461;
input n_17;
input n_1391;
input n_1947;
input n_225;
input n_1599;
input n_1876;
input n_1006;
input n_1830;
input n_575;
input n_546;
input n_503;
input n_2527;
input n_1112;
input n_700;
input n_1159;
input n_772;
input n_1216;
input n_1245;
input n_1669;
input n_1675;
input n_2466;
input n_676;
input n_42;
input n_2038;
input n_2263;
input n_2116;
input n_2271;
input n_2145;
input n_2326;
input n_1838;
input n_1594;
input n_680;
input n_1935;
input n_287;
input n_1716;
input n_302;
input n_1872;
input n_380;
input n_1585;
input n_2281;
input n_1432;
input n_94;
input n_2245;
input n_4;
input n_249;
input n_1108;
input n_355;
input n_212;
input n_65;
input n_123;
input n_444;
input n_851;
input n_1590;
input n_1351;
input n_2216;
input n_1274;
input n_257;
input n_2426;
input n_652;
input n_1819;
input n_475;
input n_135;
input n_947;
input n_2134;
input n_930;
input n_1260;
input n_1179;
input n_468;
input n_102;
input n_182;
input n_696;
input n_1442;
input n_482;
input n_798;
input n_577;
input n_1833;
input n_407;
input n_1691;
input n_27;
input n_916;
input n_1386;
input n_912;
input n_1884;
input n_460;
input n_1555;
input n_1842;
input n_2499;
input n_2549;
input n_366;
input n_762;
input n_1253;
input n_1468;
input n_1661;
input n_555;
input n_804;
input n_1656;
input n_1382;
input n_966;
input n_992;
input n_955;
input n_1182;
input n_794;
input n_78;
input n_2166;
input n_1692;
input n_1562;
input n_514;
input n_418;
input n_2185;
input n_2398;
input n_1376;
input n_513;
input n_288;
input n_179;
input n_1292;
input n_1178;
input n_1972;
input n_2015;
input n_1435;
input n_1750;
input n_1026;
input n_1506;
input n_1610;
input n_2202;
input n_2072;
input n_306;
input n_2415;
input n_92;
input n_203;
input n_436;
input n_150;
input n_324;
input n_2087;
input n_669;
input n_931;
input n_1491;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_967;
input n_1083;
input n_2161;
input n_1418;
input n_746;
input n_1357;
input n_292;
input n_1079;
input n_1787;
input n_2462;
input n_1389;
input n_2155;
input n_615;
input n_1139;
input n_76;
input n_2439;
input n_517;
input n_1312;
input n_1717;
input n_0;
input n_1812;
input n_824;
input n_428;
input n_159;
input n_2172;
input n_892;
input n_1880;
input n_959;
input n_30;
input n_2365;
input n_2257;
input n_1399;
input n_1101;
input n_1567;
input n_1343;
input n_563;
input n_2219;
input n_1855;
input n_2100;
input n_2333;
input n_144;
input n_990;
input n_1623;
input n_1903;
input n_867;
input n_2147;
input n_2435;
input n_1226;
input n_2224;
input n_944;
input n_749;
input n_1932;
input n_1780;
input n_1970;
input n_1920;
input n_2083;
input n_815;
input n_542;
input n_2167;
input n_2293;
input n_1340;
input n_470;
input n_1240;
input n_1087;
input n_2400;
input n_632;
input n_477;
input n_650;
input n_2388;
input n_425;
input n_2273;
input n_1433;
input n_1911;
input n_1825;
input n_1908;
input n_1155;
input n_1071;
input n_712;
input n_976;
input n_909;
input n_1392;
input n_767;
input n_1832;
input n_1841;
input n_1680;
input n_2066;
input n_2302;
input n_964;
input n_1627;
input n_2220;
input n_382;
input n_489;
input n_2294;
input n_80;
input n_2274;
input n_251;
input n_974;
input n_506;
input n_1731;
input n_799;
input n_1147;
input n_2378;
input n_397;
input n_2467;
input n_471;
input n_351;
input n_965;
input n_1914;
input n_155;
input n_2253;
input n_934;
input n_2213;
input n_1447;
input n_2363;
input n_1220;
input n_356;
input n_2019;
input n_698;
input n_2130;
input n_1674;
input n_2021;
input n_2025;
input n_2160;
input n_1992;
input n_124;
input n_307;
input n_1209;
input n_1020;
input n_1563;
input n_646;
input n_2507;
input n_2142;
input n_1633;
input n_34;
input n_404;
input n_172;
input n_1913;
input n_2069;
input n_2495;
input n_1058;
input n_2328;
input n_347;
input n_2434;
input n_1042;
input n_183;
input n_1234;
input n_2311;
input n_479;
input n_1578;
input n_2261;
input n_1455;
input n_2287;
input n_299;
input n_836;
input n_2223;
input n_1279;
input n_2473;
input n_2144;
input n_2511;
input n_564;
input n_133;
input n_66;
input n_205;
input n_1029;
input n_1247;
input n_760;
input n_522;
input n_2438;
input n_1568;
input n_20;
input n_1483;
input n_1363;
input n_367;
input n_1111;
input n_970;
input n_1689;
input n_2535;
input n_713;
input n_1255;
input n_1646;
input n_598;
input n_345;
input n_2262;
input n_1237;
input n_927;
input n_261;
input n_1095;
input n_1728;
input n_2335;
input n_370;
input n_706;
input n_2120;
input n_286;
input n_1401;
input n_1419;
input n_1531;
input n_776;
input n_424;
input n_2041;
input n_2113;
input n_1933;
input n_1651;
input n_85;
input n_130;
input n_1387;
input n_466;
input n_1263;
input n_346;
input n_1817;
input n_2404;
input n_2168;
input n_348;
input n_552;
input n_2312;
input n_670;
input n_1826;
input n_379;
input n_138;
input n_162;
input n_264;
input n_2483;
input n_441;
input n_1951;
input n_2490;
input n_1032;
input n_1217;
input n_1496;
input n_637;
input n_1592;
input n_73;
input n_327;
input n_1259;
input n_1177;
input n_1231;
input n_2132;
input n_980;
input n_1618;
input n_1869;
input n_1743;
input n_905;
input n_207;
input n_720;
input n_926;
input n_41;
input n_1943;
input n_2296;
input n_194;
input n_1802;
input n_2178;
input n_2112;
input n_1163;
input n_186;
input n_1795;
input n_1384;
input n_2237;
input n_145;
input n_2146;
input n_1868;
input n_59;
input n_1501;
input n_2241;
input n_2373;
input n_1173;
input n_2350;
input n_1068;
input n_1198;
input n_2531;
input n_1570;
input n_2099;
input n_487;
input n_1518;
input n_1456;
input n_90;
input n_1879;
input n_1886;
input n_1648;
input n_2187;
input n_1413;
input n_2481;
input n_2129;
input n_855;
input n_2327;
input n_158;
input n_808;
input n_1365;
input n_2476;
input n_553;
input n_2059;
input n_2437;
input n_1439;
input n_814;
input n_578;
input n_2074;
input n_1665;
input n_1287;
input n_405;
input n_1611;
input n_2122;
input n_120;
input n_2399;
input n_320;
input n_1414;
input n_1134;
input n_2067;
input n_1484;
input n_1901;
input n_647;
input n_2055;
input n_2027;
input n_1423;
input n_2117;
input n_481;
input n_600;
input n_1053;
input n_1609;
input n_1939;
input n_2308;
input n_2242;
input n_1906;
input n_529;
input n_1899;
input n_2195;
input n_502;
input n_2194;
input n_218;
input n_1467;
input n_247;
input n_1828;
input n_2159;
input n_1798;
input n_1304;
input n_1608;
input n_1744;
input n_2267;
input n_1105;
input n_547;
input n_439;
input n_604;
input n_677;
input n_478;
input n_703;
input n_1349;
input n_1709;
input n_1061;
input n_2102;
input n_326;
input n_681;
input n_227;
input n_874;
input n_2286;
input n_2023;
input n_1278;
input n_707;
input n_11;
input n_129;
input n_126;
input n_983;
input n_590;
input n_699;
input n_727;
input n_301;
input n_1726;
input n_2075;
input n_2523;
input n_1945;
input n_545;
input n_1015;
input n_2418;
input n_1377;
input n_1162;
input n_536;
input n_1614;
input n_2031;
input n_2496;
input n_2118;
input n_325;
input n_1740;
input n_1602;
input n_688;
input n_636;
input n_427;
input n_1098;
input n_1490;
input n_2338;
input n_442;
input n_777;
input n_1553;
input n_1080;
input n_920;
input n_1760;
input n_1086;
input n_1092;
input n_2225;
input n_986;
input n_1104;
input n_1963;
input n_729;
input n_887;
input n_2057;
input n_2218;
input n_1122;
input n_1205;
input n_1408;
input n_163;
input n_1693;
input n_2125;
input n_1132;
input n_390;
input n_1156;
input n_501;
input n_2184;
input n_314;
input n_1823;
input n_1120;
input n_1202;
input n_627;
input n_2254;
input n_1188;
input n_1498;
input n_1371;
input n_2033;
input n_233;
input n_957;
input n_388;
input n_1402;
input n_1242;
input n_1607;
input n_1489;
input n_1218;
input n_2217;
input n_221;
input n_321;
input n_86;
input n_2226;
input n_1586;
input n_861;
input n_1543;
input n_1431;
input n_877;
input n_1119;
input n_1863;
input n_1763;
input n_1666;
input n_1500;
input n_616;
input n_2214;
input n_1055;
input n_1395;
input n_1346;
input n_2256;
input n_1189;
input n_1089;
input n_281;
input n_1859;
input n_262;
input n_1502;
input n_1523;
input n_2190;
input n_1478;
input n_1883;
input n_2516;
input n_1969;
input n_735;
input n_297;
input n_1005;
input n_527;
input n_2379;
input n_46;
input n_84;
input n_1294;
input n_1667;
input n_845;
input n_888;
input n_2300;
input n_1649;
input n_2452;
input n_1677;
input n_2470;
input n_1927;
input n_1297;
input n_178;
input n_551;
input n_417;
input n_1708;
input n_70;
input n_343;
input n_1222;
input n_2284;
input n_1844;
input n_2283;
input n_582;
input n_2526;
input n_1957;
input n_1953;
input n_755;
input n_1097;
input n_1219;
input n_1711;
input n_710;
input n_1919;
input n_534;
input n_1791;
input n_2508;
input n_2124;
input n_1894;
input n_1460;
input n_1239;
input n_278;
input n_2266;
input n_2449;
input n_560;
input n_890;
input n_842;
input n_148;
input n_1898;
input n_451;
input n_745;
input n_1741;
input n_1572;
input n_1907;
input n_1793;
input n_61;
input n_742;
input n_1081;
input n_1373;
input n_1975;
input n_1388;
input n_1266;
input n_1540;
input n_1719;
input n_2119;
input n_769;
input n_1797;
input n_2366;
input n_2493;
input n_13;
input n_1753;
input n_1990;
input n_1372;
input n_476;
input n_832;
input n_55;
input n_535;
input n_744;
input n_1895;
input n_2474;
input n_982;
input n_1800;
input n_915;
input n_215;
input n_1075;
input n_2008;
input n_454;
input n_298;
input n_1331;
input n_1890;
input n_1529;
input n_1227;
input n_2127;
input n_655;
input n_1734;
input n_1860;
input n_403;
input n_2460;
input n_1007;
input n_1580;
input n_1319;
input n_657;
input n_837;
input n_812;
input n_2448;
input n_2211;
input n_2292;
input n_2480;
input n_606;
input n_951;
input n_862;
input n_1700;
input n_659;
input n_1332;
input n_2306;
input n_509;
input n_1854;
input n_666;
input n_1747;
input n_2071;
input n_2424;
input n_430;
input n_1206;
input n_1729;
input n_722;
input n_1508;
input n_2414;
input n_2082;
input n_1532;
input n_1171;
input n_1030;
input n_785;
input n_2389;
input n_1309;
input n_999;
input n_2280;
input n_1766;
input n_1338;
input n_1342;
input n_456;
input n_1867;
input n_852;
input n_1394;
input n_704;
input n_1060;
input n_1044;
input n_1714;
input n_521;
input n_2140;
input n_873;
input n_1301;
input n_1748;
input n_2157;
input n_1966;
input n_1243;
input n_2171;
input n_2468;
input n_1400;
input n_342;
input n_2035;
input n_1466;
input n_1513;
input n_1527;
input n_358;
input n_1783;
input n_608;
input n_2494;
input n_1538;
input n_2457;
input n_2128;
input n_1037;
input n_1329;
input n_317;
input n_1993;
input n_1545;
input n_134;
input n_1257;
input n_1480;
input n_1954;
input n_1668;
input n_1878;
input n_2540;
input n_1605;
input n_1078;
input n_266;
input n_2486;
input n_1897;
input n_157;
input n_2520;
input n_2137;
input n_1161;
input n_2489;
input n_811;
input n_624;
input n_791;
input n_876;
input n_618;
input n_1191;
input n_2492;
input n_736;
input n_1025;
input n_1215;
input n_241;
input n_1449;
input n_2337;
input n_2265;
input n_687;
input n_797;
input n_2026;
input n_1786;
input n_480;
input n_1327;
input n_1475;
input n_211;
input n_642;
input n_1804;
input n_2106;
input n_97;
input n_408;
input n_1406;
input n_595;
input n_1405;
input n_602;
input n_2272;
input n_1757;
input n_592;
input n_1499;
input n_854;
input n_1318;
input n_2091;
input n_393;
input n_1632;
input n_1769;
input n_474;
input n_1929;
input n_1950;
input n_2264;
input n_805;
input n_2032;
input n_2090;
input n_295;
input n_1658;
input n_190;
input n_2249;
input n_1072;
input n_695;
input n_1526;
input n_1305;
input n_64;
input n_180;
input n_730;
input n_386;
input n_1596;
input n_2348;
input n_1281;
input n_516;
input n_2364;
input n_1997;
input n_1137;
input n_1873;
input n_1258;
input n_197;
input n_640;
input n_463;
input n_1476;
input n_1524;
input n_1733;
input n_1856;
input n_2016;
input n_943;
input n_1118;
input n_678;
input n_651;
input n_1874;
input n_1293;
input n_961;
input n_469;
input n_1046;
input n_1807;
input n_726;
input n_1123;
input n_1657;
input n_878;
input n_1784;
input n_771;
input n_1321;
input n_752;
input n_2307;
input n_71;
input n_1488;
input n_985;
input n_421;
input n_1330;
input n_906;
input n_1180;
input n_1697;
input n_2295;
input n_283;
input n_806;
input n_1984;
input n_1350;
input n_1556;
input n_649;
input n_1561;
input n_2412;
input n_374;
input n_1352;
input n_2405;
input n_1824;
input n_643;
input n_1492;
input n_226;
input n_2383;
input n_1441;
input n_1822;
input n_682;
input n_36;
input n_1616;
input n_2416;
input n_819;
input n_2386;
input n_1971;
input n_586;
input n_1324;
input n_1429;
input n_2064;
input n_2353;
input n_2528;
input n_1778;
input n_1776;
input n_686;
input n_605;
input n_1154;
input n_584;
input n_1557;
input n_1759;
input n_1829;
input n_2325;
input n_1130;
input n_1450;
input n_349;
input n_756;
input n_2022;
input n_1016;
input n_2298;
input n_1149;
input n_1505;
input n_2408;
input n_2320;
input n_979;
input n_2329;
input n_1642;
input n_2417;
input n_2;
input n_2525;
input n_1815;
input n_897;
input n_2546;
input n_949;
input n_2454;
input n_1493;
input n_515;
input n_807;
input n_891;
input n_885;
input n_1659;
input n_2354;
input n_198;
input n_1864;
input n_1887;
input n_1208;
input n_1987;
input n_396;
input n_2368;
input n_802;
input n_23;
input n_1151;
input n_554;
input n_960;
input n_2352;
input n_2502;
input n_1256;
input n_87;
input n_714;
input n_2170;
input n_790;
input n_2244;
input n_2143;
input n_2393;
input n_354;
input n_140;
input n_725;
input n_2377;
input n_1577;
input n_151;
input n_1448;
input n_2198;
input n_28;
input n_1009;
input n_230;
input n_1133;
input n_154;
input n_883;
input n_142;
input n_473;
input n_1852;
input n_801;
input n_1286;
input n_818;
input n_1685;
input n_779;
input n_2410;
input n_2314;
input n_2477;
input n_2279;
input n_594;
input n_2222;
input n_1995;
input n_1877;
input n_1397;
input n_35;
input n_1052;
input n_272;
input n_1333;
input n_1306;
input n_1849;
input n_2076;
input n_2133;
input n_2203;
input n_833;
input n_1426;
input n_2250;
input n_2497;
input n_2247;
input n_2230;
input n_879;
input n_1117;
input n_38;
input n_422;
input n_1269;
input n_1303;
input n_1547;
input n_1438;
input n_1541;
input n_597;
input n_75;
input n_2001;
input n_1047;
input n_95;
input n_2506;
input n_1472;
input n_2413;
input n_1593;
input n_1050;
input n_566;
input n_2158;
input n_2285;
input n_152;
input n_169;
input n_106;
input n_1201;
input n_1288;
input n_173;
input n_858;
input n_1185;
input n_2475;
input n_2173;
input n_335;
input n_1035;
input n_1143;
input n_344;
input n_2070;
input n_2136;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_1090;
input n_2403;
input n_1367;
input n_2044;
input n_166;
input n_253;
input n_928;
input n_1153;
input n_271;
input n_465;
input n_825;
input n_1103;
input n_732;
input n_1565;
input n_1192;
input n_128;
input n_224;
input n_82;
input n_894;
input n_1380;
input n_1624;
input n_1801;
input n_420;
input n_1291;
input n_562;
input n_2020;
input n_748;
input n_2310;
input n_510;
input n_1045;
input n_256;
input n_1160;
input n_1882;
input n_1976;
input n_1023;
input n_1881;
input n_988;
input n_330;
input n_914;
input n_400;
input n_689;
input n_1116;
input n_282;
input n_328;
input n_368;
input n_1958;
input n_467;
input n_1511;
input n_2177;
input n_1422;
input n_1965;
input n_644;
input n_1197;
input n_276;
input n_497;
input n_1165;
input n_1641;
input n_168;
input n_81;
input n_538;
input n_1517;
input n_2036;
input n_576;
input n_843;
input n_511;
input n_455;
input n_429;
input n_588;
input n_638;
input n_2003;
input n_2533;
input n_2210;
input n_1307;
input n_1128;
input n_2053;
input n_1671;
input n_1417;
input n_1048;
input n_2343;
input n_775;
input n_667;
input n_2419;
input n_1049;
input n_2330;
input n_14;
input n_869;
input n_141;
input n_846;
input n_1398;
input n_1921;
input n_2450;
input n_2411;
input n_1356;
input n_1341;
input n_2234;
input n_2309;
input n_1504;
input n_1955;
input n_2110;
input n_2431;
input n_1773;
input n_1440;
input n_1370;
input n_1603;
input n_305;
input n_312;
input n_56;
input n_60;
input n_728;
input n_413;
input n_2401;
input n_715;
input n_889;
input n_1066;
input n_1549;
input n_2331;
input n_935;
input n_2478;
input n_685;
input n_911;
input n_361;
input n_89;
input n_623;
input n_1712;
input n_1403;
input n_1065;
input n_453;
input n_1534;
input n_1948;
input n_74;
input n_810;
input n_19;
input n_40;
input n_1290;
input n_181;
input n_1959;
input n_617;
input n_2396;
input n_543;
input n_1362;
input n_1559;
input n_2121;
input n_236;
input n_601;
input n_683;
input n_565;
input n_628;
input n_1300;
input n_1960;
input n_2068;
input n_743;
input n_1194;
input n_1647;
input n_1546;
input n_1420;
input n_2553;
input n_907;
input n_1454;
input n_660;
input n_464;
input n_2459;
input n_962;
input n_941;
input n_1210;
input n_847;
input n_747;
input n_1622;
input n_1135;
input n_918;
input n_1968;
input n_107;
input n_1885;
input n_639;
input n_452;
input n_673;
input n_2196;
input n_1038;
input n_2371;
input n_1978;
input n_414;
input n_571;
input n_1521;
input n_1694;
input n_1940;
input n_6;
input n_284;
input n_593;
input n_1695;
input n_1164;
input n_37;
input n_58;
input n_2313;
input n_609;
input n_1193;
input n_1345;
input n_613;
input n_1022;
input n_1336;
input n_1033;
input n_1774;
input n_409;
input n_171;
input n_519;
input n_384;
input n_1166;
input n_1056;
input n_2007;
input n_526;
input n_1994;
input n_1767;
input n_1040;
input n_674;
input n_1158;
input n_316;
input n_125;
input n_1973;
input n_1444;
input n_1803;
input n_820;
input n_1749;
input n_43;
input n_872;
input n_1653;
input n_254;
input n_2303;
input n_1157;
input n_1584;
input n_234;
input n_848;
input n_1664;
input n_280;
input n_629;
input n_1739;
input n_161;
input n_1814;
input n_532;
input n_2154;
input n_2441;
input n_2236;
input n_1789;
input n_763;
input n_1986;
input n_2174;
input n_99;
input n_540;
input n_216;
input n_692;
input n_5;
input n_2054;
input n_1857;
input n_2315;
input n_984;
input n_1687;
input n_2073;
input n_223;
input n_2150;
input n_1552;
input n_750;
input n_834;
input n_1612;
input n_2498;
input n_800;
input n_2046;
input n_1816;
input n_1910;
input n_1756;
input n_1606;
input n_2189;
input n_395;
input n_621;
input n_1587;
input n_213;
input n_2093;
input n_2340;
input n_2018;
input n_1772;
input n_67;
input n_2444;
input n_1014;
input n_724;
input n_2204;
input n_1427;
input n_1481;
input n_2040;
input n_493;
input n_1311;
input n_2199;
input n_1956;
input n_1589;
input n_114;
input n_2151;
input n_1100;
input n_585;
input n_875;
input n_1617;
input n_2455;
input n_827;
input n_2231;
input n_697;
input n_622;
input n_1626;
input n_1962;
input n_1335;
input n_1715;
input n_296;
input n_2305;
input n_880;
input n_793;
input n_2114;
input n_1175;
input n_2289;
input n_132;
input n_2530;
input n_2299;
input n_751;
input n_1027;
input n_1070;
input n_2406;
input n_1621;
input n_739;
input n_1485;
input n_1028;
input n_1221;
input n_530;
input n_1785;
input n_792;
input n_1262;
input n_1942;
input n_2180;
input n_580;
input n_1579;
input n_494;
input n_2181;
input n_434;
input n_2014;
input n_975;
input n_229;
input n_394;
input n_923;
input n_1645;
input n_1124;
input n_1381;
input n_1494;
input n_932;
input n_1893;
input n_1183;
input n_1326;
input n_2276;
input n_1805;
input n_2282;
input n_981;
input n_2141;
input n_1110;
input n_1758;
input n_2503;
input n_2270;
input n_243;
input n_2443;
input n_1407;
input n_185;
input n_2465;
input n_1204;
input n_1554;
input n_994;
input n_2428;
input n_1360;
input n_973;
input n_268;
input n_972;
input n_2251;
input n_164;
input n_184;
input n_856;
input n_1248;
input n_1176;
input n_1564;
input n_2010;
input n_1054;
input n_508;
input n_118;
input n_121;
input n_1679;
input n_2126;
input n_1952;
input n_2425;
input n_2394;
input n_1858;
input n_353;
input n_1678;
input n_1482;
input n_1361;
input n_2356;
input n_1601;
input n_1057;
input n_191;
input n_2487;
input n_1834;
input n_978;
input n_1011;
input n_1520;
input n_2534;
input n_2488;
input n_1509;
input n_828;
input n_322;
input n_1411;
input n_1359;
input n_558;
input n_1721;
input n_116;
input n_39;
input n_653;
input n_1445;
input n_1317;
input n_2050;
input n_2197;
input n_783;
input n_2550;
input n_556;
input n_1127;
input n_170;
input n_1536;
input n_1471;
input n_2385;
input n_160;
input n_119;
input n_2387;
input n_1008;
input n_332;
input n_581;
input n_294;
input n_1024;
input n_830;
input n_176;
input n_2291;
input n_1980;
input n_2518;
input n_987;
input n_936;
input n_2510;
input n_1620;
input n_2501;
input n_2542;
input n_1385;
input n_1525;
input n_1998;
input n_2165;
input n_541;
input n_499;
input n_1775;
input n_788;
input n_12;
input n_908;
input n_1036;
input n_2169;
input n_341;
input n_1270;
input n_109;
input n_1167;
input n_1272;
input n_549;
input n_591;
input n_969;
input n_2028;
input n_919;
input n_1663;
input n_50;
input n_2092;
input n_2175;
input n_1625;
input n_2086;
input n_1926;
input n_2402;
input n_318;
input n_1458;
input n_103;
input n_244;
input n_679;
input n_1630;
input n_220;
input n_663;
input n_1720;
input n_2409;
input n_443;
input n_2176;
input n_1412;
input n_1738;
input n_1550;
input n_528;
input n_1358;
input n_1200;
input n_387;
input n_406;
input n_826;
input n_139;
input n_2453;
input n_2344;
input n_1922;
input n_1735;
input n_1788;
input n_391;
input n_940;
input n_2392;
input n_1537;
input n_2138;
input n_2065;
input n_2543;
input n_2321;
input n_1077;
input n_607;
input n_956;
input n_445;
input n_1930;
input n_765;
input n_1809;
input n_1843;
input n_1904;
input n_122;
input n_2000;
input n_1268;
input n_385;
input n_2395;
input n_917;
input n_1271;
input n_372;
input n_2096;
input n_2440;
input n_2186;
input n_15;
input n_1530;
input n_2215;
input n_631;
input n_399;
input n_1170;
input n_2258;
input n_1261;
input n_2471;
input n_702;
input n_857;
input n_898;
input n_363;
input n_968;
input n_1067;
input n_1235;
input n_1323;
input n_2375;
input n_1462;
input n_1937;
input n_2012;
input n_1064;
input n_633;
input n_900;
input n_1446;
input n_1282;
input n_1701;
input n_1093;
input n_1551;
input n_2039;
input n_1755;
input n_1285;
input n_193;
input n_733;
input n_761;
input n_2212;
input n_731;
input n_336;
input n_1813;
input n_315;
input n_2268;
input n_311;
input n_1452;
input n_1573;
input n_8;
input n_668;
input n_758;
input n_2252;
input n_2111;
input n_2420;
input n_1996;
input n_1106;
input n_2009;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_816;
input n_1322;
input n_1473;
input n_835;
input n_446;
input n_1076;
input n_2024;
input n_1348;
input n_753;
input n_2445;
input n_1770;
input n_701;
input n_1003;
input n_2469;
input n_1125;
input n_2103;
input n_2358;
input n_1710;
input n_1865;
input n_2522;
input n_2463;
input n_309;
input n_1344;
input n_115;
input n_2355;
input n_1390;
input n_401;
input n_485;
input n_1792;
input n_504;
input n_2062;
input n_483;
input n_435;
input n_1141;
input n_1629;
input n_291;
input n_1640;
input n_822;
input n_1094;
input n_840;
input n_1459;
input n_2153;
input n_2324;
input n_1510;
input n_2505;
input n_2139;
input n_1099;
input n_839;
input n_79;
input n_1754;
input n_3;
input n_759;
input n_567;
input n_2397;
input n_91;
input n_2521;
input n_240;
input n_369;
input n_1727;
input n_2235;
input n_44;
input n_1991;
input n_1575;
input n_1848;
input n_1892;
input n_1172;
input n_614;
input n_1212;
input n_831;
input n_778;
input n_48;
input n_1619;
input n_2351;
input n_188;
input n_2260;
input n_323;
input n_550;
input n_1315;
input n_1660;
input n_1902;
input n_997;
input n_635;
input n_2206;
input n_2541;
input n_694;
input n_1643;
input n_1320;
input n_1113;
input n_2347;
input n_248;
input n_1152;
input n_2447;
input n_2034;
input n_1845;
input n_2538;
input n_1934;
input n_2101;
input n_921;
input n_2362;
input n_1615;
input n_1236;
input n_228;
input n_2104;
input n_1265;
input n_1576;
input n_2105;
input n_1470;
input n_671;
input n_1533;
input n_1806;
input n_2372;
input n_2552;
input n_1;
input n_1409;
input n_1148;
input n_1588;
input n_1684;
input n_1673;
input n_2422;
input n_1334;
input n_654;
input n_2290;
input n_2088;
input n_1275;
input n_488;
input n_904;
input n_505;
input n_88;
input n_2005;
input n_2048;
input n_1696;
input n_498;
input n_1875;
input n_1059;
input n_684;
input n_2429;
input n_2108;
input n_1039;
input n_2246;
input n_539;
input n_1150;
input n_977;
input n_449;
input n_2339;
input n_392;
input n_1628;
input n_1289;
input n_1831;
input n_2532;
input n_2191;
input n_1497;
input n_1866;
input n_2472;
input n_2056;
input n_459;
input n_1136;
input n_2515;
input n_1782;
input n_458;
input n_1190;
input n_1600;
input n_1144;
input n_383;
input n_838;
input n_1558;
input n_1941;
input n_1316;
input n_175;
input n_2519;
input n_950;
input n_1017;
input n_711;
input n_734;
input n_1915;
input n_2360;
input n_723;
input n_1393;
input n_2240;
input n_658;
input n_630;
input n_1369;
input n_53;
input n_362;
input n_310;
input n_1781;
input n_709;
input n_2544;
input n_24;
input n_809;
input n_2085;
input n_2432;
input n_1686;
input n_1964;
input n_235;
input n_881;
input n_1019;
input n_1477;
input n_1777;
input n_2188;
input n_1982;
input n_2097;
input n_662;
input n_641;
input n_2430;
input n_2504;
input n_910;
input n_290;
input n_741;
input n_939;
input n_1410;
input n_2297;
input n_371;
input n_199;
input n_217;
input n_1114;
input n_1325;
input n_1742;
input n_708;
input n_308;
input n_1223;
input n_2545;
input n_201;
input n_1768;
input n_2513;
input n_2193;
input n_2369;
input n_572;
input n_1199;
input n_865;
input n_10;
input n_1273;
input n_1983;
input n_1041;
input n_2451;
input n_2115;
input n_993;
input n_1862;
input n_948;
input n_2017;
input n_922;
input n_1004;
input n_1810;
input n_448;
input n_1347;
input n_860;
input n_1043;
input n_255;
input n_450;
input n_1923;
input n_1764;
input n_896;
input n_1737;
input n_1479;
input n_1613;
input n_902;
input n_1031;
input n_1723;
input n_1638;
input n_853;
input n_716;
input n_1571;
input n_1698;
input n_196;
input n_1337;
input n_774;
input n_1946;
input n_2148;
input n_933;
input n_1779;
input n_596;
input n_954;
input n_2051;
input n_1168;
input n_1821;
input n_219;
input n_1310;
input n_231;
input n_656;
input n_492;
input n_574;
input n_252;
input n_664;
input n_1591;
input n_1229;
input n_1683;
input n_2548;
input n_68;
input n_1896;
input n_2164;
input n_1732;
input n_415;
input n_2381;
input n_1967;
input n_2384;
input n_2179;
input n_63;
input n_1280;
input n_544;
input n_1516;
input n_1186;
input n_1705;
input n_599;
input n_768;
input n_1091;
input n_2052;
input n_2485;
input n_537;
input n_1063;
input n_25;
input n_991;
input n_2183;
input n_2205;
input n_83;
input n_2275;
input n_389;
input n_1724;
input n_1670;
input n_1707;
input n_1799;
input n_2080;
input n_2058;
input n_1126;
input n_2357;
input n_2029;
input n_195;
input n_1846;
input n_1912;
input n_938;
input n_1891;
input n_1328;
input n_895;
input n_110;
input n_304;
input n_1639;
input n_583;
input n_2209;
input n_2421;
input n_1302;
input n_1000;
input n_313;
input n_626;
input n_378;
input n_1581;
input n_1928;
input n_98;
input n_946;
input n_757;
input n_2047;
input n_375;
input n_113;
input n_1655;
input n_1818;
input n_33;
input n_1146;
input n_1634;
input n_1203;
input n_998;
input n_1699;
input n_1598;
input n_2269;
input n_472;
input n_937;
input n_1474;
input n_2081;
input n_2536;
input n_2524;
input n_265;
input n_1583;
input n_1604;
input n_208;
input n_1631;
input n_1702;
input n_156;
input n_174;
input n_275;
input n_100;
input n_1794;
input n_1375;
input n_147;
input n_204;
input n_1232;
input n_996;
input n_1211;
input n_1368;
input n_963;
input n_1264;
input n_51;
input n_1082;
input n_1725;
input n_496;
input n_2318;
input n_1827;
input n_866;
input n_26;
input n_246;
input n_925;
input n_1752;
input n_1313;
input n_1001;
input n_1722;
input n_2361;
input n_1115;
input n_2229;
input n_1339;
input n_1002;
input n_1644;
input n_105;
input n_1051;
input n_2551;
input n_719;
input n_131;
input n_263;
input n_1102;
input n_360;
input n_2255;
input n_1129;
input n_1252;
input n_2239;
input n_250;
input n_1464;
input n_1296;
input n_773;
input n_2316;
input n_165;
input n_2464;
input n_1010;
input n_882;
input n_2304;
input n_1249;
input n_101;
input n_803;
input n_1871;
input n_2514;
input n_329;
input n_718;
input n_1434;
input n_340;
input n_1905;
input n_1569;
input n_289;
input n_9;
input n_112;
input n_45;
input n_548;
input n_2336;
input n_523;
input n_1662;
input n_457;
input n_1299;
input n_1870;
input n_177;
input n_2063;
input n_1925;
input n_782;
input n_364;
input n_258;
input n_431;
input n_2491;
input n_1861;
input n_2079;
input n_1228;
input n_2319;
input n_2152;
input n_2517;
input n_1931;
input n_1244;
input n_1796;
input n_411;
input n_484;
input n_2259;
input n_849;
input n_2095;
input n_22;
input n_1820;
input n_29;
input n_357;
input n_412;
input n_1251;
input n_1989;
input n_447;
input n_1421;
input n_2208;
input n_2423;
input n_1762;
input n_1233;
input n_1808;
input n_1574;
input n_1672;
input n_2228;
input n_1635;
input n_1704;
input n_893;
input n_1582;
input n_841;
input n_2479;
input n_886;
input n_1069;
input n_1981;
input n_2037;
input n_359;
input n_1308;
input n_573;
input n_796;
input n_127;
input n_531;
input n_2345;
input n_1730;
input n_1374;
input n_1451;
input n_2089;
input n_1487;
input n_675;

output n_14705;

wire n_3527;
wire n_2752;
wire n_4474;
wire n_9872;
wire n_9604;
wire n_10943;
wire n_10453;
wire n_12407;
wire n_7329;
wire n_4030;
wire n_12343;
wire n_13909;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_14469;
wire n_11913;
wire n_8165;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_12760;
wire n_11172;
wire n_12018;
wire n_14470;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_10678;
wire n_5402;
wire n_11190;
wire n_13957;
wire n_6581;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_11458;
wire n_11999;
wire n_3264;
wire n_5717;
wire n_10649;
wire n_13176;
wire n_10794;
wire n_12945;
wire n_2993;
wire n_4283;
wire n_9297;
wire n_11627;
wire n_2879;
wire n_4403;
wire n_10557;
wire n_13125;
wire n_8139;
wire n_11453;
wire n_4962;
wire n_14456;
wire n_7832;
wire n_8438;
wire n_12806;
wire n_12244;
wire n_11135;
wire n_11306;
wire n_2729;
wire n_4302;
wire n_14658;
wire n_12589;
wire n_5791;
wire n_7127;
wire n_13109;
wire n_4547;
wire n_14209;
wire n_13718;
wire n_5090;
wire n_3765;
wire n_8321;
wire n_5302;
wire n_10000;
wire n_12103;
wire n_7922;
wire n_7805;
wire n_9807;
wire n_2790;
wire n_7542;
wire n_12354;
wire n_11783;
wire n_7053;
wire n_11614;
wire n_9892;
wire n_5712;
wire n_11143;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_10704;
wire n_14334;
wire n_11431;
wire n_11799;
wire n_8699;
wire n_9263;
wire n_9734;
wire n_8037;
wire n_5479;
wire n_2646;
wire n_8257;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_11246;
wire n_10213;
wire n_11377;
wire n_13029;
wire n_3115;
wire n_9886;
wire n_5263;
wire n_4028;
wire n_10904;
wire n_5565;
wire n_9096;
wire n_6358;
wire n_8546;
wire n_6293;
wire n_8997;
wire n_13215;
wire n_14066;
wire n_9985;
wire n_9665;
wire n_14300;
wire n_12233;
wire n_11349;
wire n_7001;
wire n_10169;
wire n_10903;
wire n_13875;
wire n_11906;
wire n_6129;
wire n_13755;
wire n_14335;
wire n_14473;
wire n_13910;
wire n_4321;
wire n_10574;
wire n_13066;
wire n_5590;
wire n_10468;
wire n_2621;
wire n_14226;
wire n_6524;
wire n_9241;
wire n_9286;
wire n_4853;
wire n_8744;
wire n_9592;
wire n_5229;
wire n_12574;
wire n_6313;
wire n_12260;
wire n_7464;
wire n_8449;
wire n_9683;
wire n_10380;
wire n_10968;
wire n_4260;
wire n_13491;
wire n_7626;
wire n_9939;
wire n_3348;
wire n_12315;
wire n_10688;
wire n_3261;
wire n_9358;
wire n_9466;
wire n_8953;
wire n_11756;
wire n_7965;
wire n_13636;
wire n_7368;
wire n_9787;
wire n_8399;
wire n_2807;
wire n_6664;
wire n_8598;
wire n_10276;
wire n_7562;
wire n_11604;
wire n_9997;
wire n_7534;
wire n_13196;
wire n_7428;
wire n_12581;
wire n_4512;
wire n_6190;
wire n_8460;
wire n_12085;
wire n_4132;
wire n_13980;
wire n_7373;
wire n_8068;
wire n_6891;
wire n_4500;
wire n_9318;
wire n_10281;
wire n_13715;
wire n_12089;
wire n_8734;
wire n_12671;
wire n_14592;
wire n_8720;
wire n_2663;
wire n_10528;
wire n_8097;
wire n_5481;
wire n_6539;
wire n_12993;
wire n_13120;
wire n_8114;
wire n_4824;
wire n_8422;
wire n_12728;
wire n_7467;
wire n_14572;
wire n_8126;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_9714;
wire n_14405;
wire n_14598;
wire n_10399;
wire n_4741;
wire n_7526;
wire n_8664;
wire n_10131;
wire n_11721;
wire n_14378;
wire n_11736;
wire n_4143;
wire n_14430;
wire n_10634;
wire n_4273;
wire n_11444;
wire n_11891;
wire n_13058;
wire n_4136;
wire n_14094;
wire n_9809;
wire n_11492;
wire n_3144;
wire n_14636;
wire n_9613;
wire n_9354;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_12647;
wire n_9897;
wire n_9295;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_10595;
wire n_11767;
wire n_13180;
wire n_6253;
wire n_9119;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_9058;
wire n_6197;
wire n_7200;
wire n_8326;
wire n_11807;
wire n_3639;
wire n_3254;
wire n_11944;
wire n_13090;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_11474;
wire n_11819;
wire n_8504;
wire n_3015;
wire n_5744;
wire n_8920;
wire n_3870;
wire n_12080;
wire n_6808;
wire n_3749;
wire n_5691;
wire n_7937;
wire n_8985;
wire n_3482;
wire n_7490;
wire n_13069;
wire n_6295;
wire n_11409;
wire n_5403;
wire n_11692;
wire n_13138;
wire n_12599;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_6992;
wire n_3960;
wire n_10644;
wire n_12863;
wire n_3975;
wire n_8035;
wire n_11856;
wire n_5830;
wire n_9516;
wire n_13996;
wire n_13064;
wire n_4018;
wire n_8660;
wire n_3325;
wire n_6681;
wire n_4227;
wire n_5158;
wire n_9917;
wire n_12185;
wire n_5152;
wire n_8939;
wire n_11737;
wire n_11652;
wire n_11038;
wire n_5092;
wire n_13991;
wire n_6542;
wire n_13466;
wire n_9202;
wire n_13689;
wire n_13896;
wire n_11925;
wire n_14115;
wire n_6161;
wire n_3612;
wire n_4505;
wire n_11974;
wire n_12457;
wire n_6452;
wire n_10426;
wire n_5247;
wire n_9512;
wire n_9923;
wire n_8469;
wire n_8715;
wire n_5464;
wire n_7306;
wire n_10070;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_12792;
wire n_7507;
wire n_13458;
wire n_8176;
wire n_9677;
wire n_2956;
wire n_5210;
wire n_7441;
wire n_7215;
wire n_7379;
wire n_5292;
wire n_8327;
wire n_12556;
wire n_8991;
wire n_7438;
wire n_11200;
wire n_8855;
wire n_4119;
wire n_4443;
wire n_9811;
wire n_4000;
wire n_13762;
wire n_9508;
wire n_13441;
wire n_13532;
wire n_2686;
wire n_5086;
wire n_6136;
wire n_14236;
wire n_3458;
wire n_11597;
wire n_5843;
wire n_7874;
wire n_11309;
wire n_14156;
wire n_8539;
wire n_13118;
wire n_8630;
wire n_9308;
wire n_14587;
wire n_8533;
wire n_13830;
wire n_11233;
wire n_7108;
wire n_3511;
wire n_9638;
wire n_11047;
wire n_11068;
wire n_3012;
wire n_13912;
wire n_13768;
wire n_4529;
wire n_3850;
wire n_11476;
wire n_8435;
wire n_7695;
wire n_10245;
wire n_6156;
wire n_11611;
wire n_13111;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_8204;
wire n_11957;
wire n_5060;
wire n_13290;
wire n_12509;
wire n_12663;
wire n_9199;
wire n_12155;
wire n_13379;
wire n_7162;
wire n_4432;
wire n_11210;
wire n_3518;
wire n_2800;
wire n_9808;
wire n_7331;
wire n_10457;
wire n_5913;
wire n_8958;
wire n_13838;
wire n_4530;
wire n_11333;
wire n_11682;
wire n_9821;
wire n_13692;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_10715;
wire n_11381;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_11922;
wire n_5249;
wire n_13126;
wire n_12068;
wire n_10579;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_10707;
wire n_3539;
wire n_5757;
wire n_9265;
wire n_6872;
wire n_12332;
wire n_12858;
wire n_6644;
wire n_11352;
wire n_9143;
wire n_5062;
wire n_3862;
wire n_12641;
wire n_4912;
wire n_12140;
wire n_9845;
wire n_4226;
wire n_10112;
wire n_14505;
wire n_10556;
wire n_14150;
wire n_4311;
wire n_3284;
wire n_8542;
wire n_8572;
wire n_5046;
wire n_7607;
wire n_14292;
wire n_13330;
wire n_7642;
wire n_8373;
wire n_8424;
wire n_13417;
wire n_8442;
wire n_9304;
wire n_14492;
wire n_6236;
wire n_7104;
wire n_8147;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_11152;
wire n_13505;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_10080;
wire n_2791;
wire n_3212;
wire n_11022;
wire n_4871;
wire n_11025;
wire n_12517;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_11251;
wire n_3549;
wire n_13821;
wire n_3914;
wire n_10766;
wire n_13787;
wire n_6398;
wire n_11222;
wire n_5586;
wire n_14065;
wire n_7461;
wire n_8519;
wire n_11650;
wire n_14310;
wire n_2611;
wire n_8075;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_7638;
wire n_10781;
wire n_11091;
wire n_13243;
wire n_13531;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_8642;
wire n_11713;
wire n_8648;
wire n_10217;
wire n_7224;
wire n_6966;
wire n_9791;
wire n_5056;
wire n_9449;
wire n_9934;
wire n_9149;
wire n_9686;
wire n_13063;
wire n_13186;
wire n_14639;
wire n_13463;
wire n_7259;
wire n_7838;
wire n_8556;
wire n_5984;
wire n_12961;
wire n_14039;
wire n_11398;
wire n_9844;
wire n_5204;
wire n_6705;
wire n_6724;
wire n_12389;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_11208;
wire n_9458;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_7840;
wire n_8585;
wire n_9717;
wire n_11858;
wire n_12595;
wire n_11487;
wire n_14194;
wire n_2745;
wire n_8455;
wire n_8444;
wire n_13237;
wire n_9128;
wire n_10638;
wire n_14559;
wire n_14255;
wire n_11745;
wire n_10239;
wire n_12368;
wire n_13353;
wire n_6624;
wire n_7888;
wire n_8560;
wire n_12816;
wire n_11525;
wire n_6710;
wire n_6883;
wire n_9558;
wire n_8108;
wire n_8158;
wire n_3172;
wire n_4033;
wire n_2659;
wire n_10464;
wire n_13054;
wire n_3747;
wire n_10446;
wire n_6553;
wire n_9715;
wire n_14166;
wire n_4905;
wire n_10219;
wire n_9016;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_6261;
wire n_6659;
wire n_9399;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_12967;
wire n_14458;
wire n_12907;
wire n_14353;
wire n_3116;
wire n_12020;
wire n_4141;
wire n_13877;
wire n_3784;
wire n_6893;
wire n_12377;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_3559;
wire n_12007;
wire n_13272;
wire n_11087;
wire n_8814;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_10394;
wire n_6337;
wire n_5680;
wire n_6210;
wire n_7583;
wire n_14368;
wire n_2825;
wire n_5685;
wire n_13394;
wire n_5974;
wire n_10776;
wire n_14032;
wire n_14375;
wire n_10917;
wire n_5723;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_13536;
wire n_9094;
wire n_13524;
wire n_8130;
wire n_11483;
wire n_14075;
wire n_3496;
wire n_14093;
wire n_4364;
wire n_3493;
wire n_12944;
wire n_9510;
wire n_11049;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_12706;
wire n_12973;
wire n_12319;
wire n_4307;
wire n_14178;
wire n_2795;
wire n_14053;
wire n_6044;
wire n_12388;
wire n_6206;
wire n_7893;
wire n_2954;
wire n_11031;
wire n_9429;
wire n_11599;
wire n_4438;
wire n_11292;
wire n_6538;
wire n_11568;
wire n_7966;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_9653;
wire n_4367;
wire n_5134;
wire n_11468;
wire n_13815;
wire n_7599;
wire n_9648;
wire n_7231;
wire n_14626;
wire n_10240;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_12470;
wire n_12711;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_8675;
wire n_12216;
wire n_9095;
wire n_7900;
wire n_11203;
wire n_5708;
wire n_8123;
wire n_9003;
wire n_9048;
wire n_12879;
wire n_14228;
wire n_13801;
wire n_3010;
wire n_5454;
wire n_14472;
wire n_13659;
wire n_4254;
wire n_10578;
wire n_11206;
wire n_12649;
wire n_12093;
wire n_13473;
wire n_8913;
wire n_9932;
wire n_3438;
wire n_8220;
wire n_12165;
wire n_2625;
wire n_11779;
wire n_13497;
wire n_9309;
wire n_8355;
wire n_12724;
wire n_9661;
wire n_14557;
wire n_9799;
wire n_12447;
wire n_5373;
wire n_7403;
wire n_6665;
wire n_8883;
wire n_3147;
wire n_13822;
wire n_3661;
wire n_7168;
wire n_10427;
wire n_3320;
wire n_4179;
wire n_11609;
wire n_11927;
wire n_10626;
wire n_11676;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_10138;
wire n_6860;
wire n_9063;
wire n_2919;
wire n_7322;
wire n_10364;
wire n_6060;
wire n_10532;
wire n_3108;
wire n_5983;
wire n_5788;
wire n_9895;
wire n_10288;
wire n_6709;
wire n_11602;
wire n_13843;
wire n_2632;
wire n_11865;
wire n_12566;
wire n_5557;
wire n_12383;
wire n_6914;
wire n_8816;
wire n_4314;
wire n_8418;
wire n_2980;
wire n_5951;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_12035;
wire n_3239;
wire n_2631;
wire n_12212;
wire n_9110;
wire n_3311;
wire n_11427;
wire n_3516;
wire n_11613;
wire n_4442;
wire n_10668;
wire n_4857;
wire n_8739;
wire n_9969;
wire n_11375;
wire n_8927;
wire n_10398;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_4637;
wire n_5523;
wire n_11870;
wire n_2697;
wire n_12053;
wire n_13250;
wire n_8243;
wire n_3704;
wire n_8798;
wire n_13228;
wire n_7963;
wire n_13893;
wire n_6382;
wire n_8423;
wire n_13869;
wire n_14326;
wire n_9028;
wire n_4296;
wire n_2677;
wire n_14699;
wire n_13100;
wire n_9654;
wire n_10683;
wire n_14232;
wire n_10249;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_9810;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_12852;
wire n_12123;
wire n_9701;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_9270;
wire n_11373;
wire n_11878;
wire n_3589;
wire n_6418;
wire n_8548;
wire n_9437;
wire n_8996;
wire n_13185;
wire n_9483;
wire n_6263;
wire n_14593;
wire n_6731;
wire n_8156;
wire n_5138;
wire n_8845;
wire n_4588;
wire n_6048;
wire n_13738;
wire n_7185;
wire n_10229;
wire n_12268;
wire n_5149;
wire n_9256;
wire n_4970;
wire n_5280;
wire n_3054;
wire n_10889;
wire n_11070;
wire n_6234;
wire n_4153;
wire n_8992;
wire n_5052;
wire n_5137;
wire n_3601;
wire n_7141;
wire n_11107;
wire n_14116;
wire n_3881;
wire n_13195;
wire n_12298;
wire n_6224;
wire n_12930;
wire n_8510;
wire n_5089;
wire n_11394;
wire n_5775;
wire n_9854;
wire n_3759;
wire n_9737;
wire n_8961;
wire n_12890;
wire n_14551;
wire n_9964;
wire n_11154;
wire n_3323;
wire n_4643;
wire n_9719;
wire n_6142;
wire n_10826;
wire n_2617;
wire n_6119;
wire n_10358;
wire n_12301;
wire n_13886;
wire n_6619;
wire n_11973;
wire n_13200;
wire n_2814;
wire n_4133;
wire n_11073;
wire n_13876;
wire n_2636;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_6768;
wire n_5031;
wire n_7092;
wire n_7233;
wire n_4543;
wire n_14442;
wire n_4337;
wire n_9679;
wire n_9669;
wire n_11186;
wire n_12382;
wire n_5082;
wire n_4788;
wire n_10835;
wire n_13095;
wire n_12996;
wire n_4555;
wire n_5230;
wire n_4486;
wire n_10416;
wire n_3465;
wire n_12661;
wire n_8402;
wire n_8978;
wire n_14097;
wire n_7191;
wire n_14279;
wire n_6189;
wire n_5796;
wire n_13907;
wire n_9105;
wire n_13085;
wire n_14411;
wire n_9699;
wire n_11360;
wire n_5296;
wire n_5398;
wire n_6761;
wire n_14304;
wire n_9673;
wire n_10860;
wire n_11823;
wire n_4780;
wire n_4640;
wire n_8685;
wire n_10997;
wire n_9240;
wire n_7202;
wire n_14033;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_7445;
wire n_5858;
wire n_9212;
wire n_13889;
wire n_5985;
wire n_8595;
wire n_10602;
wire n_12088;
wire n_11181;
wire n_9040;
wire n_9478;
wire n_10261;
wire n_10817;
wire n_12062;
wire n_12277;
wire n_14045;
wire n_4157;
wire n_9742;
wire n_11806;
wire n_3477;
wire n_7868;
wire n_10124;
wire n_13386;
wire n_3370;
wire n_7654;
wire n_3949;
wire n_8779;
wire n_5192;
wire n_4247;
wire n_5051;
wire n_10132;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_8520;
wire n_4583;
wire n_14305;
wire n_8555;
wire n_12421;
wire n_10730;
wire n_9456;
wire n_6366;
wire n_11321;
wire n_6304;
wire n_4292;
wire n_9146;
wire n_11702;
wire n_7176;
wire n_14233;
wire n_8565;
wire n_8334;
wire n_13605;
wire n_7547;
wire n_5552;
wire n_6074;
wire n_12133;
wire n_11970;
wire n_3764;
wire n_13283;
wire n_4773;
wire n_5028;
wire n_13596;
wire n_3025;
wire n_9573;
wire n_3051;
wire n_11286;
wire n_2802;
wire n_8030;
wire n_8513;
wire n_14511;
wire n_13746;
wire n_13327;
wire n_14550;
wire n_9379;
wire n_10948;
wire n_9219;
wire n_13534;
wire n_14056;
wire n_10927;
wire n_11496;
wire n_14151;
wire n_13149;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_8245;
wire n_13727;
wire n_13992;
wire n_7942;
wire n_4344;
wire n_5242;
wire n_12186;
wire n_3130;
wire n_8753;
wire n_7527;
wire n_9706;
wire n_4856;
wire n_2618;
wire n_7948;
wire n_7096;
wire n_11863;
wire n_4216;
wire n_9206;
wire n_2707;
wire n_14139;
wire n_8485;
wire n_5596;
wire n_6482;
wire n_10118;
wire n_8106;
wire n_2849;
wire n_8325;
wire n_2756;
wire n_3781;
wire n_14619;
wire n_10875;
wire n_4864;
wire n_11225;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_10731;
wire n_4313;
wire n_14071;
wire n_11355;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_9434;
wire n_3713;
wire n_6229;
wire n_5933;
wire n_13198;
wire n_5536;
wire n_13097;
wire n_4798;
wire n_10350;
wire n_10654;
wire n_7293;
wire n_9874;
wire n_11261;
wire n_11862;
wire n_13369;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_12579;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_5810;
wire n_3750;
wire n_10564;
wire n_3424;
wire n_12342;
wire n_13653;
wire n_3356;
wire n_14691;
wire n_11584;
wire n_9082;
wire n_7144;
wire n_12877;
wire n_3931;
wire n_12256;
wire n_4991;
wire n_11893;
wire n_10262;
wire n_13360;
wire n_11500;
wire n_11044;
wire n_7316;
wire n_7508;
wire n_13785;
wire n_9596;
wire n_3070;
wire n_8677;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_11109;
wire n_12909;
wire n_13044;
wire n_3245;
wire n_12859;
wire n_10729;
wire n_2894;
wire n_9559;
wire n_9709;
wire n_10973;
wire n_4182;
wire n_8626;
wire n_12822;
wire n_2827;
wire n_7869;
wire n_13217;
wire n_3214;
wire n_13943;
wire n_10069;
wire n_10810;
wire n_12468;
wire n_8166;
wire n_9356;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_12267;
wire n_3710;
wire n_12170;
wire n_12426;
wire n_6943;
wire n_10791;
wire n_12900;
wire n_10553;
wire n_14555;
wire n_6631;
wire n_5889;
wire n_12846;
wire n_8602;
wire n_9609;
wire n_7151;
wire n_10284;
wire n_3944;
wire n_7762;
wire n_13469;
wire n_13840;
wire n_13836;
wire n_5632;
wire n_12855;
wire n_11501;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_13569;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_9342;
wire n_14229;
wire n_4800;
wire n_14425;
wire n_7075;
wire n_13076;
wire n_5427;
wire n_12234;
wire n_4440;
wire n_4425;
wire n_6770;
wire n_14317;
wire n_5450;
wire n_7611;
wire n_11437;
wire n_7796;
wire n_6508;
wire n_14682;
wire n_7989;
wire n_13082;
wire n_8047;
wire n_12120;
wire n_13320;
wire n_2821;
wire n_3696;
wire n_9233;
wire n_10474;
wire n_7936;
wire n_10694;
wire n_10529;
wire n_13117;
wire n_4781;
wire n_12042;
wire n_6031;
wire n_3531;
wire n_14328;
wire n_5124;
wire n_4237;
wire n_8751;
wire n_5297;
wire n_11722;
wire n_4828;
wire n_3333;
wire n_12568;
wire n_12149;
wire n_14444;
wire n_8800;
wire n_4652;
wire n_12278;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_10622;
wire n_9435;
wire n_3135;
wire n_13318;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_9557;
wire n_11639;
wire n_9551;
wire n_8955;
wire n_8039;
wire n_8193;
wire n_12116;
wire n_12231;
wire n_9073;
wire n_13677;
wire n_7546;
wire n_8432;
wire n_14422;
wire n_5904;
wire n_11997;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_8684;
wire n_10270;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_13158;
wire n_7407;
wire n_12014;
wire n_13230;
wire n_9388;
wire n_3277;
wire n_10463;
wire n_9721;
wire n_11731;
wire n_14061;
wire n_4863;
wire n_10880;
wire n_11610;
wire n_12097;
wire n_14612;
wire n_12363;
wire n_13115;
wire n_13427;
wire n_5463;
wire n_2978;
wire n_6328;
wire n_11498;
wire n_6929;
wire n_12008;
wire n_11509;
wire n_4859;
wire n_4568;
wire n_8628;
wire n_14401;
wire n_14034;
wire n_13559;
wire n_3617;
wire n_6012;
wire n_2958;
wire n_7481;
wire n_11447;
wire n_4429;
wire n_6484;
wire n_5435;
wire n_11706;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_11055;
wire n_14498;
wire n_10689;
wire n_9507;
wire n_5476;
wire n_5483;
wire n_12534;
wire n_9539;
wire n_8617;
wire n_14297;
wire n_14517;
wire n_7605;
wire n_8591;
wire n_8090;
wire n_9268;
wire n_5511;
wire n_9718;
wire n_8661;
wire n_13512;
wire n_10068;
wire n_3486;
wire n_6639;
wire n_11258;
wire n_9672;
wire n_12748;
wire n_11168;
wire n_9890;
wire n_12272;
wire n_9187;
wire n_9572;
wire n_12148;
wire n_2992;
wire n_10363;
wire n_6124;
wire n_12142;
wire n_12615;
wire n_13201;
wire n_9527;
wire n_3197;
wire n_11234;
wire n_9949;
wire n_13388;
wire n_14484;
wire n_7423;
wire n_13674;
wire n_3256;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_8189;
wire n_8811;
wire n_13858;
wire n_9952;
wire n_11612;
wire n_7736;
wire n_6435;
wire n_13949;
wire n_10888;
wire n_12714;
wire n_13782;
wire n_14486;
wire n_3646;
wire n_5829;
wire n_14580;
wire n_7419;
wire n_13612;
wire n_6600;
wire n_14087;
wire n_13681;
wire n_7010;
wire n_13700;
wire n_14421;
wire n_14193;
wire n_10277;
wire n_5881;
wire n_9798;
wire n_3864;
wire n_4694;
wire n_11895;
wire n_8192;
wire n_9251;
wire n_4664;
wire n_6201;
wire n_10537;
wire n_14684;
wire n_3450;
wire n_14653;
wire n_8573;
wire n_14703;
wire n_4633;
wire n_13770;
wire n_10807;
wire n_4050;
wire n_3173;
wire n_14048;
wire n_13920;
wire n_7918;
wire n_9546;
wire n_10331;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_13130;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_9602;
wire n_9181;
wire n_12812;
wire n_3266;
wire n_3102;
wire n_13377;
wire n_11455;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_10981;
wire n_5894;
wire n_13750;
wire n_9635;
wire n_11868;
wire n_4511;
wire n_3422;
wire n_12189;
wire n_12639;
wire n_14063;
wire n_14343;
wire n_14521;
wire n_4675;
wire n_13701;
wire n_11934;
wire n_13518;
wire n_2991;
wire n_5419;
wire n_8339;
wire n_11969;
wire n_13668;
wire n_4289;
wire n_4972;
wire n_11571;
wire n_2723;
wire n_6036;
wire n_7346;
wire n_9405;
wire n_3925;
wire n_12428;
wire n_12069;
wire n_14384;
wire n_4689;
wire n_5165;
wire n_8775;
wire n_10780;
wire n_10158;
wire n_11481;
wire n_2850;
wire n_5077;
wire n_6102;
wire n_14276;
wire n_12057;
wire n_3780;
wire n_12050;
wire n_13587;
wire n_9726;
wire n_13488;
wire n_8804;
wire n_9577;
wire n_6650;
wire n_10024;
wire n_6573;
wire n_11774;
wire n_6904;
wire n_12214;
wire n_3753;
wire n_6329;
wire n_13805;
wire n_7385;
wire n_9802;
wire n_6244;
wire n_4846;
wire n_9540;
wire n_6204;
wire n_9250;
wire n_13365;
wire n_13767;
wire n_13972;
wire n_12381;
wire n_10191;
wire n_5225;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_12157;
wire n_7148;
wire n_13938;
wire n_3142;
wire n_9171;
wire n_7169;
wire n_3129;
wire n_13443;
wire n_9350;
wire n_3495;
wire n_3843;
wire n_11257;
wire n_12330;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_9441;
wire n_7600;
wire n_9124;
wire n_10675;
wire n_5826;
wire n_8697;
wire n_11598;
wire n_9626;
wire n_14011;
wire n_14645;
wire n_4822;
wire n_11327;
wire n_6946;
wire n_12926;
wire n_7947;
wire n_8645;
wire n_5931;
wire n_8820;
wire n_8146;
wire n_9408;
wire n_4635;
wire n_8154;
wire n_7847;
wire n_12824;
wire n_12392;
wire n_13094;
wire n_5532;
wire n_14545;
wire n_7311;
wire n_6804;
wire n_3740;
wire n_5441;
wire n_6179;
wire n_14103;
wire n_6059;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_2911;
wire n_8063;
wire n_3313;
wire n_13798;
wire n_14677;
wire n_8406;
wire n_6427;
wire n_14474;
wire n_14459;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_12070;
wire n_3726;
wire n_8480;
wire n_11265;
wire n_14037;
wire n_11788;
wire n_14112;
wire n_9754;
wire n_10477;
wire n_4419;
wire n_14296;
wire n_11904;
wire n_8849;
wire n_13071;
wire n_5405;
wire n_9750;
wire n_10296;
wire n_7660;
wire n_13676;
wire n_13735;
wire n_14127;
wire n_5365;
wire n_9566;
wire n_5772;
wire n_3345;
wire n_3560;
wire n_9529;
wire n_10339;
wire n_11901;
wire n_12848;
wire n_6442;
wire n_8241;
wire n_10307;
wire n_10606;
wire n_6188;
wire n_12161;
wire n_3421;
wire n_10066;
wire n_11755;
wire n_4906;
wire n_3548;
wire n_11754;
wire n_6846;
wire n_13825;
wire n_10054;
wire n_4630;
wire n_8261;
wire n_10343;
wire n_6840;
wire n_6645;
wire n_8535;
wire n_8348;
wire n_4829;
wire n_13985;
wire n_6749;
wire n_12238;
wire n_6915;
wire n_12956;
wire n_12320;
wire n_7831;
wire n_8138;
wire n_13342;
wire n_2612;
wire n_11413;
wire n_13953;
wire n_10652;
wire n_13040;
wire n_5259;
wire n_3236;
wire n_8702;
wire n_11601;
wire n_7455;
wire n_8273;
wire n_14250;
wire n_10944;
wire n_6247;
wire n_5921;
wire n_10367;
wire n_11129;
wire n_11710;
wire n_4966;
wire n_14602;
wire n_8235;
wire n_13685;
wire n_6104;
wire n_3321;
wire n_9940;
wire n_8294;
wire n_12476;
wire n_4188;
wire n_10016;
wire n_9036;
wire n_9165;
wire n_7509;
wire n_9283;
wire n_6205;
wire n_11010;
wire n_8349;
wire n_4825;
wire n_2610;
wire n_3715;
wire n_9822;
wire n_10036;
wire n_2626;
wire n_9443;
wire n_9607;
wire n_7497;
wire n_10749;
wire n_7315;
wire n_10166;
wire n_8429;
wire n_13765;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_7887;
wire n_10419;
wire n_2804;
wire n_9298;
wire n_5884;
wire n_5006;
wire n_14200;
wire n_4882;
wire n_3206;
wire n_10006;
wire n_5728;
wire n_13334;
wire n_3475;
wire n_4878;
wire n_8486;
wire n_11240;
wire n_9052;
wire n_6706;
wire n_13123;
wire n_12154;
wire n_7431;
wire n_8140;
wire n_11734;
wire n_14450;
wire n_3842;
wire n_12645;
wire n_14477;
wire n_4202;
wire n_6909;
wire n_13933;
wire n_5679;
wire n_6487;
wire n_8117;
wire n_12668;
wire n_3886;
wire n_10348;
wire n_13884;
wire n_2619;
wire n_7521;
wire n_10058;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_8129;
wire n_10355;
wire n_11156;
wire n_7253;
wire n_5208;
wire n_9535;
wire n_13511;
wire n_5113;
wire n_10304;
wire n_12928;
wire n_3987;
wire n_11955;
wire n_5205;
wire n_4249;
wire n_9943;
wire n_7569;
wire n_12538;
wire n_13745;
wire n_12151;
wire n_3160;
wire n_10966;
wire n_14697;
wire n_13112;
wire n_2968;
wire n_13646;
wire n_12130;
wire n_14608;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_12409;
wire n_13031;
wire n_6551;
wire n_3386;
wire n_12350;
wire n_7972;
wire n_8672;
wire n_13455;
wire n_7505;
wire n_13993;
wire n_3921;
wire n_14280;
wire n_13946;
wire n_6516;
wire n_14567;
wire n_2766;
wire n_10060;
wire n_7524;
wire n_13931;
wire n_4196;
wire n_11270;
wire n_8934;
wire n_11020;
wire n_7318;
wire n_2613;
wire n_9977;
wire n_10722;
wire n_7411;
wire n_13314;
wire n_7326;
wire n_13378;
wire n_5667;
wire n_9555;
wire n_13618;
wire n_10957;
wire n_2647;
wire n_14277;
wire n_8847;
wire n_8005;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_11344;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_6500;
wire n_11303;
wire n_5027;
wire n_12847;
wire n_3380;
wire n_14340;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_9030;
wire n_11216;
wire n_8221;
wire n_13638;
wire n_7573;
wire n_6630;
wire n_5759;
wire n_5629;
wire n_10409;
wire n_13167;
wire n_4631;
wire n_8191;
wire n_6798;
wire n_13758;
wire n_5999;
wire n_9590;
wire n_14646;
wire n_11511;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_10322;
wire n_11339;
wire n_11346;
wire n_11829;
wire n_12680;
wire n_5377;
wire n_6180;
wire n_12530;
wire n_11581;
wire n_8225;
wire n_3822;
wire n_7453;
wire n_4355;
wire n_3818;
wire n_12163;
wire n_14131;
wire n_7932;
wire n_9651;
wire n_7890;
wire n_5599;
wire n_10825;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_9583;
wire n_9944;
wire n_9763;
wire n_10349;
wire n_13709;
wire n_13035;
wire n_6652;
wire n_9888;
wire n_7183;
wire n_4155;
wire n_4278;
wire n_10040;
wire n_10636;
wire n_4710;
wire n_10844;
wire n_12738;
wire n_6275;
wire n_6403;
wire n_3497;
wire n_6395;
wire n_9862;
wire n_14622;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_9966;
wire n_10242;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_9936;
wire n_3927;
wire n_6141;
wire n_8559;
wire n_11165;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_9617;
wire n_10727;
wire n_4060;
wire n_9341;
wire n_6194;
wire n_8689;
wire n_11231;
wire n_3396;
wire n_9749;
wire n_5517;
wire n_9629;
wire n_13654;
wire n_5807;
wire n_11448;
wire n_12227;
wire n_5426;
wire n_6475;
wire n_12525;
wire n_10679;
wire n_4093;
wire n_11132;
wire n_10524;
wire n_12282;
wire n_5693;
wire n_13426;
wire n_5695;
wire n_12932;
wire n_4123;
wire n_13799;
wire n_14207;
wire n_4294;
wire n_8330;
wire n_10011;
wire n_12037;
wire n_3683;
wire n_6502;
wire n_10030;
wire n_6944;
wire n_11410;
wire n_14365;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_8304;
wire n_9349;
wire n_13480;
wire n_5587;
wire n_4722;
wire n_11267;
wire n_13780;
wire n_6318;
wire n_10119;
wire n_11348;
wire n_11940;
wire n_13613;
wire n_10845;
wire n_8163;
wire n_6805;
wire n_11947;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_7240;
wire n_8907;
wire n_2963;
wire n_14227;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_9423;
wire n_5584;
wire n_12424;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_6075;
wire n_10063;
wire n_12942;
wire n_6559;
wire n_4088;
wire n_9038;
wire n_8777;
wire n_11149;
wire n_2669;
wire n_8698;
wire n_10709;
wire n_6068;
wire n_3911;
wire n_3802;
wire n_12236;
wire n_4366;
wire n_6248;
wire n_6541;
wire n_11436;
wire n_9034;
wire n_5125;
wire n_4922;
wire n_11909;
wire n_12547;
wire n_13554;
wire n_6066;
wire n_6080;
wire n_14372;
wire n_13421;
wire n_4733;
wire n_7927;
wire n_8928;
wire n_13967;
wire n_13150;
wire n_13014;
wire n_7219;
wire n_10526;
wire n_11439;
wire n_8081;
wire n_12192;
wire n_4041;
wire n_12747;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_6638;
wire n_11462;
wire n_14564;
wire n_7063;
wire n_7402;
wire n_9676;
wire n_6351;
wire n_4509;
wire n_4935;
wire n_7382;
wire n_10861;
wire n_8384;
wire n_13795;
wire n_5238;
wire n_4004;
wire n_8650;
wire n_3630;
wire n_11272;
wire n_14044;
wire n_12989;
wire n_5906;
wire n_7767;
wire n_5732;
wire n_4194;
wire n_2672;
wire n_11759;
wire n_10494;
wire n_14431;
wire n_2602;
wire n_5780;
wire n_10478;
wire n_11061;
wire n_11653;
wire n_2931;
wire n_3433;
wire n_8284;
wire n_10534;
wire n_8374;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_13662;
wire n_13864;
wire n_5743;
wire n_6481;
wire n_10078;
wire n_5633;
wire n_4111;
wire n_11478;
wire n_7510;
wire n_12273;
wire n_9041;
wire n_3786;
wire n_9995;
wire n_12200;
wire n_6022;
wire n_6991;
wire n_10629;
wire n_2828;
wire n_13863;
wire n_7434;
wire n_5950;
wire n_9035;
wire n_13926;
wire n_9011;
wire n_14240;
wire n_4204;
wire n_7691;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_11748;
wire n_14165;
wire n_9135;
wire n_6744;
wire n_3645;
wire n_9776;
wire n_5705;
wire n_12660;
wire n_11867;
wire n_14192;
wire n_6927;
wire n_14678;
wire n_7335;
wire n_12400;
wire n_13072;
wire n_10472;
wire n_10695;
wire n_10286;
wire n_9413;
wire n_4996;
wire n_9107;
wire n_4411;
wire n_2883;
wire n_4317;
wire n_7735;
wire n_8531;
wire n_6116;
wire n_9548;
wire n_8074;
wire n_14246;
wire n_3550;
wire n_8780;
wire n_7956;
wire n_5510;
wire n_7495;
wire n_7651;
wire n_4785;
wire n_2870;
wire n_9775;
wire n_13857;
wire n_12922;
wire n_13033;
wire n_8580;
wire n_4068;
wire n_5440;
wire n_12193;
wire n_9288;
wire n_4163;
wire n_3294;
wire n_3610;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_3279;
wire n_12243;
wire n_5513;
wire n_10218;
wire n_5875;
wire n_14671;
wire n_8358;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_10441;
wire n_2843;
wire n_3714;
wire n_9305;
wire n_9093;
wire n_11764;
wire n_7671;
wire n_13696;
wire n_12950;
wire n_10043;
wire n_4832;
wire n_8033;
wire n_3676;
wire n_5197;
wire n_6485;
wire n_13041;
wire n_5848;
wire n_5834;
wire n_14269;
wire n_7926;
wire n_3109;
wire n_11882;
wire n_5784;
wire n_13418;
wire n_3125;
wire n_12250;
wire n_5128;
wire n_10628;
wire n_13498;
wire n_14290;
wire n_8643;
wire n_11787;
wire n_12403;
wire n_5618;
wire n_11539;
wire n_10440;
wire n_10134;
wire n_12904;
wire n_6495;
wire n_7528;
wire n_14669;
wire n_12444;
wire n_11163;
wire n_6209;
wire n_4672;
wire n_8094;
wire n_2564;
wire n_3558;
wire n_11695;
wire n_9425;
wire n_13489;
wire n_14520;
wire n_13373;
wire n_3034;
wire n_10317;
wire n_13739;
wire n_11730;
wire n_13101;
wire n_11916;
wire n_13723;
wire n_3502;
wire n_13000;
wire n_13556;
wire n_4053;
wire n_11311;
wire n_14525;
wire n_7413;
wire n_14435;
wire n_7993;
wire n_11980;
wire n_7821;
wire n_11151;
wire n_14238;
wire n_7620;
wire n_3963;
wire n_13153;
wire n_12837;
wire n_12356;
wire n_3091;
wire n_13091;
wire n_13937;
wire n_13032;
wire n_6274;
wire n_5157;
wire n_12764;
wire n_14654;
wire n_4496;
wire n_9347;
wire n_12269;
wire n_14556;
wire n_12079;
wire n_14687;
wire n_13508;
wire n_10706;
wire n_4596;
wire n_5178;
wire n_9420;
wire n_13350;
wire n_13901;
wire n_12972;
wire n_3105;
wire n_6237;
wire n_13635;
wire n_4628;
wire n_6802;
wire n_13224;
wire n_7343;
wire n_5982;
wire n_8477;
wire n_13306;
wire n_9344;
wire n_14657;
wire n_7109;
wire n_12438;
wire n_8028;
wire n_14245;
wire n_14254;
wire n_12125;
wire n_4083;
wire n_12554;
wire n_10297;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_9530;
wire n_6809;
wire n_10160;
wire n_6099;
wire n_10849;
wire n_3225;
wire n_10605;
wire n_11296;
wire n_13259;
wire n_8530;
wire n_14217;
wire n_10379;
wire n_9446;
wire n_3621;
wire n_5529;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_11081;
wire n_8500;
wire n_13278;
wire n_6716;
wire n_8713;
wire n_12860;
wire n_3565;
wire n_7885;
wire n_14554;
wire n_8297;
wire n_14100;
wire n_6905;
wire n_8926;
wire n_9865;
wire n_8456;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_11230;
wire n_5824;
wire n_8025;
wire n_10282;
wire n_5354;
wire n_7898;
wire n_11357;
wire n_3331;
wire n_11027;
wire n_13179;
wire n_10458;
wire n_12206;
wire n_11393;
wire n_6203;
wire n_12947;
wire n_6407;
wire n_14468;
wire n_4230;
wire n_3040;
wire n_11892;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_3360;
wire n_3585;
wire n_7070;
wire n_9025;
wire n_5276;
wire n_11105;
wire n_4037;
wire n_9713;
wire n_11160;
wire n_13043;
wire n_3804;
wire n_14675;
wire n_4659;
wire n_8293;
wire n_13962;
wire n_3211;
wire n_7299;
wire n_5196;
wire n_10382;
wire n_2556;
wire n_8029;
wire n_13468;
wire n_9314;
wire n_3847;
wire n_12270;
wire n_6960;
wire n_4073;
wire n_14235;
wire n_8880;
wire n_7249;
wire n_9660;
wire n_5763;
wire n_3633;
wire n_13018;
wire n_12739;
wire n_6061;
wire n_13831;
wire n_9769;
wire n_4001;
wire n_2584;
wire n_8471;
wire n_5701;
wire n_7002;
wire n_14529;
wire n_12906;
wire n_12490;
wire n_9902;
wire n_6273;
wire n_14424;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_12751;
wire n_11397;
wire n_8726;
wire n_10640;
wire n_8977;
wire n_2997;
wire n_7018;
wire n_11897;
wire n_10522;
wire n_6746;
wire n_3258;
wire n_10691;
wire n_12650;
wire n_10764;
wire n_10244;
wire n_10914;
wire n_13348;
wire n_3691;
wire n_8316;
wire n_6174;
wire n_10272;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_14690;
wire n_13415;
wire n_5907;
wire n_4339;
wire n_7297;
wire n_7730;
wire n_10980;
wire n_12279;
wire n_13265;
wire n_8134;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_5895;
wire n_9410;
wire n_9588;
wire n_2651;
wire n_12242;
wire n_2733;
wire n_4169;
wire n_4024;
wire n_3316;
wire n_8610;
wire n_4023;
wire n_10071;
wire n_4253;
wire n_7637;
wire n_3632;
wire n_12588;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_13382;
wire n_10176;
wire n_6113;
wire n_9740;
wire n_3457;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_6575;
wire n_11719;
wire n_5283;
wire n_9910;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_7613;
wire n_9061;
wire n_7995;
wire n_9941;
wire n_8113;
wire n_9579;
wire n_5686;
wire n_6391;
wire n_10254;
wire n_2740;
wire n_14446;
wire n_8724;
wire n_14121;
wire n_10332;
wire n_7140;
wire n_12775;
wire n_12173;
wire n_4066;
wire n_10938;
wire n_10257;
wire n_9668;
wire n_6252;
wire n_6426;
wire n_14031;
wire n_4681;
wire n_12167;
wire n_8253;
wire n_11956;
wire n_9258;
wire n_9228;
wire n_3303;
wire n_13461;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_10214;
wire n_11874;
wire n_5094;
wire n_10195;
wire n_3232;
wire n_13979;
wire n_9598;
wire n_10354;
wire n_7741;
wire n_12060;
wire n_3768;
wire n_4295;
wire n_10436;
wire n_11450;
wire n_4100;
wire n_11723;
wire n_6668;
wire n_9311;
wire n_11982;
wire n_14062;
wire n_3445;
wire n_12179;
wire n_11822;
wire n_14448;
wire n_11522;
wire n_4087;
wire n_8232;
wire n_12842;
wire n_8803;
wire n_10866;
wire n_4473;
wire n_4619;
wire n_12499;
wire n_6670;
wire n_5371;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_8818;
wire n_12693;
wire n_10811;
wire n_7698;
wire n_10073;
wire n_6962;
wire n_14187;
wire n_6779;
wire n_9608;
wire n_5286;
wire n_10164;
wire n_4449;
wire n_13172;
wire n_3285;
wire n_4607;
wire n_10205;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_10515;
wire n_7800;
wire n_12326;
wire n_4266;
wire n_6336;
wire n_13713;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_12542;
wire n_13650;
wire n_6049;
wire n_5885;
wire n_11499;
wire n_3628;
wire n_14390;
wire n_9818;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_11034;
wire n_7415;
wire n_8823;
wire n_5399;
wire n_8536;
wire n_9433;
wire n_14004;
wire n_11746;
wire n_11698;
wire n_8795;
wire n_2846;
wire n_3371;
wire n_10430;
wire n_12934;
wire n_10338;
wire n_11560;
wire n_9599;
wire n_8674;
wire n_9186;
wire n_14054;
wire n_4918;
wire n_5856;
wire n_8016;
wire n_13941;
wire n_3872;
wire n_5760;
wire n_12483;
wire n_7747;
wire n_9935;
wire n_14263;
wire n_12404;
wire n_12258;
wire n_4415;
wire n_5110;
wire n_8966;
wire n_11871;
wire n_14694;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_10018;
wire n_9537;
wire n_10500;
wire n_9552;
wire n_9421;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_13209;
wire n_5844;
wire n_10359;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_3441;
wire n_3020;
wire n_12823;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_6609;
wire n_10548;
wire n_7635;
wire n_4408;
wire n_12905;
wire n_10291;
wire n_8567;
wire n_8259;
wire n_10667;
wire n_12274;
wire n_12849;
wire n_11167;
wire n_11297;
wire n_4976;
wire n_9473;
wire n_6525;
wire n_10208;
wire n_11183;
wire n_3555;
wire n_9469;
wire n_11285;
wire n_5938;
wire n_14270;
wire n_7274;
wire n_3534;
wire n_11740;
wire n_8578;
wire n_10757;
wire n_4548;
wire n_7819;
wire n_8495;
wire n_14679;
wire n_2670;
wire n_13975;
wire n_6494;
wire n_3556;
wire n_4574;
wire n_8160;
wire n_8980;
wire n_2644;
wire n_6132;
wire n_10631;
wire n_10864;
wire n_11136;
wire n_4557;
wire n_3071;
wire n_11434;
wire n_8336;
wire n_11133;
wire n_13711;
wire n_5548;
wire n_7788;
wire n_6974;
wire n_13477;
wire n_10748;
wire n_4663;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_9909;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_12303;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_12002;
wire n_8600;
wire n_8229;
wire n_12442;
wire n_4686;
wire n_9236;
wire n_9751;
wire n_10751;
wire n_14649;
wire n_7794;
wire n_13579;
wire n_3707;
wire n_3895;
wire n_10434;
wire n_9369;
wire n_3149;
wire n_3934;
wire n_13634;
wire n_4338;
wire n_13987;
wire n_12597;
wire n_5917;
wire n_9757;
wire n_12419;
wire n_6965;
wire n_11886;
wire n_3231;
wire n_14210;
wire n_8761;
wire n_14316;
wire n_7630;
wire n_11804;
wire n_13262;
wire n_4161;
wire n_14673;
wire n_9076;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_3058;
wire n_5355;
wire n_9729;
wire n_3709;
wire n_3398;
wire n_11531;
wire n_12943;
wire n_13543;
wire n_6284;
wire n_3592;
wire n_12039;
wire n_10663;
wire n_14393;
wire n_5321;
wire n_14144;
wire n_7454;
wire n_10263;
wire n_12295;
wire n_3399;
wire n_8473;
wire n_9366;
wire n_4772;
wire n_11883;
wire n_6931;
wire n_6521;
wire n_8351;
wire n_5915;
wire n_7276;
wire n_11792;
wire n_6379;
wire n_9647;
wire n_12410;
wire n_7085;
wire n_6306;
wire n_12938;
wire n_4120;
wire n_7753;
wire n_12891;
wire n_13493;
wire n_12304;
wire n_6834;
wire n_2880;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_8948;
wire n_13166;
wire n_13541;
wire n_12572;
wire n_10318;
wire n_13551;
wire n_14356;
wire n_5116;
wire n_3771;
wire n_10740;
wire n_7225;
wire n_11634;
wire n_7541;
wire n_3158;
wire n_11039;
wire n_3221;
wire n_10062;
wire n_7913;
wire n_10128;
wire n_8020;
wire n_7946;
wire n_8944;
wire n_2830;
wire n_10717;
wire n_11965;
wire n_5500;
wire n_13890;
wire n_9275;
wire n_4622;
wire n_4757;
wire n_9520;
wire n_6949;
wire n_6471;
wire n_11477;
wire n_5669;
wire n_5672;
wire n_5621;
wire n_3334;
wire n_4016;
wire n_9493;
wire n_6760;
wire n_2940;
wire n_3427;
wire n_8875;
wire n_3162;
wire n_5966;
wire n_4591;
wire n_5569;
wire n_9102;
wire n_14128;
wire n_5515;
wire n_11588;
wire n_11818;
wire n_6589;
wire n_11592;
wire n_3083;
wire n_4570;
wire n_10721;
wire n_7014;
wire n_10945;
wire n_12290;
wire n_9801;
wire n_11742;
wire n_13902;
wire n_12718;
wire n_7920;
wire n_11312;
wire n_5559;
wire n_8649;
wire n_5337;
wire n_11235;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_14185;
wire n_7841;
wire n_9424;
wire n_10013;
wire n_7324;
wire n_7160;
wire n_9333;
wire n_8205;
wire n_11505;
wire n_12469;
wire n_6046;
wire n_11673;
wire n_7054;
wire n_4493;
wire n_8975;
wire n_6055;
wire n_7161;
wire n_9004;
wire n_6364;
wire n_8919;
wire n_6091;
wire n_6348;
wire n_9987;
wire n_8440;
wire n_11555;
wire n_13917;
wire n_4896;
wire n_8041;
wire n_4851;
wire n_6848;
wire n_9860;
wire n_10565;
wire n_14327;
wire n_7837;
wire n_9670;
wire n_6788;
wire n_13548;
wire n_13903;
wire n_11241;
wire n_6144;
wire n_10389;
wire n_9200;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_12336;
wire n_13080;
wire n_9417;
wire n_11059;
wire n_6896;
wire n_5753;
wire n_8076;
wire n_5358;
wire n_12248;
wire n_12931;
wire n_14047;
wire n_11066;
wire n_4901;
wire n_3480;
wire n_8757;
wire n_10020;
wire n_7201;
wire n_13408;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_9386;
wire n_12713;
wire n_8897;
wire n_12810;
wire n_7676;
wire n_8177;
wire n_11683;
wire n_13733;
wire n_14311;
wire n_5467;
wire n_7241;
wire n_3181;
wire n_14147;
wire n_5493;
wire n_9207;
wire n_13592;
wire n_6285;
wire n_10356;
wire n_12717;
wire n_13915;
wire n_7644;
wire n_9276;
wire n_4602;
wire n_7816;
wire n_8829;
wire n_12119;
wire n_14186;
wire n_2818;
wire n_14149;
wire n_4900;
wire n_10110;
wire n_3578;
wire n_3745;
wire n_6748;
wire n_11275;
wire n_7430;
wire n_14540;
wire n_13589;
wire n_3487;
wire n_3668;
wire n_11329;
wire n_8638;
wire n_14272;
wire n_13189;
wire n_13260;
wire n_5901;
wire n_9980;
wire n_2837;
wire n_11923;
wire n_11718;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_10501;
wire n_7269;
wire n_12003;
wire n_7047;
wire n_2671;
wire n_12292;
wire n_2702;
wire n_10908;
wire n_9176;
wire n_6937;
wire n_4363;
wire n_12405;
wire n_3561;
wire n_9728;
wire n_11809;
wire n_4103;
wire n_10777;
wire n_8101;
wire n_13712;
wire n_5439;
wire n_8687;
wire n_6115;
wire n_3154;
wire n_9866;
wire n_14685;
wire n_8721;
wire n_8749;
wire n_12780;
wire n_13349;
wire n_9465;
wire n_13277;
wire n_3938;
wire n_11975;
wire n_8937;
wire n_6272;
wire n_7067;
wire n_12087;
wire n_13233;
wire n_13808;
wire n_14478;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_12662;
wire n_10965;
wire n_4416;
wire n_7879;
wire n_8730;
wire n_11441;
wire n_12416;
wire n_9702;
wire n_10998;
wire n_13503;
wire n_6607;
wire n_12854;
wire n_4439;
wire n_4985;
wire n_12936;
wire n_9000;
wire n_13056;
wire n_3382;
wire n_13300;
wire n_7117;
wire n_11743;
wire n_3930;
wire n_3808;
wire n_12765;
wire n_9610;
wire n_5471;
wire n_13087;
wire n_4660;
wire n_8503;
wire n_10082;
wire n_10870;
wire n_12796;
wire n_11914;
wire n_3081;
wire n_6446;
wire n_10756;
wire n_5497;
wire n_9139;
wire n_13287;
wire n_5519;
wire n_6071;
wire n_2579;
wire n_12028;
wire n_8315;
wire n_11175;
wire n_10411;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_6807;
wire n_2844;
wire n_11753;
wire n_8197;
wire n_13726;
wire n_11790;
wire n_9407;
wire n_12294;
wire n_6616;
wire n_6719;
wire n_14621;
wire n_10423;
wire n_4814;
wire n_8019;
wire n_8801;
wire n_12190;
wire n_14396;
wire n_6178;
wire n_11249;
wire n_8707;
wire n_6677;
wire n_11791;
wire n_12786;
wire n_7875;
wire n_5502;
wire n_8962;
wire n_13665;
wire n_8931;
wire n_8248;
wire n_14177;
wire n_7550;
wire n_14533;
wire n_8554;
wire n_2838;
wire n_13242;
wire n_11879;
wire n_13900;
wire n_10782;
wire n_13837;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_12386;
wire n_13121;
wire n_13680;
wire n_13679;
wire n_9357;
wire n_9477;
wire n_11911;
wire n_13734;
wire n_14591;
wire n_7238;
wire n_6862;
wire n_8501;
wire n_3657;
wire n_5706;
wire n_11842;
wire n_12746;
wire n_14023;
wire n_2634;
wire n_13047;
wire n_11304;
wire n_11320;
wire n_2746;
wire n_7292;
wire n_13146;
wire n_7804;
wire n_10251;
wire n_12128;
wire n_11776;
wire n_14544;
wire n_11471;
wire n_5098;
wire n_13475;
wire n_6000;
wire n_6774;
wire n_9289;
wire n_11794;
wire n_6443;
wire n_9828;
wire n_8263;
wire n_5145;
wire n_6072;
wire n_13236;
wire n_2878;
wire n_7248;
wire n_10737;
wire n_3830;
wire n_10475;
wire n_3252;
wire n_6647;
wire n_11198;
wire n_8040;
wire n_13336;
wire n_5466;
wire n_14465;
wire n_6941;
wire n_7239;
wire n_9797;
wire n_6552;
wire n_7826;
wire n_10665;
wire n_9981;
wire n_3315;
wire n_6094;
wire n_12761;
wire n_14482;
wire n_3523;
wire n_12113;
wire n_8102;
wire n_3999;
wire n_14440;
wire n_10541;
wire n_13393;
wire n_9793;
wire n_11419;
wire n_14214;
wire n_13202;
wire n_8196;
wire n_11171;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_8822;
wire n_5213;
wire n_12017;
wire n_3474;
wire n_5738;
wire n_14483;
wire n_9514;
wire n_7971;
wire n_12139;
wire n_8885;
wire n_11564;
wire n_5592;
wire n_11078;
wire n_5620;
wire n_12802;
wire n_3150;
wire n_5491;
wire n_10633;
wire n_4831;
wire n_12592;
wire n_4782;
wire n_9825;
wire n_2859;
wire n_10573;
wire n_5216;
wire n_3412;
wire n_11218;
wire n_5953;
wire n_8474;
wire n_5703;
wire n_10258;
wire n_6886;
wire n_7078;
wire n_4597;
wire n_12791;
wire n_9501;
wire n_12352;
wire n_13811;
wire n_12296;
wire n_11459;
wire n_9043;
wire n_8152;
wire n_12491;
wire n_11998;
wire n_8269;
wire n_4546;
wire n_11775;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_11288;
wire n_4147;
wire n_12454;
wire n_10042;
wire n_12162;
wire n_10570;
wire n_13151;
wire n_3073;
wire n_6531;
wire n_9481;
wire n_3571;
wire n_11768;
wire n_7577;
wire n_4576;
wire n_12992;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_11456;
wire n_11708;
wire n_14330;
wire n_12960;
wire n_8144;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_11662;
wire n_13617;
wire n_7513;
wire n_10098;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_9351;
wire n_9766;
wire n_13935;
wire n_13930;
wire n_6935;
wire n_2899;
wire n_6984;
wire n_10106;
wire n_6778;
wire n_8058;
wire n_11877;
wire n_12046;
wire n_8909;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_5526;
wire n_3877;
wire n_5202;
wire n_12074;
wire n_14380;
wire n_3817;
wire n_6345;
wire n_9242;
wire n_10754;
wire n_6386;
wire n_2722;
wire n_6596;
wire n_3728;
wire n_12749;
wire n_14630;
wire n_5107;
wire n_7165;
wire n_9777;
wire n_4680;
wire n_5067;
wire n_11932;
wire n_11821;
wire n_12485;
wire n_14464;
wire n_9522;
wire n_14560;
wire n_6830;
wire n_2685;
wire n_9748;
wire n_5987;
wire n_12488;
wire n_14028;
wire n_12252;
wire n_10851;
wire n_9005;
wire n_12090;
wire n_11395;
wire n_2788;
wire n_10387;
wire n_6642;
wire n_6291;
wire n_9666;
wire n_6510;
wire n_10615;
wire n_5264;
wire n_14081;
wire n_14281;
wire n_2595;
wire n_10790;
wire n_3084;
wire n_10028;
wire n_10555;
wire n_12896;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_11532;
wire n_8024;
wire n_7123;
wire n_14670;
wire n_4562;
wire n_3860;
wire n_10222;
wire n_2909;
wire n_3554;
wire n_12868;
wire n_6509;
wire n_10671;
wire n_2717;
wire n_6376;
wire n_8107;
wire n_9605;
wire n_2981;
wire n_10498;
wire n_13959;
wire n_9947;
wire n_9930;
wire n_13292;
wire n_4995;
wire n_5873;
wire n_6514;
wire n_10420;
wire n_4498;
wire n_6741;
wire n_10083;
wire n_10520;
wire n_6434;
wire n_9662;
wire n_5741;
wire n_2743;
wire n_2969;
wire n_3429;
wire n_9768;
wire n_6593;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_12583;
wire n_8748;
wire n_14420;
wire n_8452;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_3485;
wire n_4109;
wire n_10255;
wire n_8742;
wire n_3777;
wire n_8393;
wire n_9835;
wire n_11117;
wire n_11494;
wire n_9656;
wire n_11643;
wire n_14613;
wire n_3767;
wire n_12462;
wire n_12618;
wire n_14090;
wire n_14604;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_9475;
wire n_3692;
wire n_3234;
wire n_14347;
wire n_11475;
wire n_8122;
wire n_11004;
wire n_9724;
wire n_6947;
wire n_8403;
wire n_8912;
wire n_10612;
wire n_4850;
wire n_10007;
wire n_9154;
wire n_12127;
wire n_13651;
wire n_3716;
wire n_11223;
wire n_11570;
wire n_7157;
wire n_2926;
wire n_10937;
wire n_4937;
wire n_8740;
wire n_10493;
wire n_13631;
wire n_5574;
wire n_13264;
wire n_13678;
wire n_8310;
wire n_3391;
wire n_5877;
wire n_14406;
wire n_10104;
wire n_6375;
wire n_11212;
wire n_10552;
wire n_7781;
wire n_13294;
wire n_4786;
wire n_6042;
wire n_8238;
wire n_5203;
wire n_7908;
wire n_10295;
wire n_8296;
wire n_10954;
wire n_7091;
wire n_9788;
wire n_9833;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_9589;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_14590;
wire n_8850;
wire n_9861;
wire n_2855;
wire n_2848;
wire n_7886;
wire n_7675;
wire n_11122;
wire n_6775;
wire n_8943;
wire n_3306;
wire n_4345;
wire n_8993;
wire n_11159;
wire n_12329;
wire n_9205;
wire n_11631;
wire n_9418;
wire n_9946;
wire n_10376;
wire n_7774;
wire n_8634;
wire n_12611;
wire n_11715;
wire n_13625;
wire n_8831;
wire n_6970;
wire n_13034;
wire n_9979;
wire n_12205;
wire n_13122;
wire n_6948;
wire n_3460;
wire n_14324;
wire n_13210;
wire n_5155;
wire n_8676;
wire n_14337;
wire n_11889;
wire n_14509;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_10087;
wire n_5408;
wire n_10341;
wire n_11278;
wire n_12606;
wire n_14692;
wire n_8758;
wire n_11671;
wire n_5812;
wire n_9973;
wire n_5540;
wire n_11782;
wire n_7381;
wire n_5804;
wire n_9007;
wire n_8544;
wire n_3240;
wire n_7999;
wire n_5066;
wire n_14253;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_9020;
wire n_10027;
wire n_9260;
wire n_5130;
wire n_14212;
wire n_4175;
wire n_10154;
wire n_6241;
wire n_13597;
wire n_9619;
wire n_14392;
wire n_13510;
wire n_5200;
wire n_9235;
wire n_3393;
wire n_10161;
wire n_13003;
wire n_8652;
wire n_9112;
wire n_12365;
wire n_2836;
wire n_12423;
wire n_7873;
wire n_12843;
wire n_2864;
wire n_4456;
wire n_11372;
wire n_9691;
wire n_5992;
wire n_8646;
wire n_13573;
wire n_2601;
wire n_12518;
wire n_12861;
wire n_9133;
wire n_5684;
wire n_13708;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_9752;
wire n_6632;
wire n_8999;
wire n_4948;
wire n_3629;
wire n_10902;
wire n_5413;
wire n_7713;
wire n_6623;
wire n_9395;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_6933;
wire n_10294;
wire n_3724;
wire n_9353;
wire n_11155;
wire n_3287;
wire n_11714;
wire n_12293;
wire n_13947;
wire n_3046;
wire n_2921;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_8031;
wire n_3257;
wire n_11590;
wire n_9804;
wire n_12450;
wire n_5737;
wire n_9125;
wire n_8015;
wire n_8412;
wire n_3730;
wire n_8439;
wire n_8575;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_13648;
wire n_5097;
wire n_10323;
wire n_2695;
wire n_7084;
wire n_11976;
wire n_13274;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_4003;
wire n_8499;
wire n_9397;
wire n_10969;
wire n_13015;
wire n_13472;
wire n_13322;
wire n_13870;
wire n_6390;
wire n_7640;
wire n_12000;
wire n_6799;
wire n_8772;
wire n_10806;
wire n_9767;
wire n_12903;
wire n_3014;
wire n_7912;
wire n_6278;
wire n_11430;
wire n_7195;
wire n_12309;
wire n_5640;
wire n_3342;
wire n_13401;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_8557;
wire n_13891;
wire n_3796;
wire n_9384;
wire n_3884;
wire n_4492;
wire n_13850;
wire n_3625;
wire n_13835;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_10666;
wire n_12895;
wire n_5661;
wire n_3760;
wire n_7641;
wire n_4975;
wire n_11638;
wire n_3515;
wire n_12687;
wire n_12023;
wire n_14460;
wire n_5306;
wire n_5905;
wire n_13908;
wire n_8815;
wire n_7949;
wire n_6112;
wire n_11659;
wire n_2728;
wire n_9906;
wire n_8679;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_11948;
wire n_4022;
wire n_7115;
wire n_9310;
wire n_11843;
wire n_10659;
wire n_11689;
wire n_7764;
wire n_8446;
wire n_9163;
wire n_11535;
wire n_12022;
wire n_12624;
wire n_4336;
wire n_11808;
wire n_8789;
wire n_8128;
wire n_7520;
wire n_5314;
wire n_9322;
wire n_12719;
wire n_7616;
wire n_14493;
wire n_10793;
wire n_14491;
wire n_8359;
wire n_5231;
wire n_5064;
wire n_6412;
wire n_6271;
wire n_11108;
wire n_9377;
wire n_7235;
wire n_6572;
wire n_9224;
wire n_10211;
wire n_10837;
wire n_3981;
wire n_14381;
wire n_12664;
wire n_13020;
wire n_11577;
wire n_7271;
wire n_9055;
wire n_13749;
wire n_13311;
wire n_2681;
wire n_7222;
wire n_8678;
wire n_9971;
wire n_8605;
wire n_12981;
wire n_13945;
wire n_3031;
wire n_10976;
wire n_9624;
wire n_6930;
wire n_10045;
wire n_14172;
wire n_10289;
wire n_5482;
wire n_9145;
wire n_12716;
wire n_10232;
wire n_13079;
wire n_11098;
wire n_3215;
wire n_8443;
wire n_8525;
wire n_12166;
wire n_12507;
wire n_3138;
wire n_8312;
wire n_10819;
wire n_2860;
wire n_8901;
wire n_13786;
wire n_13645;
wire n_6584;
wire n_4494;
wire n_9887;
wire n_12044;
wire n_6387;
wire n_9373;
wire n_4201;
wire n_14374;
wire n_6470;
wire n_7206;
wire n_8869;
wire n_11279;
wire n_11729;
wire n_14012;
wire n_9770;
wire n_11514;
wire n_5287;
wire n_8272;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_6625;
wire n_14569;
wire n_4074;
wire n_7383;
wire n_12430;
wire n_3994;
wire n_4636;
wire n_11606;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_10306;
wire n_12902;
wire n_12257;
wire n_11727;
wire n_13299;
wire n_10103;
wire n_14664;
wire n_11337;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_10183;
wire n_12839;
wire n_13693;
wire n_5623;
wire n_11778;
wire n_12925;
wire n_11658;
wire n_10710;
wire n_8870;
wire n_9753;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_10931;
wire n_9468;
wire n_11433;
wire n_8178;
wire n_5524;
wire n_7854;
wire n_9517;
wire n_9544;
wire n_5735;
wire n_7959;
wire n_14338;
wire n_8234;
wire n_6363;
wire n_13434;
wire n_6588;
wire n_11369;
wire n_4243;
wire n_2765;
wire n_7897;
wire n_12759;
wire n_11720;
wire n_14418;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_13500;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_8488;
wire n_11840;
wire n_6865;
wire n_11284;
wire n_12553;
wire n_13113;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_9774;
wire n_7132;
wire n_11987;
wire n_12016;
wire n_12496;
wire n_11052;
wire n_7533;
wire n_9586;
wire n_10670;
wire n_13655;
wire n_10150;
wire n_3377;
wire n_6722;
wire n_9780;
wire n_13476;
wire n_11177;
wire n_6420;
wire n_10004;
wire n_4907;
wire n_11169;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_8862;
wire n_13229;
wire n_14092;
wire n_8184;
wire n_13950;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_11221;
wire n_14219;
wire n_13344;
wire n_10151;
wire n_10353;
wire n_11095;
wire n_10187;
wire n_10171;
wire n_11211;
wire n_7129;
wire n_12138;
wire n_7080;
wire n_4870;
wire n_3374;
wire n_6981;
wire n_7776;
wire n_4818;
wire n_8001;
wire n_10406;
wire n_8695;
wire n_12230;
wire n_12521;
wire n_11236;
wire n_11931;
wire n_7436;
wire n_8767;
wire n_11036;
wire n_12562;
wire n_8571;
wire n_7020;
wire n_11600;
wire n_5935;
wire n_8064;
wire n_14117;
wire n_14588;
wire n_6696;
wire n_13721;
wire n_4916;
wire n_8472;
wire n_13302;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_6045;
wire n_5376;
wire n_12217;
wire n_13535;
wire n_14261;
wire n_3508;
wire n_6300;
wire n_13704;
wire n_6653;
wire n_6372;
wire n_13969;
wire n_4129;
wire n_14016;
wire n_7120;
wire n_11114;
wire n_10479;
wire n_7978;
wire n_10033;
wire n_5488;
wire n_9099;
wire n_6900;
wire n_10034;
wire n_5727;
wire n_11336;
wire n_3599;
wire n_6660;
wire n_8787;
wire n_11009;
wire n_9543;
wire n_8131;
wire n_5988;
wire n_6424;
wire n_10696;
wire n_14633;
wire n_11480;
wire n_5646;
wire n_14538;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_7694;
wire n_8771;
wire n_9245;
wire n_5832;
wire n_13269;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_7142;
wire n_10360;
wire n_6423;
wire n_6526;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_8150;
wire n_9168;
wire n_11423;
wire n_12691;
wire n_5328;
wire n_3819;
wire n_9074;
wire n_12159;
wire n_6011;
wire n_4616;
wire n_5016;
wire n_3222;
wire n_12259;
wire n_11665;
wire n_12975;
wire n_9330;
wire n_9367;
wire n_7465;
wire n_11556;
wire n_11685;
wire n_13402;
wire n_14231;
wire n_5470;
wire n_10230;
wire n_11801;
wire n_12117;
wire n_8917;
wire n_12587;
wire n_11573;
wire n_4374;
wire n_3205;
wire n_6176;
wire n_9300;
wire n_14489;
wire n_13619;
wire n_14663;
wire n_3868;
wire n_11589;
wire n_11667;
wire n_14395;
wire n_8230;
wire n_10414;
wire n_6222;
wire n_13110;
wire n_12422;
wire n_8352;
wire n_7760;
wire n_2593;
wire n_9918;
wire n_12977;
wire n_6969;
wire n_13060;
wire n_2741;
wire n_2714;
wire n_9496;
wire n_13177;
wire n_8914;
wire n_10953;
wire n_14082;
wire n_8821;
wire n_11446;
wire n_13853;
wire n_8465;
wire n_6587;
wire n_6688;
wire n_8360;
wire n_6505;
wire n_13586;
wire n_9837;
wire n_12772;
wire n_5362;
wire n_8209;
wire n_8986;
wire n_14701;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_3611;
wire n_11633;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_11011;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_7629;
wire n_12145;
wire n_10787;
wire n_6987;
wire n_3995;
wire n_7567;
wire n_8743;
wire n_11342;
wire n_8963;
wire n_9191;
wire n_3908;
wire n_11812;
wire n_6453;
wire n_9114;
wire n_6308;
wire n_11142;
wire n_13074;
wire n_10896;
wire n_8396;
wire n_3892;
wire n_13773;
wire n_8514;
wire n_12196;
wire n_13482;
wire n_8550;
wire n_7449;
wire n_11959;
wire n_8151;
wire n_13927;
wire n_14688;
wire n_3501;
wire n_12889;
wire n_13096;
wire n_2555;
wire n_3568;
wire n_3216;
wire n_12493;
wire n_9913;
wire n_2708;
wire n_6187;
wire n_11626;
wire n_6597;
wire n_13810;
wire n_11178;
wire n_12440;
wire n_4844;
wire n_9329;
wire n_6220;
wire n_13684;
wire n_14452;
wire n_12608;
wire n_4049;
wire n_2661;
wire n_10598;
wire n_13008;
wire n_13800;
wire n_7479;
wire n_7882;
wire n_13607;
wire n_11750;
wire n_13742;
wire n_7517;
wire n_9627;
wire n_3551;
wire n_13412;
wire n_11283;
wire n_10271;
wire n_11338;
wire n_5037;
wire n_11295;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_8070;
wire n_4525;
wire n_8866;
wire n_10402;
wire n_6149;
wire n_11191;
wire n_10064;
wire n_3364;
wire n_11661;
wire n_13329;
wire n_10137;
wire n_2643;
wire n_9585;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_9376;
wire n_4369;
wire n_12515;
wire n_3826;
wire n_5648;
wire n_11644;
wire n_12249;
wire n_6439;
wire n_4324;
wire n_11354;
wire n_13537;
wire n_8797;
wire n_14247;
wire n_14462;
wire n_6547;
wire n_13075;
wire n_11126;
wire n_9524;
wire n_7177;
wire n_7902;
wire n_11408;
wire n_12623;
wire n_5160;
wire n_12971;
wire n_2742;
wire n_13051;
wire n_3671;
wire n_12674;
wire n_5762;
wire n_9606;
wire n_14419;
wire n_10800;
wire n_5484;
wire n_12026;
wire n_13038;
wire n_14514;
wire n_13812;
wire n_10019;
wire n_10762;
wire n_14135;
wire n_7353;
wire n_4104;
wire n_11935;
wire n_8054;
wire n_3791;
wire n_10047;
wire n_6478;
wire n_11037;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_13977;
wire n_3199;
wire n_8841;
wire n_11396;
wire n_9084;
wire n_14681;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_14453;
wire n_6906;
wire n_3016;
wire n_6739;
wire n_3367;
wire n_3669;
wire n_10995;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_4528;
wire n_2772;
wire n_14036;
wire n_10597;
wire n_10561;
wire n_7818;
wire n_12345;
wire n_7645;
wire n_5385;
wire n_7482;
wire n_3990;
wire n_13841;
wire n_14312;
wire n_11726;
wire n_12346;
wire n_5622;
wire n_14522;
wire n_14110;
wire n_10523;
wire n_8618;
wire n_10377;
wire n_10243;
wire n_5635;
wire n_4069;
wire n_8538;
wire n_3582;
wire n_8590;
wire n_13883;
wire n_7907;
wire n_9204;
wire n_8970;
wire n_4280;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_8791;
wire n_13724;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_10165;
wire n_9616;
wire n_5380;
wire n_9708;
wire n_7862;
wire n_10153;
wire n_9130;
wire n_9988;
wire n_3735;
wire n_8703;
wire n_12265;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_3656;
wire n_12147;
wire n_7721;
wire n_4524;
wire n_9209;
wire n_8061;
wire n_2831;
wire n_10775;
wire n_10173;
wire n_10585;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_12075;
wire n_8754;
wire n_8864;
wire n_5941;
wire n_10985;
wire n_4891;
wire n_11300;
wire n_14294;
wire n_8837;
wire n_12108;
wire n_10999;
wire n_13425;
wire n_2629;
wire n_3369;
wire n_13791;
wire n_8915;
wire n_10587;
wire n_8784;
wire n_11219;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_11857;
wire n_5597;
wire n_11735;
wire n_11986;
wire n_9086;
wire n_8768;
wire n_12102;
wire n_6999;
wire n_8072;
wire n_8086;
wire n_9014;
wire n_5469;
wire n_6019;
wire n_3685;
wire n_7539;
wire n_14611;
wire n_9010;
wire n_11637;
wire n_13925;
wire n_6440;
wire n_4977;
wire n_8774;
wire n_14417;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_11072;
wire n_12183;
wire n_2939;
wire n_3425;
wire n_13432;
wire n_4876;
wire n_5021;
wire n_12519;
wire n_2900;
wire n_12955;
wire n_9044;
wire n_2912;
wire n_13538;
wire n_14176;
wire n_5936;
wire n_14650;
wire n_8307;
wire n_3813;
wire n_13774;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_9694;
wire n_11421;
wire n_13323;
wire n_10718;
wire n_13214;
wire n_10951;
wire n_10412;
wire n_8470;
wire n_5928;
wire n_7830;
wire n_8050;
wire n_3124;
wire n_3811;
wire n_10310;
wire n_4200;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_10655;
wire n_9633;
wire n_6165;
wire n_10133;
wire n_12793;
wire n_3463;
wire n_11989;
wire n_10942;
wire n_2785;
wire n_4938;
wire n_2574;
wire n_6114;
wire n_13192;
wire n_2928;
wire n_13392;
wire n_5505;
wire n_13433;
wire n_12865;
wire n_14662;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_9261;
wire n_11331;
wire n_12285;
wire n_5504;
wire n_7348;
wire n_9345;
wire n_11953;
wire n_4118;
wire n_6829;
wire n_11820;
wire n_12478;
wire n_3857;
wire n_3110;
wire n_9375;
wire n_4239;
wire n_9472;
wire n_9764;
wire n_10509;
wire n_8010;
wire n_3157;
wire n_13059;
wire n_12522;
wire n_13451;
wire n_2730;
wire n_9448;
wire n_6464;
wire n_8802;
wire n_8950;
wire n_5129;
wire n_13199;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_8603;
wire n_9487;
wire n_10639;
wire n_13588;
wire n_5494;
wire n_5970;
wire n_11358;
wire n_12413;
wire n_6838;
wire n_13191;
wire n_2700;
wire n_6368;
wire n_14133;
wire n_10690;
wire n_12369;
wire n_12681;
wire n_7935;
wire n_11118;
wire n_8143;
wire n_11844;
wire n_9271;
wire n_3640;
wire n_5663;
wire n_12084;
wire n_5161;
wire n_14132;
wire n_7933;
wire n_12152;
wire n_12726;
wire n_12784;
wire n_7155;
wire n_6640;
wire n_9851;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_6850;
wire n_4343;
wire n_3879;
wire n_12520;
wire n_12511;
wire n_4764;
wire n_7743;
wire n_5389;
wire n_11861;
wire n_12705;
wire n_13899;
wire n_4990;
wire n_2986;
wire n_8584;
wire n_14443;
wire n_11370;
wire n_13017;
wire n_9101;
wire n_6550;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_3591;
wire n_8574;
wire n_12832;
wire n_2760;
wire n_4919;
wire n_13422;
wire n_7043;
wire n_7986;
wire n_3317;
wire n_8049;
wire n_9927;
wire n_12207;
wire n_13666;
wire n_12782;
wire n_7266;
wire n_13042;
wire n_10621;
wire n_11884;
wire n_5653;
wire n_4835;
wire n_4420;
wire n_7996;
wire n_14513;
wire n_12970;
wire n_10789;
wire n_4251;
wire n_5266;
wire n_10496;
wire n_12384;
wire n_4559;
wire n_4742;
wire n_12605;
wire n_5038;
wire n_3566;
wire n_10319;
wire n_5800;
wire n_14021;
wire n_8509;
wire n_12408;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_9850;
wire n_4162;
wire n_5766;
wire n_10499;
wire n_14223;
wire n_11717;
wire n_5293;
wire n_10224;
wire n_13234;
wire n_4790;
wire n_7035;
wire n_10970;
wire n_4173;
wire n_8354;
wire n_12651;
wire n_5309;
wire n_6047;
wire n_9432;
wire n_3573;
wire n_2943;
wire n_12160;
wire n_13829;
wire n_11464;
wire n_3319;
wire n_11243;
wire n_9824;
wire n_14582;
wire n_8277;
wire n_7442;
wire n_4727;
wire n_10827;
wire n_6568;
wire n_3654;
wire n_11473;
wire n_14508;
wire n_5627;
wire n_3783;
wire n_10055;
wire n_12638;
wire n_12698;
wire n_4008;
wire n_11654;
wire n_13878;
wire n_10783;
wire n_14562;
wire n_8583;
wire n_3643;
wire n_3184;
wire n_7153;
wire n_8681;
wire n_6258;
wire n_8644;
wire n_10148;
wire n_7939;
wire n_9884;
wire n_7715;
wire n_11534;
wire n_3982;
wire n_10465;
wire n_14040;
wire n_14361;
wire n_11749;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_10610;
wire n_8609;
wire n_13955;
wire n_9144;
wire n_3973;
wire n_8052;
wire n_12481;
wire n_4799;
wire n_8733;
wire n_9758;
wire n_12078;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_12815;
wire n_4534;
wire n_12129;
wire n_5636;
wire n_4960;
wire n_9931;
wire n_7699;
wire n_9693;
wire n_11546;
wire n_12502;
wire n_10830;
wire n_9273;
wire n_9196;
wire n_5707;
wire n_5594;
wire n_9029;
wire n_10086;
wire n_3738;
wire n_5697;
wire n_13763;
wire n_7580;
wire n_5606;
wire n_11785;
wire n_6727;
wire n_5911;
wire n_12697;
wire n_7340;
wire n_8080;
wire n_13437;
wire n_3600;
wire n_10279;
wire n_7303;
wire n_10932;
wire n_11440;
wire n_9967;
wire n_12908;
wire n_8819;
wire n_7870;
wire n_6139;
wire n_7568;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_8487;
wire n_13293;
wire n_3027;
wire n_6454;
wire n_11545;
wire n_4011;
wire n_11697;
wire n_3695;
wire n_13487;
wire n_3800;
wire n_13555;
wire n_13239;
wire n_3462;
wire n_10487;
wire n_14579;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_9881;
wire n_2820;
wire n_3733;
wire n_11645;
wire n_3967;
wire n_12512;
wire n_11263;
wire n_12199;
wire n_6333;
wire n_11937;
wire n_7004;
wire n_12584;
wire n_13854;
wire n_13361;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_10910;
wire n_5058;
wire n_8382;
wire n_9733;
wire n_3096;
wire n_8517;
wire n_7207;
wire n_8827;
wire n_13558;
wire n_9075;
wire n_11324;
wire n_13954;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_11763;
wire n_13803;
wire n_7167;
wire n_5849;
wire n_3233;
wire n_11853;
wire n_3322;
wire n_12988;
wire n_14537;
wire n_8906;
wire n_5841;
wire n_10109;
wire n_7146;
wire n_7030;
wire n_14542;
wire n_10857;
wire n_4478;
wire n_8203;
wire n_2935;
wire n_9442;
wire n_4246;
wire n_7618;
wire n_14625;
wire n_2863;
wire n_13244;
wire n_4632;
wire n_13305;
wire n_12284;
wire n_11364;
wire n_11941;
wire n_9630;
wire n_4061;
wire n_11359;
wire n_12031;
wire n_14203;
wire n_9898;
wire n_11323;
wire n_11504;
wire n_11704;
wire n_2920;
wire n_11587;
wire n_11620;
wire n_13697;
wire n_3344;
wire n_8340;
wire n_4754;
wire n_12652;
wire n_9582;
wire n_8268;
wire n_10865;
wire n_8171;
wire n_4375;
wire n_12850;
wire n_9877;
wire n_14578;
wire n_10179;
wire n_12969;
wire n_10925;
wire n_12607;
wire n_12379;
wire n_3368;
wire n_9986;
wire n_13743;
wire n_13951;
wire n_14222;
wire n_13695;
wire n_8008;
wire n_7633;
wire n_10246;
wire n_9636;
wire n_3117;
wire n_4684;
wire n_10439;
wire n_13376;
wire n_14377;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_8553;
wire n_2592;
wire n_8824;
wire n_11902;
wire n_3490;
wire n_7280;
wire n_8369;
wire n_5043;
wire n_12701;
wire n_14008;
wire n_7339;
wire n_7597;
wire n_8884;
wire n_12898;
wire n_4241;
wire n_2751;
wire n_3113;
wire n_9225;
wire n_4183;
wire n_7768;
wire n_11282;
wire n_5645;
wire n_6455;
wire n_5020;
wire n_13639;
wire n_2842;
wire n_7615;
wire n_12475;
wire n_3603;
wire n_10182;
wire n_8271;
wire n_9091;
wire n_3720;
wire n_6183;
wire n_13772;
wire n_14643;
wire n_12027;
wire n_8392;
wire n_8309;
wire n_6107;
wire n_12218;
wire n_10795;
wire n_13602;
wire n_6476;
wire n_5232;
wire n_10046;
wire n_2560;
wire n_4256;
wire n_9412;
wire n_11834;
wire n_8874;
wire n_8228;
wire n_12174;
wire n_5035;
wire n_11405;
wire n_11028;
wire n_3037;
wire n_11663;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_8483;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_12385;
wire n_14407;
wire n_3363;
wire n_6636;
wire n_9525;
wire n_11071;
wire n_12289;
wire n_11625;
wire n_11187;
wire n_12041;
wire n_12565;
wire n_3522;
wire n_12882;
wire n_13736;
wire n_13254;
wire n_12819;
wire n_8172;
wire n_4455;
wire n_13341;
wire n_3241;
wire n_6554;
wire n_3899;
wire n_9575;
wire n_5631;
wire n_3481;
wire n_6994;
wire n_7401;
wire n_10413;
wire n_10456;
wire n_11566;
wire n_11271;
wire n_12164;
wire n_12433;
wire n_11649;
wire n_12224;
wire n_13061;
wire n_5101;
wire n_9738;
wire n_10735;
wire n_6020;
wire n_13328;
wire n_9252;
wire n_12550;
wire n_6185;
wire n_8344;
wire n_12800;
wire n_14568;
wire n_14259;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_12561;
wire n_8738;
wire n_8936;
wire n_10822;
wire n_9739;
wire n_6785;
wire n_2803;
wire n_9727;
wire n_2887;
wire n_10508;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_13281;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_8226;
wire n_6695;
wire n_7529;
wire n_5608;
wire n_3354;
wire n_6501;
wire n_11308;
wire n_11739;
wire n_11593;
wire n_9148;
wire n_10858;
wire n_6466;
wire n_10736;
wire n_11828;
wire n_9958;
wire n_3437;
wire n_6467;
wire n_9323;
wire n_14138;
wire n_4212;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_9779;
wire n_8088;
wire n_5702;
wire n_14244;
wire n_9545;
wire n_8930;
wire n_9155;
wire n_12563;
wire n_8662;
wire n_13114;
wire n_11291;
wire n_3574;
wire n_11425;
wire n_13566;
wire n_9046;
wire n_9430;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_9625;
wire n_11890;
wire n_13621;
wire n_8783;
wire n_12398;
wire n_13624;
wire n_5182;
wire n_4217;
wire n_8663;
wire n_14015;
wire n_10928;
wire n_5277;
wire n_6507;
wire n_10842;
wire n_12941;
wire n_6618;
wire n_9447;
wire n_13407;
wire n_2951;
wire n_4048;
wire n_3807;
wire n_13404;
wire n_6213;
wire n_8364;
wire n_9485;
wire n_4949;
wire n_2974;
wire n_8490;
wire n_8981;
wire n_9129;
wire n_12461;
wire n_11832;
wire n_7872;
wire n_6873;
wire n_3969;
wire n_7958;
wire n_4605;
wire n_8118;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_8671;
wire n_7101;
wire n_12095;
wire n_14191;
wire n_8785;
wire n_11294;
wire n_11744;
wire n_10210;
wire n_11470;
wire n_13994;
wire n_7843;
wire n_12998;
wire n_9047;
wire n_13219;
wire n_10057;
wire n_6063;
wire n_13737;
wire n_2858;
wire n_12630;
wire n_11641;
wire n_3076;
wire n_7578;
wire n_12789;
wire n_12679;
wire n_14146;
wire n_3410;
wire n_13372;
wire n_5415;
wire n_14084;
wire n_7261;
wire n_8982;
wire n_10739;
wire n_4592;
wire n_4999;
wire n_12327;
wire n_6993;
wire n_9745;
wire n_14288;
wire n_12038;
wire n_13932;
wire n_10533;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_13978;
wire n_11875;
wire n_8100;
wire n_10878;
wire n_2589;
wire n_4086;
wire n_10988;
wire n_8522;
wire n_13563;
wire n_13141;
wire n_12338;
wire n_10993;
wire n_13249;
wire n_8381;
wire n_9320;
wire n_8835;
wire n_6767;
wire n_11014;
wire n_4656;
wire n_4862;
wire n_12030;
wire n_14553;
wire n_5687;
wire n_6558;
wire n_13517;
wire n_6755;
wire n_9108;
wire n_9457;
wire n_9907;
wire n_10959;
wire n_6153;
wire n_11310;
wire n_3536;
wire n_7263;
wire n_11062;
wire n_3782;
wire n_10940;
wire n_12067;
wire n_13783;
wire n_12675;
wire n_6608;
wire n_11400;
wire n_11040;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_13968;
wire n_12870;
wire n_14038;
wire n_3594;
wire n_12291;
wire n_5383;
wire n_6635;
wire n_7245;
wire n_7925;
wire n_7310;
wire n_9567;
wire n_6359;
wire n_11773;
wire n_14385;
wire n_5690;
wire n_10583;
wire n_14027;
wire n_11332;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_7585;
wire n_8356;
wire n_13279;
wire n_5029;
wire n_13731;
wire n_12013;
wire n_13007;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_9852;
wire n_10881;
wire n_12395;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_14049;
wire n_13160;
wire n_2985;
wire n_11943;
wire n_5218;
wire n_10544;
wire n_12933;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_13895;
wire n_14403;
wire n_13213;
wire n_8736;
wire n_3114;
wire n_10491;
wire n_12131;
wire n_13507;
wire n_6082;
wire n_11144;
wire n_13385;
wire n_10926;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_11841;
wire n_8918;
wire n_11766;
wire n_12766;
wire n_10839;
wire n_3047;
wire n_10603;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_9022;
wire n_13790;
wire n_7514;
wire n_12399;
wire n_8616;
wire n_6105;
wire n_12762;
wire n_10400;
wire n_11518;
wire n_5512;
wire n_13567;
wire n_7738;
wire n_14346;
wire n_2808;
wire n_8838;
wire n_8908;
wire n_13687;
wire n_3520;
wire n_11960;
wire n_7609;
wire n_13580;
wire n_9161;
wire n_3272;
wire n_12241;
wire n_10792;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_11274;
wire n_6548;
wire n_8607;
wire n_13779;
wire n_8213;
wire n_14487;
wire n_13722;
wire n_13225;
wire n_14615;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_10994;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_13514;
wire n_13806;
wire n_2676;
wire n_9903;
wire n_9831;
wire n_14595;
wire n_10032;
wire n_8436;
wire n_7282;
wire n_13261;
wire n_8551;
wire n_14638;
wire n_13039;
wire n_2770;
wire n_4550;
wire n_9238;
wire n_12137;
wire n_14167;
wire n_4347;
wire n_11624;
wire n_10580;
wire n_7921;
wire n_5193;
wire n_4933;
wire n_4144;
wire n_10512;
wire n_9248;
wire n_12495;
wire n_5514;
wire n_11917;
wire n_5611;
wire n_3278;
wire n_12790;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_9867;
wire n_12106;
wire n_11130;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_10005;
wire n_11053;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_11872;
wire n_12434;
wire n_5188;
wire n_6674;
wire n_13669;
wire n_5049;
wire n_12710;
wire n_7489;
wire n_9056;
wire n_6331;
wire n_5308;
wire n_9106;
wire n_4434;
wire n_13303;
wire n_5068;
wire n_12881;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_14496;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_10596;
wire n_12920;
wire n_4019;
wire n_4199;
wire n_14260;
wire n_7968;
wire n_11220;
wire n_10061;
wire n_10507;
wire n_6023;
wire n_7820;
wire n_8437;
wire n_7833;
wire n_12086;
wire n_11887;
wire n_3829;
wire n_14189;
wire n_12281;
wire n_12991;
wire n_4510;
wire n_14552;
wire n_7750;
wire n_5057;
wire n_9071;
wire n_6196;
wire n_12995;
wire n_5425;
wire n_5273;
wire n_10136;
wire n_5839;
wire n_7588;
wire n_10967;
wire n_11551;
wire n_14339;
wire n_13368;
wire n_10369;
wire n_3546;
wire n_7697;
wire n_10025;
wire n_10708;
wire n_11703;
wire n_5887;
wire n_13948;
wire n_7808;
wire n_3068;
wire n_9519;
wire n_9027;
wire n_7603;
wire n_13598;
wire n_6321;
wire n_14180;
wire n_5683;
wire n_8704;
wire n_14341;
wire n_3002;
wire n_8984;
wire n_9786;
wire n_10194;
wire n_7192;
wire n_12807;
wire n_5248;
wire n_4899;
wire n_11153;
wire n_10833;
wire n_3146;
wire n_10685;
wire n_3038;
wire n_10513;
wire n_4156;
wire n_8613;
wire n_13611;
wire n_11030;
wire n_14704;
wire n_3693;
wire n_13178;
wire n_14293;
wire n_10223;
wire n_5880;
wire n_13495;
wire n_8012;
wire n_12012;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_8881;
wire n_5531;
wire n_9404;
wire n_13777;
wire n_3681;
wire n_5666;
wire n_13301;
wire n_3970;
wire n_11368;
wire n_12098;
wire n_7988;
wire n_12025;
wire n_12669;
wire n_13205;
wire n_3188;
wire n_4448;
wire n_10410;
wire n_13049;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_8763;
wire n_6450;
wire n_9370;
wire n_6995;
wire n_13009;
wire n_4193;
wire n_4579;
wire n_6347;
wire n_13748;
wire n_13338;
wire n_6496;
wire n_13747;
wire n_4776;
wire n_8387;
wire n_9352;
wire n_11716;
wire n_14083;
wire n_8105;
wire n_10984;
wire n_13485;
wire n_10144;
wire n_12019;
wire n_2704;
wire n_6745;
wire n_7943;
wire n_6698;
wire n_3729;
wire n_4471;
wire n_6968;
wire n_13416;
wire n_11967;
wire n_7377;
wire n_12255;
wire n_8900;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_9681;
wire n_14439;
wire n_8353;
wire n_12503;
wire n_9051;
wire n_7723;
wire n_3028;
wire n_4691;
wire n_7904;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_5461;
wire n_9098;
wire n_12415;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_8323;
wire n_13053;
wire n_13752;
wire n_10459;
wire n_12951;
wire n_14125;
wire n_6164;
wire n_11426;
wire n_8711;
wire n_13273;
wire n_3616;
wire n_11628;
wire n_4753;
wire n_12704;
wire n_9484;
wire n_4803;
wire n_8731;
wire n_3874;
wire n_5730;
wire n_10155;
wire n_11367;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_5754;
wire n_11418;
wire n_2852;
wire n_8597;
wire n_6330;
wire n_7178;
wire n_11026;
wire n_7045;
wire n_11576;
wire n_3637;
wire n_9853;
wire n_8534;
wire n_8655;
wire n_9210;
wire n_12884;
wire n_13324;
wire n_4893;
wire n_10915;
wire n_13414;
wire n_13894;
wire n_10949;
wire n_7777;
wire n_12339;
wire n_8302;
wire n_14616;
wire n_4258;
wire n_5756;
wire n_14695;
wire n_14455;
wire n_12911;
wire n_8496;
wire n_7693;
wire n_11150;
wire n_2917;
wire n_3194;
wire n_10156;
wire n_5033;
wire n_11123;
wire n_14414;
wire n_10248;
wire n_6015;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_14449;
wire n_11733;
wire n_3461;
wire n_10215;
wire n_10624;
wire n_12915;
wire n_7682;
wire n_7300;
wire n_6861;
wire n_10152;
wire n_12888;
wire n_4203;
wire n_12105;
wire n_9756;
wire n_5789;
wire n_12034;
wire n_5400;
wire n_7558;
wire n_5347;
wire n_2957;
wire n_11188;
wire n_9166;
wire n_8103;
wire n_8719;
wire n_10877;
wire n_7798;
wire n_9778;
wire n_8879;
wire n_13906;
wire n_4767;
wire n_8969;
wire n_9141;
wire n_4569;
wire n_11209;
wire n_6528;
wire n_14441;
wire n_13159;
wire n_9700;
wire n_10316;
wire n_8896;
wire n_5144;
wire n_3820;
wire n_11503;
wire n_6895;
wire n_3072;
wire n_10385;
wire n_8335;
wire n_2961;
wire n_13337;
wire n_4468;
wire n_5509;
wire n_3848;
wire n_7400;
wire n_14230;
wire n_11699;
wire n_13145;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_12549;
wire n_6523;
wire n_11817;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_14618;
wire n_11469;
wire n_9363;
wire n_11971;
wire n_4698;
wire n_14199;
wire n_3674;
wire n_5349;
wire n_14101;
wire n_6472;
wire n_3763;
wire n_9532;
wire n_10823;
wire n_12237;
wire n_14001;
wire n_6389;
wire n_14586;
wire n_3499;
wire n_14623;
wire n_14635;
wire n_10680;
wire n_5534;
wire n_9307;
wire n_13922;
wire n_9876;
wire n_12220;
wire n_3910;
wire n_3947;
wire n_12564;
wire n_10814;
wire n_12375;
wire n_13333;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_6073;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_8462;
wire n_9959;
wire n_3228;
wire n_8834;
wire n_9989;
wire n_10651;
wire n_14495;
wire n_8286;
wire n_8417;
wire n_13872;
wire n_12809;
wire n_2678;
wire n_8964;
wire n_10611;
wire n_6869;
wire n_4761;
wire n_4627;
wire n_10549;
wire n_10370;
wire n_11621;
wire n_7672;
wire n_10770;
wire n_14171;
wire n_4556;
wire n_6137;
wire n_9467;
wire n_11558;
wire n_12043;
wire n_3088;
wire n_12513;
wire n_5254;
wire n_3590;
wire n_12337;
wire n_10393;
wire n_5079;
wire n_8247;
wire n_2761;
wire n_9406;
wire n_10089;
wire n_11417;
wire n_11113;
wire n_14182;
wire n_4520;
wire n_10543;
wire n_13355;
wire n_8639;
wire n_12504;
wire n_11301;
wire n_9160;
wire n_3295;
wire n_5751;
wire n_11051;
wire n_12489;
wire n_10321;
wire n_12886;
wire n_13308;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_6885;
wire n_7681;
wire n_5039;
wire n_6613;
wire n_6580;
wire n_8727;
wire n_8566;
wire n_4265;
wire n_8482;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_13923;
wire n_11018;
wire n_13905;
wire n_10259;
wire n_7491;
wire n_12836;
wire n_14243;
wire n_13936;
wire n_10909;
wire n_10094;
wire n_8599;
wire n_4612;
wire n_14386;
wire n_5997;
wire n_10302;
wire n_11328;
wire n_8781;
wire n_5375;
wire n_5438;
wire n_9167;
wire n_11276;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_6602;
wire n_6530;
wire n_7915;
wire n_4149;
wire n_4958;
wire n_6135;
wire n_12655;
wire n_10623;
wire n_8839;
wire n_11326;
wire n_13627;
wire n_14359;
wire n_5563;
wire n_3030;
wire n_4538;
wire n_3505;
wire n_3075;
wire n_13882;
wire n_12779;
wire n_8365;
wire n_13144;
wire n_14085;
wire n_6942;
wire n_7860;
wire n_14108;
wire n_6892;
wire n_4730;
wire n_7357;
wire n_8112;
wire n_8489;
wire n_13364;
wire n_8859;
wire n_8060;
wire n_9290;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_3697;
wire n_8244;
wire n_13134;
wire n_13340;
wire n_6977;
wire n_7229;
wire n_12688;
wire n_11732;
wire n_10485;
wire n_8096;
wire n_11946;
wire n_7336;
wire n_5932;
wire n_11334;
wire n_6598;
wire n_10105;
wire n_6795;
wire n_6121;
wire n_11855;
wire n_12321;
wire n_3430;
wire n_5919;
wire n_8346;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_11781;
wire n_13310;
wire n_14548;
wire n_14306;
wire n_11080;
wire n_9705;
wire n_4967;
wire n_8367;
wire n_4696;
wire n_9113;
wire n_10761;
wire n_12104;
wire n_14074;
wire n_3484;
wire n_6001;
wire n_13445;
wire n_14043;
wire n_4971;
wire n_9521;
wire n_9682;
wire n_14676;
wire n_7493;
wire n_9278;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_14355;
wire n_2590;
wire n_4661;
wire n_3041;
wire n_2797;
wire n_5823;
wire n_8898;
wire n_8658;
wire n_9222;
wire n_5944;
wire n_8905;
wire n_5422;
wire n_6989;
wire n_8145;
wire n_8237;
wire n_6299;
wire n_11445;
wire n_12643;
wire n_10592;
wire n_9813;
wire n_7424;
wire n_10216;
wire n_5246;
wire n_8562;
wire n_4376;
wire n_9863;
wire n_3832;
wire n_10616;
wire n_11350;
wire n_14527;
wire n_12799;
wire n_3525;
wire n_13833;
wire n_3712;
wire n_12202;
wire n_12694;
wire n_11057;
wire n_9394;
wire n_10170;
wire n_11182;
wire n_4305;
wire n_11140;
wire n_2953;
wire n_2823;
wire n_11082;
wire n_7273;
wire n_9663;
wire n_7901;
wire n_3684;
wire n_14371;
wire n_5725;
wire n_10146;
wire n_5404;
wire n_10175;
wire n_11949;
wire n_13576;
wire n_12055;
wire n_4834;
wire n_9994;
wire n_5332;
wire n_7149;
wire n_9723;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_4692;
wire n_11693;
wire n_12506;
wire n_8211;
wire n_3268;
wire n_2559;
wire n_8537;
wire n_8946;
wire n_5616;
wire n_8055;
wire n_10848;
wire n_4259;
wire n_5870;
wire n_7909;
wire n_12788;
wire n_12894;
wire n_6053;
wire n_11024;
wire n_6233;
wire n_10450;
wire n_10918;
wire n_12333;
wire n_13502;
wire n_4299;
wire n_13131;
wire n_5625;
wire n_13238;
wire n_14597;
wire n_6758;
wire n_5367;
wire n_9069;
wire n_12866;
wire n_6629;
wire n_5288;
wire n_13247;
wire n_11158;
wire n_2694;
wire n_6356;
wire n_8332;
wire n_5601;
wire n_4965;
wire n_3742;
wire n_7601;
wire n_8998;
wire n_13391;
wire n_14190;
wire n_11046;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_11390;
wire n_12551;
wire n_11224;
wire n_13970;
wire n_10536;
wire n_14696;
wire n_8157;
wire n_9284;
wire n_4953;
wire n_10990;
wire n_8484;
wire n_4813;
wire n_3352;
wire n_12223;
wire n_12627;
wire n_12390;
wire n_7147;
wire n_7596;
wire n_9556;
wire n_12226;
wire n_14546;
wire n_5294;
wire n_11380;
wire n_8161;
wire n_5570;
wire n_11101;
wire n_6411;
wire n_11578;
wire n_9337;
wire n_2731;
wire n_5411;
wire n_5670;
wire n_3703;
wire n_13256;
wire n_11015;
wire n_11214;
wire n_9211;
wire n_12378;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_10278;
wire n_4802;
wire n_4793;
wire n_10482;
wire n_14174;
wire n_6032;
wire n_10996;
wire n_5733;
wire n_8692;
wire n_3435;
wire n_12794;
wire n_4897;
wire n_9243;
wire n_14046;
wire n_12436;
wire n_6918;
wire n_10733;
wire n_9773;
wire n_14158;
wire n_4674;
wire n_8812;
wire n_14218;
wire n_11033;
wire n_8682;
wire n_13170;
wire n_4796;
wire n_8290;
wire n_7138;
wire n_13664;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_7976;
wire n_9928;
wire n_10975;
wire n_2750;
wire n_11950;
wire n_8890;
wire n_10484;
wire n_12962;
wire n_8747;
wire n_7617;
wire n_12094;
wire n_4575;
wire n_9784;
wire n_10641;
wire n_11115;
wire n_12964;
wire n_3665;
wire n_3063;
wire n_8062;
wire n_14120;
wire n_3281;
wire n_7137;
wire n_5061;
wire n_3535;
wire n_14652;
wire n_14412;
wire n_3858;
wire n_14499;
wire n_4653;
wire n_7700;
wire n_11709;
wire n_8275;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_10584;
wire n_14609;
wire n_8667;
wire n_4581;
wire n_3220;
wire n_9192;
wire n_10365;
wire n_14427;
wire n_6008;
wire n_10778;
wire n_4625;
wire n_11607;
wire n_11542;
wire n_7098;
wire n_6181;
wire n_14668;
wire n_5070;
wire n_4845;
wire n_13105;
wire n_4148;
wire n_9134;
wire n_12838;
wire n_13964;
wire n_3679;
wire n_5575;
wire n_6654;
wire n_11491;
wire n_7661;
wire n_4968;
wire n_7801;
wire n_8807;
wire n_9975;
wire n_13766;
wire n_9765;
wire n_11896;
wire n_13525;
wire n_6907;
wire n_4590;
wire n_5177;
wire n_4038;
wire n_3856;
wire n_11371;
wire n_11939;
wire n_5316;
wire n_7876;
wire n_2735;
wire n_14332;
wire n_4214;
wire n_13081;
wire n_10378;
wire n_5290;
wire n_13057;
wire n_10324;
wire n_11563;
wire n_2709;
wire n_3419;
wire n_7323;
wire n_13861;
wire n_10850;
wire n_5048;
wire n_11565;
wire n_13129;
wire n_13257;
wire n_5363;
wire n_14583;
wire n_11164;
wire n_12633;
wire n_5665;
wire n_6517;
wire n_11401;
wire n_11414;
wire n_4892;
wire n_6339;
wire n_10330;
wire n_12514;
wire n_14408;
wire n_14659;
wire n_9564;
wire n_14267;
wire n_9127;
wire n_11199;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_14370;
wire n_5607;
wire n_7929;
wire n_14516;
wire n_2782;
wire n_3929;
wire n_11319;
wire n_9306;
wire n_4353;
wire n_8212;
wire n_4950;
wire n_10442;
wire n_7755;
wire n_6504;
wire n_9891;
wire n_13865;
wire n_13135;
wire n_10962;
wire n_10022;
wire n_13973;
wire n_4176;
wire n_9078;
wire n_7556;
wire n_11415;
wire n_13553;
wire n_4124;
wire n_4431;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_10972;
wire n_6814;
wire n_7216;
wire n_13248;
wire n_4488;
wire n_10127;
wire n_5278;
wire n_14278;
wire n_2779;
wire n_3627;
wire n_10824;
wire n_3596;
wire n_5214;
wire n_11128;
wire n_9332;
wire n_12262;
wire n_3756;
wire n_12391;
wire n_8223;
wire n_8043;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_8159;
wire n_5845;
wire n_8868;
wire n_9889;
wire n_4608;
wire n_9294;
wire n_12731;
wire n_6691;
wire n_13623;
wire n_13775;
wire n_12235;
wire n_3948;
wire n_4839;
wire n_9174;
wire n_5969;
wire n_10375;
wire n_9132;
wire n_13464;
wire n_2650;
wire n_4454;
wire n_11669;
wire n_4184;
wire n_9547;
wire n_6343;
wire n_12406;
wire n_6005;
wire n_3883;
wire n_6686;
wire n_4032;
wire n_12929;
wire n_2571;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_14067;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_6025;
wire n_12229;
wire n_3049;
wire n_8434;
wire n_14264;
wire n_3634;
wire n_12508;
wire n_5436;
wire n_7962;
wire n_6697;
wire n_11262;
wire n_12271;
wire n_3066;
wire n_11110;
wire n_12803;
wire n_13084;
wire n_14451;
wire n_14614;
wire n_10122;
wire n_6085;
wire n_10898;
wire n_3913;
wire n_9762;
wire n_11849;
wire n_5341;
wire n_8608;
wire n_2575;
wire n_13583;
wire n_3739;
wire n_5140;
wire n_13470;
wire n_12245;
wire n_2942;
wire n_6062;
wire n_4541;
wire n_14394;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_8656;
wire n_3861;
wire n_5096;
wire n_9183;
wire n_11287;
wire n_6771;
wire n_7905;
wire n_4171;
wire n_11247;
wire n_5847;
wire n_7204;
wire n_12376;
wire n_9461;
wire n_9117;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_12773;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_10116;
wire n_10590;
wire n_10991;
wire n_11945;
wire n_11769;
wire n_4884;
wire n_3580;
wire n_12720;
wire n_12736;
wire n_8249;
wire n_4276;
wire n_5268;
wire n_5050;
wire n_9062;
wire n_5240;
wire n_5503;
wire n_5718;
wire n_7208;
wire n_9915;
wire n_7718;
wire n_10265;
wire n_13006;
wire n_11277;
wire n_12459;
wire n_11075;
wire n_5001;
wire n_12708;
wire n_6567;
wire n_11919;
wire n_12387;
wire n_13705;
wire n_5658;
wire n_4174;
wire n_9001;
wire n_13599;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_13077;
wire n_9081;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_9156;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_8717;
wire n_10159;
wire n_5174;
wire n_9024;
wire n_9198;
wire n_10178;
wire n_4801;
wire n_10571;
wire n_6079;
wire n_6260;
wire n_4582;
wire n_14268;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_13892;
wire n_14251;
wire n_12239;
wire n_14136;
wire n_12636;
wire n_14002;
wire n_3119;
wire n_6671;
wire n_11085;
wire n_9335;
wire n_4740;
wire n_10550;
wire n_9488;
wire n_7632;
wire n_4394;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_11510;
wire n_9725;
wire n_8842;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_10185;
wire n_12648;
wire n_9526;
wire n_4920;
wire n_3909;
wire n_10809;
wire n_13316;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_13140;
wire n_5541;
wire n_6314;
wire n_10660;
wire n_13162;
wire n_12501;
wire n_5610;
wire n_9962;
wire n_8576;
wire n_2810;
wire n_12755;
wire n_6703;
wire n_14262;
wire n_10657;
wire n_10627;
wire n_8799;
wire n_4378;
wire n_9667;
wire n_5166;
wire n_2683;
wire n_11256;
wire n_6065;
wire n_7265;
wire n_12441;
wire n_14018;
wire n_4180;
wire n_11516;
wire n_11520;
wire n_4459;
wire n_6878;
wire n_11461;
wire n_11137;
wire n_3624;
wire n_6725;
wire n_8181;
wire n_5808;
wire n_6527;
wire n_4594;
wire n_13604;
wire n_8447;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_14029;
wire n_13157;
wire n_2748;
wire n_11536;
wire n_11544;
wire n_14488;
wire n_10897;
wire n_4642;
wire n_13952;
wire n_14234;
wire n_9716;
wire n_6913;
wire n_7473;
wire n_7242;
wire n_9253;
wire n_6533;
wire n_11305;
wire n_14126;
wire n_7164;
wire n_2925;
wire n_8022;
wire n_10617;
wire n_12011;
wire n_3544;
wire n_6845;
wire n_10451;
wire n_5300;
wire n_8227;
wire n_14438;
wire n_10768;
wire n_7853;
wire n_3852;
wire n_11268;
wire n_13707;
wire n_5233;
wire n_12742;
wire n_10309;
wire n_5381;
wire n_9796;
wire n_5770;
wire n_7483;
wire n_13868;
wire n_8756;
wire n_5710;
wire n_10021;
wire n_9953;
wire n_2628;
wire n_7389;
wire n_10053;
wire n_3219;
wire n_10315;
wire n_5333;
wire n_5799;
wire n_10765;
wire n_6265;
wire n_4914;
wire n_12317;
wire n_8604;
wire n_12831;
wire n_8809;
wire n_13092;
wire n_8976;
wire n_11815;
wire n_13694;
wire n_3510;
wire n_10907;
wire n_7046;
wire n_13928;
wire n_7834;
wire n_10312;
wire n_11299;
wire n_4587;
wire n_3688;
wire n_11273;
wire n_8940;
wire n_5008;
wire n_9077;
wire n_12872;
wire n_13147;
wire n_12871;
wire n_3871;
wire n_13212;
wire n_12590;
wire n_14503;
wire n_14325;
wire n_3757;
wire n_11213;
wire n_13519;
wire n_8844;
wire n_6148;
wire n_8995;
wire n_8255;
wire n_5538;
wire n_3666;
wire n_6357;
wire n_8216;
wire n_8693;
wire n_12785;
wire n_3479;
wire n_5499;
wire n_13661;
wire n_9123;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_7811;
wire n_6522;
wire n_12545;
wire n_8669;
wire n_4285;
wire n_7097;
wire n_12531;
wire n_7000;
wire n_2668;
wire n_10486;
wire n_11290;
wire n_2701;
wire n_10357;
wire n_3741;
wire n_9922;
wire n_5582;
wire n_2567;
wire n_9177;
wire n_14348;
wire n_2557;
wire n_5675;
wire n_2755;
wire n_5109;
wire n_7880;
wire n_14130;
wire n_8769;
wire n_9463;
wire n_6713;
wire n_12916;
wire n_8149;
wire n_10067;
wire n_13163;
wire n_12953;
wire n_10698;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_7851;
wire n_13106;
wire n_13874;
wire n_13246;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_10135;
wire n_13776;
wire n_6108;
wire n_12222;
wire n_10260;
wire n_7664;
wire n_12370;
wire n_6100;
wire n_14329;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_11412;
wire n_2829;
wire n_7332;
wire n_14428;
wire n_8990;
wire n_5862;
wire n_7477;
wire n_14617;
wire n_10268;
wire n_8208;
wire n_7468;
wire n_11550;
wire n_12692;
wire n_13640;
wire n_5886;
wire n_9451;
wire n_7714;
wire n_7899;
wire n_8710;
wire n_12976;
wire n_6415;
wire n_8479;
wire n_6783;
wire n_14660;
wire n_4861;
wire n_13984;
wire n_12397;
wire n_8512;
wire n_14524;
wire n_13093;
wire n_9843;
wire n_3673;
wire n_3052;
wire n_9710;
wire n_12634;
wire n_13288;
wire n_9087;
wire n_4621;
wire n_14287;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_7845;
wire n_11619;
wire n_13086;
wire n_14052;
wire n_14216;
wire n_3936;
wire n_5564;
wire n_12613;
wire n_9956;
wire n_3082;
wire n_9079;
wire n_5162;
wire n_5442;
wire n_12946;
wire n_5802;
wire n_9782;
wire n_10049;
wire n_4784;
wire n_14206;
wire n_13012;
wire n_13606;
wire n_12901;
wire n_13449;
wire n_10589;
wire n_3210;
wire n_6340;
wire n_13099;
wire n_14475;
wire n_9950;
wire n_11019;
wire n_14620;
wire n_7858;
wire n_11580;
wire n_3867;
wire n_3397;
wire n_13699;
wire n_12683;
wire n_6103;
wire n_6392;
wire n_6513;
wire n_11642;
wire n_4613;
wire n_2565;
wire n_13389;
wire n_9197;
wire n_6720;
wire n_12286;
wire n_11076;
wire n_11752;
wire n_5883;
wire n_9140;
wire n_14134;
wire n_13995;
wire n_10785;
wire n_13439;
wire n_8401;
wire n_3078;
wire n_6078;
wire n_14122;
wire n_3971;
wire n_12146;
wire n_7680;
wire n_14415;
wire n_5630;
wire n_6666;
wire n_9364;
wire n_9452;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_9362;
wire n_9398;
wire n_13675;
wire n_13483;
wire n_6815;
wire n_14321;
wire n_9203;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_9712;
wire n_9536;
wire n_12054;
wire n_8450;
wire n_9848;
wire n_12081;
wire n_13614;
wire n_14095;
wire n_11202;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_9460;
wire n_7710;
wire n_8788;
wire n_5394;
wire n_14080;
wire n_8324;
wire n_11227;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_13814;
wire n_10381;
wire n_9841;
wire n_14502;
wire n_12557;
wire n_2558;
wire n_9772;
wire n_10147;
wire n_10554;
wire n_2812;
wire n_9057;
wire n_3300;
wire n_7061;
wire n_8104;
wire n_7066;
wire n_9068;
wire n_11860;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_8014;
wire n_12213;
wire n_4122;
wire n_6661;
wire n_10919;
wire n_12646;
wire n_4522;
wire n_10228;
wire n_14159;
wire n_5991;
wire n_8623;
wire n_14077;
wire n_14518;
wire n_4952;
wire n_9634;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_9348;
wire n_11125;
wire n_5920;
wire n_3946;
wire n_13011;
wire n_12737;
wire n_2640;
wire n_6125;
wire n_8651;
wire n_5000;
wire n_10699;
wire n_4634;
wire n_9632;
wire n_4932;
wire n_14358;
wire n_12092;
wire n_11951;
wire n_2983;
wire n_5211;
wire n_9257;
wire n_4089;
wire n_11451;
wire n_11816;
wire n_9500;
wire n_5132;
wire n_3498;
wire n_3513;
wire n_9747;
wire n_9470;
wire n_11508;
wire n_6414;
wire n_5535;
wire n_4506;
wire n_6097;
wire n_14467;
wire n_7783;
wire n_11232;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_10188;
wire n_9591;
wire n_11138;
wire n_14373;
wire n_9049;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_4346;
wire n_13585;
wire n_7003;
wire n_10433;
wire n_8137;
wire n_10231;
wire n_8413;
wire n_10841;
wire n_6302;
wire n_3863;
wire n_10929;
wire n_12642;
wire n_13142;
wire n_3882;
wire n_13974;
wire n_9471;
wire n_3916;
wire n_6922;
wire n_14656;
wire n_3968;
wire n_3675;
wire n_14070;
wire n_10582;
wire n_13494;
wire n_12601;
wire n_2841;
wire n_10719;
wire n_3332;
wire n_8300;
wire n_8069;
wire n_10747;
wire n_7501;
wire n_10934;
wire n_11383;
wire n_9409;
wire n_10711;
wire n_10743;
wire n_11088;
wire n_6432;
wire n_12959;
wire n_7984;
wire n_12899;
wire n_12616;
wire n_2998;
wire n_7366;
wire n_8173;
wire n_10481;
wire n_4359;
wire n_13562;
wire n_13540;
wire n_12919;
wire n_2822;
wire n_7589;
wire n_13568;
wire n_13642;
wire n_4447;
wire n_4293;
wire n_2937;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_9832;
wire n_4039;
wire n_12010;
wire n_12314;
wire n_5793;
wire n_14632;
wire n_6926;
wire n_8091;
wire n_13751;
wire n_3057;
wire n_12394;
wire n_12856;
wire n_5761;
wire n_13465;
wire n_6699;
wire n_12797;
wire n_13683;
wire n_13630;
wire n_3983;
wire n_9067;
wire n_8254;
wire n_8400;
wire n_10141;
wire n_11090;
wire n_14661;
wire n_10305;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_9858;
wire n_7511;
wire n_10936;
wire n_12134;
wire n_13824;
wire n_12730;
wire n_3773;
wire n_3494;
wire n_9482;
wire n_9033;
wire n_6957;
wire n_11429;
wire n_5074;
wire n_14624;
wire n_12735;
wire n_14510;
wire n_7917;
wire n_11908;
wire n_3788;
wire n_3939;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_8368;
wire n_6694;
wire n_9247;
wire n_3260;
wire n_8463;
wire n_9965;
wire n_10425;
wire n_3349;
wire n_6449;
wire n_10862;
wire n_12254;
wire n_14333;
wire n_4348;
wire n_7422;
wire n_9299;
wire n_13357;
wire n_3139;
wire n_8889;
wire n_3801;
wire n_5681;
wire n_9244;
wire n_9785;
wire n_11298;
wire n_14667;
wire n_5261;
wire n_12427;
wire n_12124;
wire n_9195;
wire n_8322;
wire n_11353;
wire n_12494;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_8987;
wire n_13454;
wire n_3653;
wire n_3823;
wire n_9280;
wire n_3403;
wire n_7621;
wire n_9911;
wire n_12051;
wire n_8274;
wire n_13958;
wire n_6594;
wire n_6342;
wire n_6195;
wire n_2716;
wire n_10373;
wire n_6441;
wire n_11116;
wire n_7158;
wire n_7572;
wire n_13637;
wire n_11173;
wire n_2944;
wire n_11660;
wire n_2780;
wire n_3439;
wire n_7500;
wire n_4084;
wire n_12355;
wire n_7985;
wire n_9687;
wire n_4240;
wire n_8657;
wire n_4121;
wire n_3602;
wire n_11567;
wire n_8954;
wire n_2774;
wire n_6354;
wire n_11881;
wire n_10563;
wire n_12458;
wire n_2799;
wire n_8311;
wire n_5748;
wire n_4393;
wire n_11363;
wire n_6662;
wire n_7494;
wire n_9088;
wire n_3984;
wire n_14050;
wire n_8728;
wire n_9580;
wire n_11280;
wire n_9569;
wire n_8994;
wire n_4389;
wire n_6433;
wire n_9680;
wire n_8398;
wire n_6200;
wire n_5641;
wire n_12463;
wire n_12612;
wire n_8407;
wire n_8071;
wire n_13423;
wire n_13046;
wire n_4461;
wire n_2763;
wire n_11636;
wire n_3156;
wire n_10530;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_12798;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_8528;
wire n_14088;
wire n_9227;
wire n_13644;
wire n_5657;
wire n_12510;
wire n_11313;
wire n_14364;
wire n_8475;
wire n_9951;
wire n_9855;
wire n_3579;
wire n_9072;
wire n_12635;
wire n_10102;
wire n_13545;
wire n_3896;
wire n_12537;
wire n_4067;
wire n_13197;
wire n_5244;
wire n_12076;
wire n_5765;
wire n_5114;
wire n_9054;
wire n_4551;
wire n_10117;
wire n_4521;
wire n_13252;
wire n_6956;
wire n_13139;
wire n_10126;
wire n_7587;
wire n_6451;
wire n_12874;
wire n_11920;
wire n_3005;
wire n_7704;
wire n_10604;
wire n_5420;
wire n_6497;
wire n_8511;
wire n_7865;
wire n_5206;
wire n_13356;
wire n_14447;
wire n_4387;
wire n_14237;
wire n_9584;
wire n_9287;
wire n_3186;
wire n_10344;
wire n_10568;
wire n_9459;
wire n_6701;
wire n_2594;
wire n_5298;
wire n_9490;
wire n_10209;
wire n_8867;
wire n_3417;
wire n_8246;
wire n_8558;
wire n_9655;
wire n_13769;
wire n_9846;
wire n_3626;
wire n_12048;
wire n_9593;
wire n_4598;
wire n_4464;
wire n_12072;
wire n_8925;
wire n_5106;
wire n_7881;
wire n_11317;
wire n_9147;
wire n_13339;
wire n_4789;
wire n_3180;
wire n_14433;
wire n_12829;
wire n_3423;
wire n_14672;
wire n_9678;
wire n_10803;
wire n_12132;
wire n_13626;
wire n_11903;
wire n_8641;
wire n_9658;
wire n_10299;
wire n_9560;
wire n_12528;
wire n_9578;
wire n_11813;
wire n_14195;
wire n_5080;
wire n_9396;
wire n_4565;
wire n_7032;
wire n_12745;
wire n_9303;
wire n_3392;
wire n_12371;
wire n_11811;
wire n_12841;
wire n_7198;
wire n_12417;
wire n_6884;
wire n_7752;
wire n_10618;
wire n_10836;
wire n_11378;
wire n_5081;
wire n_8201;
wire n_6921;
wire n_2904;
wire n_12180;
wire n_12049;
wire n_3353;
wire n_2946;
wire n_7953;
wire n_6106;
wire n_14434;
wire n_6876;
wire n_3512;
wire n_9553;
wire n_12603;
wire n_4552;
wire n_8046;
wire n_12978;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_14575;
wire n_10930;
wire n_6172;
wire n_14005;
wire n_9942;
wire n_9805;
wire n_13686;
wire n_4482;
wire n_5957;
wire n_4172;
wire n_12466;
wire n_13842;
wire n_4040;
wire n_8414;
wire n_3024;
wire n_5567;
wire n_8292;
wire n_9138;
wire n_9879;
wire n_5406;
wire n_8647;
wire n_11936;
wire n_6362;
wire n_9213;
wire n_12071;
wire n_4328;
wire n_12982;
wire n_8543;
wire n_14680;
wire n_13459;
wire n_11543;
wire n_11184;
wire n_11795;
wire n_5191;
wire n_11391;
wire n_6067;
wire n_2893;
wire n_11646;
wire n_6833;
wire n_4940;
wire n_9374;
wire n_3161;
wire n_13649;
wire n_14497;
wire n_8331;
wire n_8317;
wire n_7126;
wire n_12578;
wire n_12311;
wire n_11963;
wire n_5867;
wire n_14109;
wire n_13253;
wire n_12985;
wire n_12232;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_12640;
wire n_7496;
wire n_13729;
wire n_6430;
wire n_11435;
wire n_13647;
wire n_9179;
wire n_3977;
wire n_6296;
wire n_10014;
wire n_4112;
wire n_11056;
wire n_10714;
wire n_5602;
wire n_4928;
wire n_7196;
wire n_14241;
wire n_2614;
wire n_12101;
wire n_11120;
wire n_11185;
wire n_7360;
wire n_5428;
wire n_10916;
wire n_6325;
wire n_10895;
wire n_14693;
wire n_12197;
wire n_12497;
wire n_4865;
wire n_6678;
wire n_7982;
wire n_10838;
wire n_13002;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_8174;
wire n_8187;
wire n_8929;
wire n_10108;
wire n_14069;
wire n_4436;
wire n_5822;
wire n_5786;
wire n_3586;
wire n_10661;
wire n_8846;
wire n_5817;
wire n_9277;
wire n_4160;
wire n_6109;
wire n_9611;
wire n_6385;
wire n_12571;
wire n_9744;
wire n_5798;
wire n_10123;
wire n_4137;
wire n_13022;
wire n_8032;
wire n_9504;
wire n_5417;
wire n_14118;
wire n_14445;
wire n_11147;
wire n_10048;
wire n_4545;
wire n_11194;
wire n_8200;
wire n_4758;
wire n_8036;
wire n_9285;
wire n_4840;
wire n_5713;
wire n_9905;
wire n_10963;
wire n_11016;
wire n_12228;
wire n_11146;
wire n_3097;
wire n_13088;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_10788;
wire n_14142;
wire n_9190;
wire n_8586;
wire n_8524;
wire n_11924;
wire n_12540;
wire n_4535;
wire n_7518;
wire n_8828;
wire n_9639;
wire n_10422;
wire n_4385;
wire n_12001;
wire n_7779;
wire n_12059;
wire n_9664;
wire n_13275;
wire n_11830;
wire n_14577;
wire n_4731;
wire n_3748;
wire n_7575;
wire n_11489;
wire n_7073;
wire n_13026;
wire n_8092;
wire n_10471;
wire n_13760;
wire n_12479;
wire n_10979;
wire n_6309;
wire n_8370;
wire n_3732;
wire n_9109;
wire n_10189;
wire n_13820;
wire n_8135;
wire n_12702;
wire n_6519;
wire n_4671;
wire n_14366;
wire n_9741;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_4558;
wire n_10569;
wire n_13116;
wire n_13663;
wire n_10686;
wire n_14055;
wire n_14197;
wire n_8764;
wire n_14454;
wire n_7349;
wire n_9875;
wire n_8502;
wire n_10713;
wire n_11411;
wire n_4319;
wire n_9360;
wire n_6585;
wire n_12211;
wire n_14323;
wire n_7786;
wire n_10913;
wire n_9021;
wire n_8454;
wire n_2929;
wire n_12306;
wire n_4358;
wire n_11145;
wire n_9122;
wire n_7579;
wire n_10099;
wire n_7122;
wire n_12335;
wire n_12637;
wire n_10193;
wire n_14096;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_10203;
wire n_10140;
wire n_13982;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_10920;
wire n_10149;
wire n_11000;
wire n_11712;
wire n_14068;
wire n_4748;
wire n_3167;
wire n_14019;
wire n_7624;
wire n_13405;
wire n_9803;
wire n_13828;
wire n_14397;
wire n_8776;
wire n_10576;
wire n_2857;
wire n_8564;
wire n_12114;
wire n_8343;
wire n_7828;
wire n_14319;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_3050;
wire n_3919;
wire n_8718;
wire n_13102;
wire n_13550;
wire n_14301;
wire n_10682;
wire n_5506;
wire n_7543;
wire n_9659;
wire n_12204;
wire n_13643;
wire n_5475;
wire n_8042;
wire n_7727;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_9013;
wire n_5431;
wire n_9427;
wire n_12325;
wire n_8379;
wire n_8034;
wire n_12143;
wire n_7778;
wire n_5100;
wire n_10225;
wire n_2764;
wire n_9126;
wire n_7019;
wire n_5315;
wire n_2633;
wire n_5752;
wire n_3708;
wire n_2907;
wire n_8441;
wire n_9474;
wire n_14026;
wire n_14362;
wire n_7702;
wire n_14114;
wire n_5746;
wire n_10368;
wire n_4910;
wire n_4724;
wire n_10237;
wire n_14504;
wire n_9538;
wire n_3718;
wire n_6685;
wire n_3390;
wire n_8569;
wire n_9574;
wire n_10531;
wire n_12032;
wire n_4666;
wire n_4082;
wire n_3140;
wire n_12066;
wire n_14471;
wire n_8592;
wire n_8865;
wire n_3976;
wire n_3381;
wire n_2813;
wire n_7952;
wire n_11170;
wire n_7347;
wire n_9450;
wire n_3736;
wire n_10031;
wire n_4466;
wire n_6016;
wire n_9998;
wire n_13963;
wire n_3955;
wire n_5366;
wire n_11523;
wire n_5322;
wire n_11121;
wire n_12176;
wire n_5414;
wire n_11805;
wire n_3086;
wire n_13266;
wire n_7791;
wire n_3165;
wire n_8362;
wire n_6971;
wire n_10847;
wire n_3336;
wire n_8632;
wire n_10035;
wire n_14242;
wire n_14523;
wire n_7739;
wire n_12740;
wire n_7945;
wire n_9372;
wire n_9045;
wire n_8361;
wire n_9657;
wire n_7656;
wire n_11457;
wire n_5903;
wire n_7199;
wire n_10107;
wire n_3635;
wire n_11725;
wire n_3541;
wire n_10283;
wire n_5151;
wire n_5307;
wire n_3605;
wire n_4721;
wire n_9904;
wire n_12344;
wire n_9924;
wire n_9159;
wire n_8561;
wire n_6549;
wire n_8611;
wire n_9326;
wire n_8410;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_6658;
wire n_11694;
wire n_5369;
wire n_9476;
wire n_6683;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_5912;
wire n_11540;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_10050;
wire n_11058;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_8878;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_12203;
wire n_11403;
wire n_8492;
wire n_9301;
wire n_14099;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_10392;
wire n_14041;
wire n_12769;
wire n_8888;
wire n_6820;
wire n_5446;
wire n_11741;
wire n_7610;
wire n_7107;
wire n_11245;
wire n_4561;
wire n_14225;
wire n_3291;
wire n_7456;
wire n_9382;
wire n_11784;
wire n_8095;
wire n_11365;
wire n_13291;
wire n_9921;
wire n_7369;
wire n_9325;
wire n_9945;
wire n_9643;
wire n_7548;
wire n_11005;
wire n_13016;
wire n_2578;
wire n_12820;
wire n_8735;
wire n_7598;
wire n_7250;
wire n_8808;
wire n_9201;
wire n_8902;
wire n_7823;
wire n_9771;
wire n_8833;
wire n_14605;
wire n_12869;
wire n_4715;
wire n_6157;
wire n_8796;
wire n_2715;
wire n_14413;
wire n_2665;
wire n_4879;
wire n_13435;
wire n_8794;
wire n_12689;
wire n_11074;
wire n_5044;
wire n_3755;
wire n_4536;
wire n_9894;
wire n_9274;
wire n_11141;
wire n_12750;
wire n_8549;
wire n_14161;
wire n_6676;
wire n_4304;
wire n_10095;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_14285;
wire n_11102;
wire n_10716;
wire n_12171;
wire n_14000;
wire n_10088;
wire n_11238;
wire n_11406;
wire n_2854;
wire n_10443;
wire n_10488;
wire n_7525;
wire n_4418;
wire n_7924;
wire n_3341;
wire n_11103;
wire n_12420;
wire n_9232;
wire n_8690;
wire n_4125;
wire n_5390;
wire n_12954;
wire n_5351;
wire n_5267;
wire n_11852;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_12500;
wire n_8593;
wire n_11837;
wire n_10912;
wire n_13501;
wire n_10469;
wire n_13533;
wire n_9649;
wire n_11684;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_12112;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_4412;
wire n_6923;
wire n_7649;
wire n_8195;
wire n_8009;
wire n_8588;
wire n_9839;
wire n_10887;
wire n_3358;
wire n_12004;
wire n_6704;
wire n_7634;
wire n_9090;
wire n_7406;
wire n_13520;
wire n_4682;
wire n_9346;
wire n_11012;
wire n_6673;
wire n_14480;
wire n_9696;
wire n_11041;
wire n_14181;
wire n_10742;
wire n_14024;
wire n_11798;
wire n_12614;
wire n_13165;
wire n_9996;
wire n_6534;
wire n_9968;
wire n_8805;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_4957;
wire n_4855;
wire n_3289;
wire n_6127;
wire n_9383;
wire n_9498;
wire n_10405;
wire n_6246;
wire n_10390;
wire n_11978;
wire n_10989;
wire n_9836;
wire n_5005;
wire n_14570;
wire n_14702;
wire n_11827;
wire n_10328;
wire n_13315;
wire n_10692;
wire n_6126;
wire n_7372;
wire n_8596;
wire n_9938;
wire n_12912;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_10867;
wire n_6841;
wire n_11847;
wire n_10206;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_11281;
wire n_2658;
wire n_12957;
wire n_5624;
wire n_10092;
wire n_3620;
wire n_4601;
wire n_4518;
wire n_5474;
wire n_2767;
wire n_7009;
wire n_3376;
wire n_11772;
wire n_9743;
wire n_9121;
wire n_7371;
wire n_13448;
wire n_11237;
wire n_9509;
wire n_3123;
wire n_5447;
wire n_12153;
wire n_2692;
wire n_12005;
wire n_7463;
wire n_9621;
wire n_4102;
wire n_10738;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_11851;
wire n_9158;
wire n_2862;
wire n_4325;
wire n_14239;
wire n_14501;
wire n_2645;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_12586;
wire n_11993;
wire n_5962;
wire n_4413;
wire n_11131;
wire n_12221;
wire n_8627;
wire n_14318;
wire n_11432;
wire n_12302;
wire n_3307;
wire n_8945;
wire n_9142;
wire n_3251;
wire n_3288;
wire n_13628;
wire n_2833;
wire n_9216;
wire n_9189;
wire n_6723;
wire n_7398;
wire n_3723;
wire n_7941;
wire n_4135;
wire n_9563;
wire n_12757;
wire n_13010;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_13251;
wire n_8858;
wire n_12107;
wire n_11738;
wire n_11595;
wire n_3880;
wire n_13504;
wire n_13521;
wire n_14404;
wire n_12695;
wire n_11512;
wire n_5801;
wire n_14163;
wire n_3904;
wire n_12349;
wire n_6054;
wire n_13703;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_13161;
wire n_7011;
wire n_10813;
wire n_3405;
wire n_14076;
wire n_10986;
wire n_11603;
wire n_6393;
wire n_14291;
wire n_12380;
wire n_7074;
wire n_10853;
wire n_8916;
wire n_10899;
wire n_11707;
wire n_11728;
wire n_13352;
wire n_11521;
wire n_13309;
wire n_5465;
wire n_12577;
wire n_10575;
wire n_8745;
wire n_3532;
wire n_5154;
wire n_14388;
wire n_5721;
wire n_2609;
wire n_8169;
wire n_6184;
wire n_8018;
wire n_11802;
wire n_9984;
wire n_4138;
wire n_3131;
wire n_7083;
wire n_8260;
wire n_12723;
wire n_10334;
wire n_14153;
wire n_12135;
wire n_2882;
wire n_14674;
wire n_7143;
wire n_7701;
wire n_11688;
wire n_13484;
wire n_8688;
wire n_9794;
wire n_7969;
wire n_10726;
wire n_8279;
wire n_4384;
wire n_8793;
wire n_4639;
wire n_12864;
wire n_13486;
wire n_10388;
wire n_4577;
wire n_6312;
wire n_13478;
wire n_7683;
wire n_9550;
wire n_13108;
wire n_11042;
wire n_12570;
wire n_14124;
wire n_10510;
wire n_14344;
wire n_7669;
wire n_8298;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_11696;
wire n_6438;
wire n_11761;
wire n_3926;
wire n_4481;
wire n_5087;
wire n_10635;
wire n_11681;
wire n_2938;
wire n_7209;
wire n_13429;
wire n_6193;
wire n_3992;
wire n_13897;
wire n_8023;
wire n_9319;
wire n_7330;
wire n_6007;
wire n_13374;
wire n_13182;
wire n_6734;
wire n_10852;
wire n_6535;
wire n_13789;
wire n_8053;
wire n_11407;
wire n_8059;
wire n_9871;
wire n_14354;
wire n_6879;
wire n_9562;
wire n_9896;
wire n_9612;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_9698;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_9528;
wire n_10241;
wire n_4620;
wire n_5397;
wire n_6255;
wire n_6457;
wire n_13690;
wire n_9272;
wire n_13055;
wire n_14379;
wire n_9955;
wire n_9645;
wire n_4924;
wire n_4044;
wire n_8372;
wire n_6270;
wire n_14283;
wire n_8737;
wire n_9731;
wire n_10026;
wire n_5996;
wire n_13577;
wire n_5566;
wire n_9697;
wire n_3304;
wire n_7288;
wire n_10772;
wire n_4388;
wire n_13098;
wire n_10901;
wire n_7362;
wire n_7237;
wire n_7082;
wire n_8988;
wire n_3247;
wire n_10664;
wire n_7131;
wire n_6276;
wire n_12328;
wire n_13839;
wire n_9642;
wire n_8723;
wire n_11189;
wire n_12559;
wire n_9929;
wire n_9050;
wire n_4406;
wire n_4271;
wire n_12056;
wire n_13898;
wire n_7042;
wire n_9859;
wire n_8419;
wire n_2809;
wire n_10767;
wire n_10320;
wire n_5652;
wire n_13380;
wire n_8893;
wire n_5805;
wire n_7304;
wire n_11910;
wire n_6266;
wire n_3301;
wire n_12109;
wire n_2910;
wire n_14457;
wire n_9531;
wire n_10521;
wire n_3785;
wire n_5492;
wire n_8077;
wire n_11242;
wire n_5501;
wire n_12917;
wire n_6934;
wire n_13188;
wire n_14179;
wire n_13362;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_11361;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_8826;
wire n_3178;
wire n_12058;
wire n_11894;
wire n_13819;
wire n_7023;
wire n_10872;
wire n_13990;
wire n_9732;
wire n_5842;
wire n_5758;
wire n_12083;
wire n_9685;
wire n_12529;
wire n_3100;
wire n_3721;
wire n_10374;
wire n_11253;
wire n_13983;
wire n_12045;
wire n_13193;
wire n_7404;
wire n_3389;
wire n_10345;
wire n_8959;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_12471;
wire n_4973;
wire n_13802;
wire n_13781;
wire n_7981;
wire n_4792;
wire n_13037;
wire n_3537;
wire n_4402;
wire n_14252;
wire n_12188;
wire n_5473;
wire n_12575;
wire n_10601;
wire n_14698;
wire n_11623;
wire n_8712;
wire n_12473;
wire n_10372;
wire n_6352;
wire n_11124;
wire n_14295;
wire n_2941;
wire n_4286;
wire n_9378;
wire n_3638;
wire n_6211;
wire n_10448;
wire n_8109;
wire n_10301;
wire n_11977;
wire n_3576;
wire n_10074;
wire n_12040;
wire n_14025;
wire n_13127;
wire n_9389;
wire n_12598;
wire n_5562;
wire n_4858;
wire n_6093;
wire n_5370;
wire n_10001;
wire n_13561;
wire n_7378;
wire n_9623;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7877;
wire n_14336;
wire n_11351;
wire n_7787;
wire n_7836;
wire n_8515;
wire n_8725;
wire n_12626;
wire n_11094;
wire n_10960;
wire n_10712;
wire n_8007;
wire n_13911;
wire n_14313;
wire n_4318;
wire n_13961;
wire n_13343;
wire n_12546;
wire n_8910;
wire n_5227;
wire n_14091;
wire n_10100;
wire n_5902;
wire n_9164;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_11366;
wire n_2793;
wire n_5282;
wire n_9387;
wire n_8301;
wire n_6764;
wire n_7871;
wire n_14512;
wire n_13539;
wire n_10162;
wire n_2639;
wire n_9840;
wire n_7016;
wire n_4738;
wire n_12100;
wire n_2603;
wire n_8892;
wire n_11399;
wire n_9637;
wire n_5386;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_8252;
wire n_4526;
wire n_4105;
wire n_10535;
wire n_10674;
wire n_12676;
wire n_13584;
wire n_3663;
wire n_9491;
wire n_7563;
wire n_6955;
wire n_10337;
wire n_10774;
wire n_5952;
wire n_7180;
wire n_13107;
wire n_10407;
wire n_14655;
wire n_10577;
wire n_14481;
wire n_13778;
wire n_8972;
wire n_14531;
wire n_8494;
wire n_12999;
wire n_10264;
wire n_6569;
wire n_7919;
wire n_13740;
wire n_9992;
wire n_14606;
wire n_14089;
wire n_2966;
wire n_8278;
wire n_3431;
wire n_8180;
wire n_11549;
wire n_14437;
wire n_12362;
wire n_3355;
wire n_7031;
wire n_13913;
wire n_13367;
wire n_5716;
wire n_10313;
wire n_10843;
wire n_12983;
wire n_14003;
wire n_8941;
wire n_10771;
wire n_8891;
wire n_3897;
wire n_7103;
wire n_12360;
wire n_13570;
wire n_6605;
wire n_10724;
wire n_5888;
wire n_9266;
wire n_4005;
wire n_14409;
wire n_8270;
wire n_8231;
wire n_4181;
wire n_2597;
wire n_11983;
wire n_6832;
wire n_12313;
wire n_12604;
wire n_5980;
wire n_8683;
wire n_9391;
wire n_4092;
wire n_12558;
wire n_10445;
wire n_4875;
wire n_7771;
wire n_8903;
wire n_4255;
wire n_13284;
wire n_2758;
wire n_6544;
wire n_8810;
wire n_12596;
wire n_6469;
wire n_12840;
wire n_5036;
wire n_11119;
wire n_12696;
wire n_6332;
wire n_10863;
wire n_10958;
wire n_11215;
wire n_13730;
wire n_5790;
wire n_7130;
wire n_10174;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_13960;
wire n_6310;
wire n_8932;
wire n_8264;
wire n_12435;
wire n_9695;
wire n_7134;
wire n_3042;
wire n_8288;
wire n_13411;
wire n_11954;
wire n_14629;
wire n_11526;
wire n_13438;
wire n_14010;
wire n_11591;
wire n_10403;
wire n_11972;
wire n_4142;
wire n_5118;
wire n_9834;
wire n_5485;
wire n_9901;
wire n_10076;
wire n_5525;
wire n_7102;
wire n_10015;
wire n_6259;
wire n_3004;
wire n_14432;
wire n_5271;
wire n_4849;
wire n_13410;
wire n_7133;
wire n_9800;
wire n_10745;
wire n_6651;
wire n_6289;
wire n_3838;
wire n_9255;
wire n_8882;
wire n_14308;
wire n_12460;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_12733;
wire n_8388;
wire n_5445;
wire n_2734;
wire n_8067;
wire n_13600;
wire n_8385;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_8670;
wire n_4504;
wire n_10460;
wire n_14299;
wire n_14215;
wire n_3598;
wire n_4917;
wire n_7706;
wire n_7813;
wire n_8142;
wire n_13332;
wire n_14265;
wire n_13942;
wire n_7992;
wire n_9085;
wire n_7643;
wire n_11204;
wire n_6836;
wire n_12939;
wire n_3273;
wire n_9120;
wire n_2918;
wire n_6595;
wire n_10415;
wire n_11302;
wire n_9899;
wire n_12374;
wire n_9136;
wire n_12261;
wire n_6186;
wire n_11561;
wire n_10227;
wire n_2641;
wire n_13490;
wire n_14198;
wire n_2580;
wire n_7628;
wire n_13381;
wire n_5628;
wire n_5245;
wire n_9436;
wire n_4489;
wire n_14013;
wire n_11385;
wire n_12065;
wire n_13204;
wire n_5329;
wire n_12275;
wire n_8224;
wire n_5472;
wire n_6035;
wire n_9042;
wire n_10884;
wire n_13375;
wire n_7236;
wire n_9570;
wire n_4833;
wire n_3394;
wire n_9239;
wire n_6405;
wire n_8345;
wire n_11054;
wire n_11777;
wire n_9644;
wire n_5850;
wire n_9343;
wire n_8614;
wire n_8242;
wire n_6786;
wire n_4564;
wire n_8299;
wire n_9131;
wire n_13286;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_9060;
wire n_9792;
wire n_3581;
wire n_8110;
wire n_5072;
wire n_8529;
wire n_3778;
wire n_14204;
wire n_13384;
wire n_11325;
wire n_10801;
wire n_6769;
wire n_10325;
wire n_13013;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_8951;
wire n_11217;
wire n_4080;
wire n_13582;
wire n_12752;
wire n_10327;
wire n_8700;
wire n_6766;
wire n_4185;
wire n_5940;
wire n_3001;
wire n_14157;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_11651;
wire n_6232;
wire n_13255;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_7802;
wire n_7519;
wire n_10505;
wire n_3932;
wire n_2577;
wire n_12979;
wire n_14140;
wire n_7457;
wire n_11196;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_5860;
wire n_11672;
wire n_11557;
wire n_9982;
wire n_11552;
wire n_6416;
wire n_13682;
wire n_2933;
wire n_8468;
wire n_9031;
wire n_12715;
wire n_12910;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_11084;
wire n_12787;
wire n_8933;
wire n_6214;
wire n_3952;
wire n_9006;
wire n_8636;
wire n_10408;
wire n_11442;
wire n_9221;
wire n_13424;
wire n_4365;
wire n_3584;
wire n_14102;
wire n_4349;
wire n_3446;
wire n_10514;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_8378;
wire n_6143;
wire n_14603;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_10091;
wire n_11195;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_10562;
wire n_10586;
wire n_10893;
wire n_8283;
wire n_6225;
wire n_4373;
wire n_7914;
wire n_8860;
wire n_2664;
wire n_12401;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_14104;
wire n_4390;
wire n_10593;
wire n_13304;
wire n_11517;
wire n_7892;
wire n_4107;
wire n_12722;
wire n_13716;
wire n_9523;
wire n_10821;
wire n_4380;
wire n_4609;
wire n_4361;
wire n_7325;
wire n_11918;
wire n_14561;
wire n_13460;
wire n_4453;
wire n_6219;
wire n_7674;
wire n_8686;
wire n_13590;
wire n_12712;
wire n_10961;
wire n_6175;
wire n_6445;
wire n_9829;
wire n_8563;
wire n_11077;
wire n_4571;
wire n_13914;
wire n_3137;
wire n_11579;
wire n_10197;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_8493;
wire n_6198;
wire n_5172;
wire n_14119;
wire n_13670;
wire n_13148;
wire n_10950;
wire n_6499;
wire n_9411;
wire n_12209;
wire n_7983;
wire n_5311;
wire n_8765;
wire n_14168;
wire n_14494;
wire n_13452;
wire n_14506;
wire n_5164;
wire n_11640;
wire n_13688;
wire n_4964;
wire n_10180;
wire n_9153;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_10079;
wire n_7361;
wire n_11656;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_11845;
wire n_11679;
wire n_14007;
wire n_13671;
wire n_2982;
wire n_8653;
wire n_5495;
wire n_6281;
wire n_13005;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_13313;
wire n_5547;
wire n_4693;
wire n_10361;
wire n_14154;
wire n_11635;
wire n_8601;
wire n_9675;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_8333;
wire n_9571;
wire n_9097;
wire n_12323;
wire n_12835;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_10075;
wire n_11572;
wire n_9789;
wire n_2674;
wire n_13387;
wire n_5820;
wire n_13068;
wire n_11529;
wire n_9925;
wire n_7309;
wire n_7119;
wire n_14426;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_13173;
wire n_10012;
wire n_3902;
wire n_14351;
wire n_12873;
wire n_12830;
wire n_12015;
wire n_12348;
wire n_12767;
wire n_3244;
wire n_10939;
wire n_2562;
wire n_3112;
wire n_10008;
wire n_11384;
wire n_14382;
wire n_9511;
wire n_9795;
wire n_3196;
wire n_11134;
wire n_8708;
wire n_10503;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_10111;
wire n_10798;
wire n_10982;
wire n_4678;
wire n_11630;
wire n_12867;
wire n_13479;
wire n_5301;
wire n_13203;
wire n_13263;
wire n_13710;
wire n_5126;
wire n_13211;
wire n_8659;
wire n_14700;
wire n_6732;
wire n_8759;
wire n_3488;
wire n_9622;
wire n_12198;
wire n_9761;
wire n_2744;
wire n_6817;
wire n_5776;
wire n_7646;
wire n_14249;
wire n_9954;
wire n_14530;
wire n_3779;
wire n_13848;
wire n_6982;
wire n_12617;
wire n_7291;
wire n_10669;
wire n_8790;
wire n_13052;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_8832;
wire n_13282;
wire n_8305;
wire n_3834;
wire n_4303;
wire n_3923;
wire n_5603;
wire n_8453;
wire n_6560;
wire n_6634;
wire n_14275;
wire n_5348;
wire n_12666;
wire n_9847;
wire n_13818;
wire n_4868;
wire n_7017;
wire n_13846;
wire n_12845;
wire n_11617;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_13312;
wire n_4465;
wire n_9640;
wire n_8127;
wire n_13565;
wire n_2596;
wire n_5217;
wire n_8337;
wire n_9115;
wire n_5558;
wire n_3986;
wire n_3725;
wire n_7861;
wire n_12047;
wire n_10190;
wire n_12411;
wire n_9534;
wire n_4026;
wire n_13788;
wire n_4245;
wire n_11422;
wire n_5520;
wire n_7889;
wire n_13295;
wire n_3894;
wire n_12594;
wire n_10542;
wire n_14349;
wire n_5909;
wire n_4852;
wire n_7554;
wire n_3202;
wire n_11289;
wire n_8508;
wire n_4290;
wire n_4945;
wire n_11376;
wire n_5750;
wire n_7648;
wire n_8968;
wire n_10752;
wire n_5654;
wire n_11157;
wire n_10868;
wire n_11013;
wire n_2819;
wire n_9594;
wire n_11017;
wire n_7653;
wire n_11765;
wire n_6400;
wire n_12885;
wire n_11307;
wire n_7846;
wire n_3547;
wire n_4014;
wire n_8347;
wire n_5554;
wire n_9503;
wire n_12811;
wire n_3045;
wire n_9919;
wire n_13346;
wire n_13331;
wire n_5135;
wire n_7551;
wire n_11793;
wire n_11574;
wire n_4599;
wire n_13307;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_10017;
wire n_13574;
wire n_12073;
wire n_8093;
wire n_8899;
wire n_9385;
wire n_12913;
wire n_13027;
wire n_14563;
wire n_5448;
wire n_14357;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_11836;
wire n_5412;
wire n_8481;
wire n_14169;
wire n_3249;
wire n_3483;
wire n_6851;
wire n_6621;
wire n_4046;
wire n_11747;
wire n_4701;
wire n_2915;
wire n_7606;
wire n_9963;
wire n_7420;
wire n_10572;
wire n_11193;
wire n_9885;
wire n_8115;
wire n_4869;
wire n_13939;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_11670;
wire n_14042;
wire n_10642;
wire n_2719;
wire n_10115;
wire n_10517;
wire n_14429;
wire n_14098;
wire n_13289;
wire n_10247;
wire n_2876;
wire n_13851;
wire n_13852;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_12585;
wire n_12451;
wire n_12029;
wire n_12963;
wire n_13616;
wire n_6226;
wire n_14490;
wire n_9827;
wire n_12169;
wire n_3033;
wire n_12801;
wire n_9182;
wire n_10620;
wire n_8182;
wire n_9426;
wire n_9293;
wire n_2824;
wire n_10065;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_11762;
wire n_14030;
wire n_14500;
wire n_7896;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_9581;
wire n_5900;
wire n_8629;
wire n_12657;
wire n_8186;
wire n_7319;
wire n_11758;
wire n_3619;
wire n_6158;
wire n_13366;
wire n_9400;
wire n_4013;
wire n_10744;
wire n_3434;
wire n_9246;
wire n_4342;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_3853;
wire n_8233;
wire n_4382;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_9445;
wire n_8282;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_7516;
wire n_6928;
wire n_6317;
wire n_10609;
wire n_13860;
wire n_11958;
wire n_6707;
wire n_10009;
wire n_13847;
wire n_7244;
wire n_11314;
wire n_4626;
wire n_12210;
wire n_10072;
wire n_12443;
wire n_12699;
wire n_7625;
wire n_8750;
wire n_10130;
wire n_4997;
wire n_8183;
wire n_13657;
wire n_5065;
wire n_9104;
wire n_13450;
wire n_6806;
wire n_10956;
wire n_7991;
wire n_8637;
wire n_4638;
wire n_2786;
wire n_9542;
wire n_11490;
wire n_11515;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_8792;
wire n_6835;
wire n_7286;
wire n_3517;
wire n_13610;
wire n_6269;
wire n_7857;
wire n_13871;
wire n_7970;
wire n_9302;
wire n_8258;
wire n_10829;
wire n_3719;
wire n_7154;
wire n_11356;
wire n_12781;
wire n_10506;
wire n_3526;
wire n_3888;
wire n_9960;
wire n_12573;
wire n_13326;
wire n_3198;
wire n_5295;
wire n_8416;
wire n_8390;
wire n_13881;
wire n_11678;
wire n_12744;
wire n_6088;
wire n_10236;
wire n_11374;
wire n_14519;
wire n_11176;
wire n_7194;
wire n_4841;
wire n_11402;
wire n_4683;
wire n_5173;
wire n_11162;
wire n_2873;
wire n_10002;
wire n_8696;
wire n_9185;
wire n_9601;
wire n_13137;
wire n_13226;
wire n_3330;
wire n_3514;
wire n_11771;
wire n_5655;
wire n_3383;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_3905;
wire n_7163;
wire n_13431;
wire n_14402;
wire n_14507;
wire n_14020;
wire n_3797;
wire n_13552;
wire n_13164;
wire n_7027;
wire n_3416;
wire n_8552;
wire n_12006;
wire n_4600;
wire n_5861;
wire n_6964;
wire n_3943;
wire n_10855;
wire n_3145;
wire n_14389;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_9403;
wire n_14558;
wire n_11322;
wire n_6316;
wire n_8619;
wire n_7068;
wire n_11484;
wire n_9972;
wire n_11711;
wire n_13227;
wire n_2908;
wire n_8594;
wire n_9878;
wire n_14541;
wire n_10139;
wire n_14183;
wire n_4106;
wire n_9541;
wire n_10941;
wire n_14689;
wire n_12548;
wire n_8162;
wire n_9735;
wire n_9576;
wire n_14528;
wire n_4549;
wire n_7327;
wire n_12727;
wire n_12240;
wire n_13045;
wire n_6610;
wire n_13620;
wire n_5998;
wire n_8318;
wire n_4702;
wire n_5102;
wire n_9974;
wire n_4954;
wire n_10992;
wire n_4491;
wire n_2906;
wire n_8425;
wire n_6752;
wire n_13001;
wire n_6959;
wire n_9704;
wire n_6250;
wire n_13919;
wire n_11392;
wire n_12372;
wire n_3283;
wire n_11803;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_11912;
wire n_13862;
wire n_13784;
wire n_7864;
wire n_11139;
wire n_3451;
wire n_10650;
wire n_8051;
wire n_4734;
wire n_11021;
wire n_6675;
wire n_7955;
wire n_2832;
wire n_5827;
wire n_9039;
wire n_12914;
wire n_7384;
wire n_12844;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_12952;
wire n_5678;
wire n_6561;
wire n_11379;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_13271;
wire n_7512;
wire n_7814;
wire n_12276;
wire n_12096;
wire n_8389;
wire n_4515;
wire n_10417;
wire n_10029;
wire n_12150;
wire n_14271;
wire n_13595;
wire n_8620;
wire n_10125;
wire n_5555;
wire n_13757;
wire n_8886;
wire n_4809;
wire n_7152;
wire n_4012;
wire n_10253;
wire n_11899;
wire n_13761;
wire n_5212;
wire n_4760;
wire n_13190;
wire n_13136;
wire n_6823;
wire n_10693;
wire n_3606;
wire n_14461;
wire n_7062;
wire n_7090;
wire n_12449;
wire n_8202;
wire n_13633;
wire n_11966;
wire n_14205;
wire n_5815;
wire n_4320;
wire n_12118;
wire n_10599;
wire n_5084;
wire n_7223;
wire n_14266;
wire n_12770;
wire n_5251;
wire n_8755;
wire n_13174;
wire n_8668;
wire n_5965;
wire n_4980;
wire n_3324;
wire n_10977;
wire n_13528;
wire n_6796;
wire n_8979;
wire n_5407;
wire n_2988;
wire n_12814;
wire n_11553;
wire n_4560;
wire n_14064;
wire n_14322;
wire n_13220;
wire n_12009;
wire n_14466;
wire n_13456;
wire n_13916;
wire n_7761;
wire n_10947;
wire n_8141;
wire n_10386;
wire n_5042;
wire n_3230;
wire n_3793;
wire n_8199;
wire n_12826;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_10267;
wire n_6090;
wire n_5368;
wire n_10401;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_3183;
wire n_9908;
wire n_11127;
wire n_8004;
wire n_11926;
wire n_8383;
wire n_3607;
wire n_9864;
wire n_9688;
wire n_12144;
wire n_3613;
wire n_2885;
wire n_2616;
wire n_7388;
wire n_7056;
wire n_10428;
wire n_14585;
wire n_10212;
wire n_7437;
wire n_11460;
wire n_6489;
wire n_11486;
wire n_9023;
wire n_5310;
wire n_2769;
wire n_8895;
wire n_8680;
wire n_14208;
wire n_4987;
wire n_6714;
wire n_8394;
wire n_7849;
wire n_10539;
wire n_14152;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_7417;
wire n_2739;
wire n_12937;
wire n_3962;
wire n_11148;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_10728;
wire n_12312;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_6620;
wire n_6791;
wire n_4540;
wire n_9220;
wire n_13929;
wire n_6821;
wire n_9317;
wire n_12580;
wire n_13965;
wire n_13796;
wire n_5588;
wire n_3854;
wire n_8198;
wire n_9993;
wire n_10879;
wire n_13474;
wire n_8665;
wire n_12393;
wire n_6583;
wire n_10545;
wire n_3652;
wire n_12201;
wire n_7859;
wire n_3449;
wire n_13240;
wire n_13187;
wire n_13594;
wire n_3089;
wire n_4854;
wire n_9561;
wire n_10516;
wire n_14640;
wire n_9444;
wire n_10497;
wire n_8017;
wire n_11675;
wire n_5477;
wire n_2727;
wire n_10705;
wire n_7523;
wire n_12082;
wire n_13966;
wire n_11032;
wire n_5234;
wire n_14035;
wire n_12322;
wire n_6890;
wire n_9184;
wire n_10432;
wire n_11454;
wire n_7559;
wire n_14345;
wire n_9037;
wire n_7576;
wire n_6988;
wire n_8303;
wire n_10779;
wire n_11554;
wire n_5871;
wire n_11988;
wire n_13981;
wire n_4747;
wire n_14647;
wire n_8000;
wire n_11197;
wire n_14286;
wire n_3472;
wire n_14686;
wire n_6052;
wire n_7769;
wire n_11416;
wire n_9505;
wire n_9193;
wire n_14360;
wire n_7257;
wire n_3126;
wire n_12986;
wire n_2759;
wire n_6973;
wire n_10869;
wire n_8852;
wire n_5007;
wire n_8709;
wire n_4881;
wire n_10314;
wire n_10504;
wire n_6488;
wire n_4495;
wire n_3958;
wire n_10687;
wire n_13691;
wire n_4737;
wire n_9218;
wire n_11341;
wire n_9755;
wire n_4357;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_11045;
wire n_3191;
wire n_12373;
wire n_7005;
wire n_12741;
wire n_5334;
wire n_3562;
wire n_8782;
wire n_7081;
wire n_10882;
wire n_7742;
wire n_5253;
wire n_10293;
wire n_3588;
wire n_6280;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_9506;
wire n_9162;
wire n_13629;
wire n_3095;
wire n_7341;
wire n_5792;
wire n_13155;
wire n_14581;
wire n_3698;
wire n_4513;
wire n_11569;
wire n_13152;
wire n_10256;
wire n_4775;
wire n_6256;
wire n_2620;
wire n_8716;
wire n_12677;
wire n_8250;
wire n_7264;
wire n_12412;
wire n_7842;
wire n_14315;
wire n_12181;
wire n_12833;
wire n_6648;
wire n_9415;
wire n_10298;
wire n_12115;
wire n_12631;
wire n_7492;
wire n_13194;
wire n_13546;
wire n_6649;
wire n_8714;
wire n_8357;
wire n_12567;
wire n_3093;
wire n_12175;
wire n_2970;
wire n_6910;
wire n_9990;
wire n_3885;
wire n_8466;
wire n_4264;
wire n_5954;
wire n_9015;
wire n_10326;
wire n_13446;
wire n_10235;
wire n_3192;
wire n_4709;
wire n_6431;
wire n_8589;
wire n_12754;
wire n_4223;
wire n_3250;
wire n_14141;
wire n_12455;
wire n_3538;
wire n_13363;
wire n_3915;
wire n_11990;
wire n_8266;
wire n_3839;
wire n_8587;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_10725;
wire n_10274;
wire n_13728;
wire n_13601;
wire n_3875;
wire n_4029;
wire n_8876;
wire n_11541;
wire n_9214;
wire n_4206;
wire n_12340;
wire n_4099;
wire n_10799;
wire n_8922;
wire n_11680;
wire n_10090;
wire n_3120;
wire n_6512;
wire n_12686;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_9070;
wire n_8498;
wire n_4794;
wire n_9933;
wire n_4843;
wire n_12734;
wire n_5580;
wire n_5215;
wire n_12331;
wire n_4763;
wire n_3937;
wire n_10874;
wire n_9339;
wire n_11596;
wire n_9991;
wire n_12880;
wire n_9486;
wire n_8457;
wire n_6243;
wire n_14113;
wire n_5795;
wire n_10763;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_10266;
wire n_8267;
wire n_12184;
wire n_12425;
wire n_7051;
wire n_13918;
wire n_11180;
wire n_6773;
wire n_10290;
wire n_6231;
wire n_12472;
wire n_13048;
wire n_12266;
wire n_7503;
wire n_4838;
wire n_4795;
wire n_12432;
wire n_8124;
wire n_3604;
wire n_8545;
wire n_5430;
wire n_6041;
wire n_8526;
wire n_12300;
wire n_13593;
wire n_8319;
wire n_7997;
wire n_12527;
wire n_5659;
wire n_11839;
wire n_9279;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_10732;
wire n_5195;
wire n_12110;
wire n_13744;
wire n_3176;
wire n_9790;
wire n_11404;
wire n_3792;
wire n_7950;
wire n_11548;
wire n_6323;
wire n_13515;
wire n_5720;
wire n_4267;
wire n_8581;
wire n_12122;
wire n_10873;
wire n_8214;
wire n_7793;
wire n_9053;
wire n_8516;
wire n_12310;
wire n_5598;
wire n_2753;
wire n_11343;
wire n_3021;
wire n_8989;
wire n_13028;
wire n_7746;
wire n_11362;
wire n_4352;
wire n_2712;
wire n_3805;
wire n_3912;
wire n_11007;
wire n_3950;
wire n_7570;
wire n_9650;
wire n_9880;
wire n_11497;
wire n_2898;
wire n_10720;
wire n_6912;
wire n_3567;
wire n_14574;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_14014;
wire n_12827;
wire n_14078;
wire n_10220;
wire n_9217;
wire n_9499;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_13467;
wire n_13245;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_10081;
wire n_12804;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_9282;
wire n_7894;
wire n_10145;
wire n_11347;
wire n_7957;
wire n_8262;
wire n_10167;
wire n_5530;
wire n_12892;
wire n_12656;
wire n_6718;
wire n_8289;
wire n_13804;
wire n_5809;
wire n_10447;
wire n_12418;
wire n_7531;
wire n_7121;
wire n_6410;
wire n_12448;
wire n_12219;
wire n_12729;
wire n_13549;
wire n_13921;
wire n_6473;
wire n_8087;
wire n_4056;
wire n_10238;
wire n_13345;
wire n_4806;
wire n_11029;
wire n_7961;
wire n_9920;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_9948;
wire n_4462;
wire n_5299;
wire n_13216;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_11226;
wire n_8863;
wire n_9371;
wire n_4517;
wire n_2896;
wire n_8701;
wire n_4043;
wire n_13036;
wire n_3170;
wire n_9237;
wire n_13398;
wire n_6857;
wire n_8705;
wire n_14148;
wire n_9815;
wire n_3415;
wire n_10292;
wire n_12644;
wire n_6975;
wire n_10820;
wire n_7763;
wire n_13258;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_7703;
wire n_11760;
wire n_13827;
wire n_7928;
wire n_4234;
wire n_10395;
wire n_12576;
wire n_10168;
wire n_14350;
wire n_8722;
wire n_3467;
wire n_5821;
wire n_11664;
wire n_3179;
wire n_6622;
wire n_12187;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_7665;
wire n_5262;
wire n_7677;
wire n_13169;
wire n_3262;
wire n_10366;
wire n_5319;
wire n_10287;
wire n_14017;
wire n_13940;
wire n_7469;
wire n_3699;
wire n_10163;
wire n_6118;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_14145;
wire n_11006;
wire n_6532;
wire n_13406;
wire n_10431;
wire n_8622;
wire n_3816;
wire n_8099;
wire n_8729;
wire n_9479;
wire n_10876;
wire n_11485;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_9480;
wire n_12453;
wire n_12593;
wire n_4207;
wire n_11449;
wire n_8085;
wire n_4725;
wire n_2757;
wire n_9597;
wire n_10614;
wire n_10786;
wire n_13873;
wire n_13335;
wire n_14273;
wire n_9173;
wire n_10352;
wire n_7203;
wire n_8947;
wire n_9641;
wire n_13714;
wire n_7797;
wire n_9983;
wire n_9267;
wire n_14565;
wire n_5943;
wire n_6556;
wire n_10039;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_13070;
wire n_6216;
wire n_13866;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_7128;
wire n_9849;
wire n_11831;
wire n_5335;
wire n_6365;
wire n_8459;
wire n_7111;
wire n_2801;
wire n_11096;
wire n_4334;
wire n_8478;
wire n_5284;
wire n_12288;
wire n_8786;
wire n_9414;
wire n_4978;
wire n_11677;
wire n_13025;
wire n_14256;
wire n_5771;
wire n_3246;
wire n_9419;
wire n_3299;
wire n_8887;
wire n_12091;
wire n_3623;
wire n_2718;
wire n_11898;
wire n_4707;
wire n_2687;
wire n_8851;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_8540;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_8276;
wire n_7057;
wire n_13457;
wire n_9823;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_9152;
wire n_8706;
wire n_3200;
wire n_6167;
wire n_12357;
wire n_3642;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_11826;
wire n_12629;
wire n_8532;
wire n_9533;
wire n_10750;
wire n_5433;
wire n_3682;
wire n_11825;
wire n_5429;
wire n_7278;
wire n_12893;
wire n_9281;
wire n_9103;
wire n_9111;
wire n_6772;
wire n_7088;
wire n_7799;
wire n_9618;
wire n_10383;
wire n_5698;
wire n_10856;
wire n_5731;
wire n_14532;
wire n_14105;
wire n_10883;
wire n_12935;
wire n_8871;
wire n_4007;
wire n_8433;
wire n_9065;
wire n_10429;
wire n_14627;
wire n_14463;
wire n_6159;
wire n_5857;
wire n_7048;
wire n_12732;
wire n_7979;
wire n_12569;
wire n_9674;
wire n_6617;
wire n_7725;
wire n_13547;
wire n_10859;
wire n_5120;
wire n_3572;
wire n_8371;
wire n_2975;
wire n_8547;
wire n_11538;
wire n_10815;
wire n_11008;
wire n_4075;
wire n_3471;
wire n_8467;
wire n_12980;
wire n_11093;
wire n_11585;
wire n_2932;
wire n_8409;
wire n_6217;
wire n_3118;
wire n_10303;
wire n_9157;
wire n_11616;
wire n_5560;
wire n_9170;
wire n_4441;
wire n_10424;
wire n_3039;
wire n_5455;
wire n_3922;
wire n_6777;
wire n_8640;
wire n_11001;
wire n_10196;
wire n_6742;
wire n_7447;
wire n_5209;
wire n_10684;
wire n_13154;
wire n_6307;
wire n_5704;
wire n_14129;
wire n_4458;
wire n_4889;
wire n_8431;
wire n_14547;
wire n_3831;
wire n_4523;
wire n_13280;
wire n_3618;
wire n_5916;
wire n_8415;
wire n_10184;
wire n_3705;
wire n_3022;
wire n_13904;
wire n_10421;
wire n_13944;
wire n_13359;
wire n_6479;
wire n_11472;
wire n_14376;
wire n_13855;
wire n_13073;
wire n_5099;
wire n_11063;
wire n_3286;
wire n_5781;
wire n_11179;
wire n_5619;
wire n_9416;
wire n_11885;
wire n_3974;
wire n_9368;
wire n_7365;
wire n_3443;
wire n_8329;
wire n_13083;
wire n_14201;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_5022;
wire n_8089;
wire n_9208;
wire n_11657;
wire n_6370;
wire n_9223;
wire n_13124;
wire n_13771;
wire n_10329;
wire n_10924;
wire n_13845;
wire n_11921;
wire n_3996;
wire n_3761;
wire n_14224;
wire n_10285;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_12099;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_9781;
wire n_3009;
wire n_13609;
wire n_13572;
wire n_13817;
wire n_8633;
wire n_12897;
wire n_7095;
wire n_7390;
wire n_9392;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_9422;
wire n_8541;
wire n_10084;
wire n_12924;
wire n_8762;
wire n_14162;
wire n_12619;
wire n_12541;
wire n_3951;
wire n_5518;
wire n_9970;
wire n_3035;
wire n_13428;
wire n_4261;
wire n_7037;
wire n_13104;
wire n_9338;
wire n_11647;
wire n_8125;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_10077;
wire n_3942;
wire n_3023;
wire n_10964;
wire n_14367;
wire n_9492;
wire n_3290;
wire n_14566;
wire n_6693;
wire n_10759;
wire n_9226;
wire n_6712;
wire n_7530;
wire n_10129;
wire n_10101;
wire n_3957;
wire n_13844;
wire n_11757;
wire n_3418;
wire n_10566;
wire n_7471;
wire n_9328;
wire n_6465;
wire n_8188;
wire n_10192;
wire n_5673;
wire n_14363;
wire n_11846;
wire n_11519;
wire n_14571;
wire n_8615;
wire n_5814;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_8011;
wire n_12191;
wire n_10207;
wire n_6730;
wire n_11530;
wire n_13526;
wire n_13998;
wire n_6367;
wire n_8923;
wire n_11488;
wire n_3326;
wire n_11389;
wire n_8624;
wire n_8222;
wire n_11928;
wire n_12429;
wire n_12825;
wire n_6069;
wire n_2732;
wire n_6515;
wire n_8206;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_9513;
wire n_11315;
wire n_3224;
wire n_9393;
wire n_13267;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_13506;
wire n_8065;
wire n_9914;
wire n_14398;
wire n_2949;
wire n_7008;
wire n_12318;
wire n_12918;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_7540;
wire n_10886;
wire n_12923;
wire n_13632;
wire n_14600;
wire n_10804;
wire n_7581;
wire n_12077;
wire n_10362;
wire n_7139;
wire n_10384;
wire n_10437;
wire n_13834;
wire n_8935;
wire n_14213;
wire n_13444;
wire n_10885;
wire n_11962;
wire n_11002;
wire n_3803;
wire n_14331;
wire n_5239;
wire n_2994;
wire n_13885;
wire n_12805;
wire n_7782;
wire n_7432;
wire n_4913;
wire n_13067;
wire n_8155;
wire n_9334;
wire n_14059;
wire n_11648;
wire n_10093;
wire n_13924;
wire n_14289;
wire n_4428;
wire n_12808;
wire n_6483;
wire n_7770;
wire n_12853;
wire n_9684;
wire n_12591;
wire n_8397;
wire n_8568;
wire n_4463;
wire n_10600;
wire n_10480;
wire n_11994;
wire n_5357;
wire n_8175;
wire n_7173;
wire n_3648;
wire n_10892;
wire n_9254;
wire n_6810;
wire n_6576;
wire n_10003;
wire n_10796;
wire n_5421;
wire n_9083;
wire n_11250;
wire n_11050;
wire n_11316;
wire n_14485;
wire n_12987;
wire n_4396;
wire n_13717;
wire n_6708;
wire n_12251;
wire n_10252;
wire n_12948;
wire n_8026;
wire n_6667;
wire n_9175;
wire n_9838;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_11428;
wire n_12467;
wire n_12756;
wire n_2623;
wire n_11463;
wire n_6040;
wire n_10495;
wire n_6847;
wire n_8974;
wire n_6305;
wire n_8836;
wire n_10812;
wire n_4034;
wire n_12678;
wire n_14211;
wire n_4228;
wire n_14641;
wire n_12700;
wire n_11674;
wire n_11097;
wire n_11069;
wire n_7251;
wire n_10894;
wire n_3166;
wire n_12602;
wire n_14155;
wire n_12194;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_8168;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_11318;
wire n_7751;
wire n_12351;
wire n_7951;
wire n_12965;
wire n_7060;
wire n_14184;
wire n_3924;
wire n_9336;
wire n_3997;
wire n_12367;
wire n_13603;
wire n_8873;
wire n_14111;
wire n_10311;
wire n_7591;
wire n_10490;
wire n_3564;
wire n_5769;
wire n_2637;
wire n_6750;
wire n_7444;
wire n_10702;
wire n_7911;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_7790;
wire n_11586;
wire n_7426;
wire n_11786;
wire n_13571;
wire n_4400;
wire n_3953;
wire n_7502;
wire n_13492;
wire n_2959;
wire n_5434;
wire n_10906;
wire n_6855;
wire n_10840;
wire n_10891;
wire n_8170;
wire n_14257;
wire n_5181;
wire n_6239;
wire n_10181;
wire n_3208;
wire n_13673;
wire n_12036;
wire n_9554;
wire n_14589;
wire n_5768;
wire n_11330;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_8120;
wire n_12263;
wire n_9116;
wire n_9315;
wire n_9830;
wire n_8825;
wire n_14416;
wire n_9169;
wire n_2916;
wire n_7252;
wire n_11201;
wire n_5963;
wire n_9999;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_12703;
wire n_4192;
wire n_8003;
wire n_11979;
wire n_12253;
wire n_9215;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_8395;
wire n_13986;
wire n_7065;
wire n_8083;
wire n_11888;
wire n_6177;
wire n_14596;
wire n_8057;
wire n_2581;
wire n_5937;
wire n_9259;
wire n_5146;
wire n_7367;
wire n_10755;
wire n_14274;
wire n_11835;
wire n_11537;
wire n_8164;
wire n_10525;
wire n_11583;
wire n_12776;
wire n_7405;
wire n_7267;
wire n_4646;
wire n_4221;
wire n_12445;
wire n_3650;
wire n_8877;
wire n_6825;
wire n_7614;
wire n_6460;
wire n_4035;
wire n_9150;
wire n_6952;
wire n_9595;
wire n_3670;
wire n_11420;
wire n_8366;
wire n_6173;
wire n_4190;
wire n_8476;
wire n_11527;
wire n_3060;
wire n_6218;
wire n_10342;
wire n_10435;
wire n_11048;
wire n_7685;
wire n_14584;
wire n_11933;
wire n_6486;
wire n_13826;
wire n_4009;
wire n_2984;
wire n_11900;
wire n_12620;
wire n_7619;
wire n_11106;
wire n_12299;
wire n_13078;
wire n_5013;
wire n_4145;
wire n_10983;
wire n_11266;
wire n_6852;
wire n_11340;
wire n_11929;
wire n_5577;
wire n_12673;
wire n_13516;
wire n_9100;
wire n_5872;
wire n_7883;
wire n_13557;
wire n_10397;
wire n_6692;
wire n_13208;
wire n_9707;
wire n_5017;
wire n_8854;
wire n_13523;
wire n_12834;
wire n_10202;
wire n_14549;
wire n_12821;
wire n_10677;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_10648;
wire n_9262;
wire n_5976;
wire n_4717;
wire n_9249;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_11964;
wire n_12247;
wire n_13030;
wire n_8256;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_13065;
wire n_7270;
wire n_10273;
wire n_12927;
wire n_12324;
wire n_12817;
wire n_11255;
wire n_8621;
wire n_13753;
wire n_11751;
wire n_4750;
wire n_10978;
wire n_9806;
wire n_10834;
wire n_13430;
wire n_8577;
wire n_9019;
wire n_10097;
wire n_13880;
wire n_2725;
wire n_2667;
wire n_9361;
wire n_3746;
wire n_7731;
wire n_6626;
wire n_13175;
wire n_4537;
wire n_13050;
wire n_10890;
wire n_5838;
wire n_13732;
wire n_7034;
wire n_10816;
wire n_8654;
wire n_3694;
wire n_12887;
wire n_13133;
wire n_6854;
wire n_7940;
wire n_6793;
wire n_14188;
wire n_5456;
wire n_4847;
wire n_3893;
wire n_5846;
wire n_9814;
wire n_11930;
wire n_3702;
wire n_5930;
wire n_11269;
wire n_10462;
wire n_12316;
wire n_12539;
wire n_13358;
wire n_8952;
wire n_13823;
wire n_12758;
wire n_12414;
wire n_3453;
wire n_9438;
wire n_7537;
wire n_12600;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_11985;
wire n_4427;
wire n_7458;
wire n_7740;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_12949;
wire n_2945;
wire n_3543;
wire n_9856;
wire n_8421;
wire n_11205;
wire n_7179;
wire n_10832;
wire n_3448;
wire n_7433;
wire n_13499;
wire n_4279;
wire n_14057;
wire n_9327;
wire n_9313;
wire n_4330;
wire n_2936;
wire n_6334;
wire n_3609;
wire n_13560;
wire n_6257;
wire n_10142;
wire n_4152;
wire n_6874;
wire n_14073;
wire n_14079;
wire n_10300;
wire n_8911;
wire n_5537;
wire n_9518;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_10335;
wire n_2570;
wire n_2789;
wire n_5409;
wire n_10753;
wire n_14220;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_12783;
wire n_13658;
wire n_5142;
wire n_12431;
wire n_10921;
wire n_10177;
wire n_8971;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_10567;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_11915;
wire n_7987;
wire n_9291;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_9009;
wire n_9882;
wire n_6377;
wire n_10492;
wire n_14137;
wire n_12061;
wire n_5401;
wire n_4595;
wire n_7272;
wire n_11873;
wire n_8215;
wire n_5201;
wire n_5816;
wire n_12628;
wire n_5551;
wire n_9722;
wire n_5416;
wire n_14175;
wire n_4404;
wire n_14644;
wire n_7906;
wire n_2652;
wire n_11260;
wire n_5498;
wire n_5543;
wire n_12359;
wire n_4054;
wire n_9760;
wire n_6018;
wire n_7765;
wire n_14320;
wire n_6021;
wire n_11880;
wire n_11605;
wire n_13615;
wire n_4617;
wire n_14022;
wire n_12974;
wire n_13156;
wire n_10741;
wire n_4611;
wire n_10037;
wire n_8949;
wire n_3169;
wire n_12136;
wire n_5797;
wire n_9454;
wire n_10760;
wire n_6511;
wire n_13849;
wire n_12121;
wire n_7815;
wire n_12658;
wire n_11838;
wire n_13956;
wire n_4732;
wire n_10607;
wire n_5942;
wire n_5764;
wire n_13702;
wire n_8983;
wire n_4969;
wire n_11089;
wire n_14314;
wire n_8121;
wire n_5252;
wire n_11629;
wire n_11259;
wire n_5777;
wire n_11100;
wire n_13119;
wire n_8942;
wire n_7785;
wire n_11608;
wire n_13756;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_12364;
wire n_14628;
wire n_13867;
wire n_8280;
wire n_7728;
wire n_2607;
wire n_11632;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_7181;
wire n_12156;
wire n_11443;
wire n_2796;
wire n_13409;
wire n_13832;
wire n_5393;
wire n_10658;
wire n_8328;
wire n_4817;
wire n_8861;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_8427;
wire n_11161;
wire n_11770;
wire n_13509;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_14399;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2947;
wire n_5643;
wire n_11466;
wire n_10489;
wire n_9826;
wire n_9937;
wire n_10347;
wire n_12632;
wire n_3769;
wire n_11810;
wire n_7825;
wire n_13168;
wire n_4437;
wire n_6419;
wire n_7916;
wire n_13581;
wire n_10952;
wire n_3055;
wire n_8194;
wire n_10758;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_9453;
wire n_7903;
wire n_9900;
wire n_12033;
wire n_7089;
wire n_8217;
wire n_14534;
wire n_10518;
wire n_9331;
wire n_7604;
wire n_2635;
wire n_11789;
wire n_7647;
wire n_2999;
wire n_12465;
wire n_13447;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_14164;
wire n_5868;
wire n_6417;
wire n_8285;
wire n_8521;
wire n_7145;
wire n_10808;
wire n_12358;
wire n_4867;
wire n_3667;
wire n_12446;
wire n_9178;
wire n_7803;
wire n_9689;
wire n_13999;
wire n_2713;
wire n_8448;
wire n_14526;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_11690;
wire n_5986;
wire n_12684;
wire n_9355;
wire n_12851;
wire n_13725;
wire n_9489;
wire n_13319;
wire n_6932;
wire n_12307;
wire n_10971;
wire n_2934;
wire n_7258;
wire n_13019;
wire n_5104;
wire n_12341;
wire n_13807;
wire n_6961;
wire n_8732;
wire n_13297;
wire n_7622;
wire n_14610;
wire n_11968;
wire n_9359;
wire n_13395;
wire n_7839;
wire n_11854;
wire n_6792;
wire n_7720;
wire n_4368;
wire n_5794;
wire n_8136;
wire n_10404;
wire n_3141;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_11797;
wire n_8420;
wire n_13672;
wire n_4430;
wire n_8386;
wire n_6123;
wire n_3238;
wire n_5338;
wire n_7440;
wire n_10802;
wire n_9568;
wire n_6831;
wire n_4544;
wire n_3175;
wire n_14302;
wire n_2666;
wire n_5578;
wire n_12654;
wire n_4191;
wire n_4409;
wire n_12921;
wire n_11991;
wire n_7809;
wire n_3255;
wire n_10340;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_14170;
wire n_7072;
wire n_10681;
wire n_14303;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_11618;
wire n_3509;
wire n_11502;
wire n_10452;
wire n_10221;
wire n_8746;
wire n_10051;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_12498;
wire n_3770;
wire n_6458;
wire n_11465;
wire n_12768;
wire n_9401;
wire n_8857;
wire n_11335;
wire n_6986;
wire n_9495;
wire n_3456;
wire n_12625;
wire n_13221;
wire n_10987;
wire n_4532;
wire n_10551;
wire n_7564;
wire n_12063;
wire n_10396;
wire n_10646;
wire n_13471;
wire n_13021;
wire n_10955;
wire n_5863;
wire n_8185;
wire n_8313;
wire n_6633;
wire n_11382;
wire n_13062;
wire n_3790;
wire n_14298;
wire n_7775;
wire n_7118;
wire n_9234;
wire n_13706;
wire n_7960;
wire n_6152;
wire n_9431;
wire n_5734;
wire n_10308;
wire n_10023;
wire n_8281;
wire n_12347;
wire n_12543;
wire n_2566;
wire n_12958;
wire n_11254;
wire n_5095;
wire n_3101;
wire n_10538;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_12532;
wire n_7069;
wire n_11388;
wire n_5199;
wire n_13347;
wire n_6546;
wire n_14051;
wire n_4257;
wire n_4282;
wire n_11043;
wire n_7636;
wire n_4341;
wire n_10199;
wire n_6925;
wire n_10673;
wire n_7186;
wire n_10467;
wire n_8766;
wire n_13976;
wire n_4027;
wire n_12334;
wire n_4650;
wire n_4309;
wire n_5480;
wire n_6428;
wire n_6924;
wire n_12876;
wire n_3077;
wire n_4944;
wire n_8066;
wire n_11252;
wire n_9340;
wire n_12774;
wire n_12544;
wire n_13793;
wire n_9380;
wire n_7666;
wire n_12653;
wire n_6425;
wire n_12353;
wire n_11824;
wire n_10581;
wire n_14594;
wire n_3478;
wire n_14369;
wire n_3062;
wire n_10818;
wire n_9976;
wire n_4994;
wire n_10226;
wire n_7967;
wire n_5977;
wire n_14515;
wire n_8314;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_11724;
wire n_3978;
wire n_12052;
wire n_11507;
wire n_3836;
wire n_11086;
wire n_10647;
wire n_13184;
wire n_9064;
wire n_3409;
wire n_4381;
wire n_8239;
wire n_9092;
wire n_3583;
wire n_11533;
wire n_4316;
wire n_7301;
wire n_11905;
wire n_14160;
wire n_4860;
wire n_4469;
wire n_9746;
wire n_12994;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_8497;
wire n_10637;
wire n_7262;
wire n_5959;
wire n_13856;
wire n_8056;
wire n_8210;
wire n_3563;
wire n_10769;
wire n_5945;
wire n_4423;
wire n_3310;
wire n_2642;
wire n_12215;
wire n_10519;
wire n_3689;
wire n_13218;
wire n_7584;
wire n_7748;
wire n_9066;
wire n_14637;
wire n_6301;
wire n_13298;
wire n_5668;
wire n_12535;
wire n_3442;
wire n_3972;
wire n_14248;
wire n_4209;
wire n_12582;
wire n_4703;
wire n_6282;
wire n_7686;
wire n_4934;
wire n_11800;
wire n_9870;
wire n_14391;
wire n_9817;
wire n_2638;
wire n_12505;
wire n_13396;
wire n_13988;
wire n_14648;
wire n_7059;
wire n_6985;
wire n_4350;
wire n_5600;
wire n_13132;
wire n_6737;
wire n_10723;
wire n_12875;
wire n_9857;
wire n_13794;
wire n_4804;
wire n_8404;
wire n_4888;
wire n_5767;
wire n_9455;
wire n_10056;
wire n_6459;
wire n_7670;
wire n_13400;
wire n_2977;
wire n_3991;
wire n_13813;
wire n_14307;
wire n_4936;
wire n_8505;
wire n_10653;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_9916;
wire n_10157;
wire n_2600;
wire n_8606;
wire n_13542;
wire n_7443;
wire n_10701;
wire n_10470;
wire n_10923;
wire n_12828;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_12402;
wire n_14387;
wire n_3806;
wire n_9440;
wire n_4759;
wire n_10038;
wire n_9059;
wire n_11691;
wire n_9812;
wire n_14666;
wire n_5869;
wire n_5914;
wire n_6753;
wire n_9690;
wire n_13879;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_11594;
wire n_9912;
wire n_11687;
wire n_4887;
wire n_3751;
wire n_9002;
wire n_11513;
wire n_3402;
wire n_9620;
wire n_10619;
wire n_13522;
wire n_6448;
wire n_9229;
wire n_12524;
wire n_14535;
wire n_5186;
wire n_14196;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_13403;
wire n_10454;
wire n_11655;
wire n_3406;
wire n_13241;
wire n_3664;
wire n_4218;
wire n_9464;
wire n_11386;
wire n_4687;
wire n_7077;
wire n_14060;
wire n_10656;
wire n_10871;
wire n_3686;
wire n_8518;
wire n_11111;
wire n_4720;
wire n_2889;
wire n_13270;
wire n_11938;
wire n_6043;
wire n_6268;
wire n_12670;
wire n_9497;
wire n_14543;
wire n_5604;
wire n_3470;
wire n_7663;
wire n_8350;
wire n_8741;
wire n_10444;
wire n_5221;
wire n_7024;
wire n_8148;
wire n_11833;
wire n_8408;
wire n_6145;
wire n_11866;
wire n_12308;
wire n_2865;
wire n_10846;
wire n_12659;
wire n_13934;
wire n_13024;
wire n_5925;
wire n_6529;
wire n_5591;
wire n_4762;
wire n_13223;
wire n_3844;
wire n_3259;
wire n_8236;
wire n_14202;
wire n_11192;
wire n_11229;
wire n_7214;
wire n_11244;
wire n_8806;
wire n_14352;
wire n_2572;
wire n_4490;
wire n_8295;
wire n_9587;
wire n_3677;
wire n_13888;
wire n_7977;
wire n_5387;
wire n_13529;
wire n_12452;
wire n_3292;
wire n_6311;
wire n_8167;
wire n_11848;
wire n_8377;
wire n_13530;
wire n_3989;
wire n_7652;
wire n_13591;
wire n_10558;
wire n_9783;
wire n_4644;
wire n_8956;
wire n_4752;
wire n_8673;
wire n_4746;
wire n_7566;
wire n_14631;
wire n_4131;
wire n_11876;
wire n_12667;
wire n_5449;
wire n_8760;
wire n_4215;
wire n_12707;
wire n_6134;
wire n_4158;
wire n_6812;
wire n_10466;
wire n_3079;
wire n_10044;
wire n_10546;
wire n_12878;
wire n_5190;
wire n_6733;
wire n_11666;
wire n_3269;
wire n_5325;
wire n_13354;
wire n_10527;
wire n_4231;
wire n_8960;
wire n_9008;
wire n_8957;
wire n_10143;
wire n_12361;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_10233;
wire n_6262;
wire n_4926;
wire n_8207;
wire n_6938;
wire n_4872;
wire n_12709;
wire n_4778;
wire n_5876;
wire n_10461;
wire n_5344;
wire n_3177;
wire n_6160;
wire n_10186;
wire n_4667;
wire n_5813;
wire n_10113;
wire n_12721;
wire n_6235;
wire n_13023;
wire n_6212;
wire n_3440;
wire n_9381;
wire n_9194;
wire n_6816;
wire n_8904;
wire n_3658;
wire n_12264;
wire n_14683;
wire n_7374;
wire n_12464;
wire n_13268;
wire n_12753;
wire n_3404;
wire n_13887;
wire n_3346;
wire n_2816;
wire n_12968;
wire n_10120;
wire n_5892;
wire n_9549;
wire n_7678;
wire n_4837;
wire n_4210;
wire n_11248;
wire n_13660;
wire n_7110;
wire n_5714;
wire n_12111;
wire n_6953;
wire n_9652;
wire n_7975;
wire n_9957;
wire n_13481;
wire n_12609;
wire n_13143;
wire n_12482;
wire n_8451;
wire n_6089;
wire n_10591;
wire n_11780;
wire n_5634;
wire n_12966;
wire n_5133;
wire n_14607;
wire n_7553;
wire n_8527;
wire n_5305;
wire n_5990;
wire n_7732;
wire n_5689;
wire n_7086;
wire n_7891;
wire n_13383;
wire n_13419;
wire n_9089;
wire n_4578;
wire n_8840;
wire n_11424;
wire n_11467;
wire n_5644;
wire n_9137;
wire n_9390;
wire n_3644;
wire n_11995;
wire n_12178;
wire n_8038;
wire n_8190;
wire n_9439;
wire n_11701;
wire n_3059;
wire n_6138;
wire n_9080;
wire n_13351;
wire n_9296;
wire n_12997;
wire n_10625;
wire n_13544;
wire n_4877;
wire n_14173;
wire n_9312;
wire n_10662;
wire n_12818;
wire n_9151;
wire n_8179;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_9883;
wire n_13420;
wire n_14576;
wire n_8287;
wire n_10697;
wire n_8341;
wire n_8111;
wire n_13527;
wire n_8830;
wire n_13206;
wire n_13235;
wire n_4998;
wire n_10200;
wire n_14436;
wire n_5576;
wire n_13399;
wire n_2868;
wire n_10935;
wire n_7345;
wire n_9324;
wire n_13317;
wire n_9631;
wire n_8308;
wire n_10547;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_8021;
wire n_11092;
wire n_13622;
wire n_10933;
wire n_2724;
wire n_8965;
wire n_9736;
wire n_7041;
wire n_9365;
wire n_10632;
wire n_6717;
wire n_14651;
wire n_7593;
wire n_8265;
wire n_13564;
wire n_11166;
wire n_6881;
wire n_10085;
wire n_3328;
wire n_9600;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_9816;
wire n_5343;
wire n_6672;
wire n_9869;
wire n_7757;
wire n_8251;
wire n_9402;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_13276;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_8773;
wire n_12195;
wire n_14383;
wire n_14400;
wire n_5947;
wire n_6242;
wire n_14143;
wire n_6601;
wire n_8570;
wire n_12536;
wire n_10645;
wire n_3469;
wire n_10041;
wire n_12168;
wire n_2835;
wire n_5835;
wire n_10096;
wire n_12533;
wire n_8579;
wire n_3743;
wire n_8079;
wire n_5542;
wire n_9615;
wire n_11869;
wire n_14106;
wire n_2948;
wire n_5015;
wire n_13792;
wire n_3099;
wire n_12560;
wire n_5527;
wire n_2897;
wire n_9711;
wire n_9759;
wire n_4812;
wire n_8506;
wire n_8973;
wire n_13171;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_13764;
wire n_8291;
wire n_3155;
wire n_4300;
wire n_11264;
wire n_10336;
wire n_9820;
wire n_8320;
wire n_7758;
wire n_8635;
wire n_12477;
wire n_9703;
wire n_4472;
wire n_12516;
wire n_9819;
wire n_9118;
wire n_11060;
wire n_2699;
wire n_9321;
wire n_12523;
wire n_11493;
wire n_11562;
wire n_13698;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_10703;
wire n_8375;
wire n_11575;
wire n_2973;
wire n_10449;
wire n_13462;
wire n_10280;
wire n_9428;
wire n_8612;
wire n_10198;
wire n_8778;
wire n_11065;
wire n_5893;
wire n_9292;
wire n_11452;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_12486;
wire n_6462;
wire n_11345;
wire n_4519;
wire n_9018;
wire n_13741;
wire n_5025;
wire n_8872;
wire n_12743;
wire n_10371;
wire n_7333;
wire n_3878;
wire n_12297;
wire n_4197;
wire n_12246;
wire n_13440;
wire n_6669;
wire n_8006;
wire n_11495;
wire n_9565;
wire n_2721;
wire n_13325;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_8491;
wire n_8218;
wire n_13089;
wire n_13578;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_5726;
wire n_3933;
wire n_7439;
wire n_4371;
wire n_12610;
wire n_14006;
wire n_10483;
wire n_12771;
wire n_5828;
wire n_7744;
wire n_2784;
wire n_7210;
wire n_10346;
wire n_3898;
wire n_11864;
wire n_6228;
wire n_10805;
wire n_14107;
wire n_6702;
wire n_7358;
wire n_8240;
wire n_10059;
wire n_9961;
wire n_4749;
wire n_12763;
wire n_7707;
wire n_5924;
wire n_7733;
wire n_13496;
wire n_14536;
wire n_5545;
wire n_8458;
wire n_8853;
wire n_9603;
wire n_11293;
wire n_5083;
wire n_7684;
wire n_10700;
wire n_11984;
wire n_3253;
wire n_11961;
wire n_8306;
wire n_11981;
wire n_14599;
wire n_6997;
wire n_9692;
wire n_4238;
wire n_6371;
wire n_13222;
wire n_11559;
wire n_7673;
wire n_14642;
wire n_12172;
wire n_11942;
wire n_11207;
wire n_11686;
wire n_12280;
wire n_12883;
wire n_7187;
wire n_8013;
wire n_14476;
wire n_3824;
wire n_8342;
wire n_10502;
wire n_12064;
wire n_12480;
wire n_7313;
wire n_10974;
wire n_5899;
wire n_11239;
wire n_14221;
wire n_10250;
wire n_10511;
wire n_9012;
wire n_11482;
wire n_3846;
wire n_12682;
wire n_10831;
wire n_5122;
wire n_11992;
wire n_4189;
wire n_2705;
wire n_12621;
wire n_4479;
wire n_13754;
wire n_10613;
wire n_6641;
wire n_3845;
wire n_12283;
wire n_6463;
wire n_10172;
wire n_3203;
wire n_10351;
wire n_13285;
wire n_4986;
wire n_10333;
wire n_4668;
wire n_9868;
wire n_6264;
wire n_5782;
wire n_8119;
wire n_9264;
wire n_4168;
wire n_8582;
wire n_11479;
wire n_7036;
wire n_11814;
wire n_4298;
wire n_10594;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_13181;
wire n_11622;
wire n_8445;
wire n_12225;
wire n_9720;
wire n_4250;
wire n_13004;
wire n_11067;
wire n_3143;
wire n_8044;
wire n_13413;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_8363;
wire n_8464;
wire n_8921;
wire n_12208;
wire n_14072;
wire n_13608;
wire n_12126;
wire n_13397;
wire n_11083;
wire n_14282;
wire n_10010;
wire n_10588;
wire n_11907;
wire n_12396;
wire n_12984;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_9646;
wire n_11952;
wire n_7480;
wire n_13997;
wire n_12158;
wire n_8843;
wire n_13513;
wire n_5185;
wire n_8405;
wire n_13232;
wire n_2964;
wire n_13296;
wire n_13816;
wire n_8376;
wire n_13859;
wire n_5032;
wire n_11506;
wire n_6990;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_10797;
wire n_8694;
wire n_2913;
wire n_8848;
wire n_6288;
wire n_13989;
wire n_14573;
wire n_3752;
wire n_8752;
wire n_10643;
wire n_3672;
wire n_8894;
wire n_8625;
wire n_7380;
wire n_14058;
wire n_2839;
wire n_8813;
wire n_3237;
wire n_7708;
wire n_12690;
wire n_12813;
wire n_11524;
wire n_10905;
wire n_9842;
wire n_11859;
wire n_4128;
wire n_11228;
wire n_12725;
wire n_4036;
wire n_9671;
wire n_5269;
wire n_8430;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_11035;
wire n_10784;
wire n_4807;
wire n_11023;
wire n_8770;
wire n_6277;
wire n_8426;
wire n_14009;
wire n_5115;
wire n_12474;
wire n_7376;
wire n_11174;
wire n_8411;
wire n_13759;
wire n_8817;
wire n_8461;
wire n_10438;
wire n_3918;
wire n_10234;
wire n_10946;
wire n_11582;
wire n_9230;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_4383;
wire n_4830;
wire n_11705;
wire n_4391;
wire n_11796;
wire n_12484;
wire n_9893;
wire n_6409;
wire n_4095;
wire n_8391;
wire n_8507;
wire n_12021;
wire n_5927;
wire n_8691;
wire n_9188;
wire n_11003;
wire n_4485;
wire n_9032;
wire n_7657;
wire n_6388;
wire n_10275;
wire n_3593;
wire n_6839;
wire n_14284;
wire n_5163;
wire n_9614;
wire n_8967;
wire n_12990;
wire n_2582;
wire n_4356;
wire n_3327;
wire n_9628;
wire n_9231;
wire n_10854;
wire n_6864;
wire n_14309;
wire n_13652;
wire n_13207;
wire n_4890;
wire n_10204;
wire n_8084;
wire n_8856;
wire n_12778;
wire n_12685;
wire n_6679;
wire n_12862;
wire n_11528;
wire n_10734;
wire n_13442;
wire n_10201;
wire n_8631;
wire n_6051;
wire n_4224;
wire n_2563;
wire n_8219;
wire n_9730;
wire n_5507;
wire n_10608;
wire n_4573;
wire n_10746;
wire n_4943;
wire n_2875;
wire n_10676;
wire n_6599;
wire n_3519;
wire n_14423;
wire n_12177;
wire n_13128;
wire n_7504;
wire n_14086;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_5642;
wire n_12672;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_8428;
wire n_9172;
wire n_12141;
wire n_14665;
wire n_14342;
wire n_9926;
wire n_14634;
wire n_6738;
wire n_12665;
wire n_13719;
wire n_5226;
wire n_11615;
wire n_11079;
wire n_8338;
wire n_7602;
wire n_9180;
wire n_9017;
wire n_12024;
wire n_12795;
wire n_9269;
wire n_6566;
wire n_9026;
wire n_13453;
wire n_9462;
wire n_10900;
wire n_5696;
wire n_7998;
wire n_13370;
wire n_8666;
wire n_5014;
wire n_3053;
wire n_7106;
wire n_6346;
wire n_11438;
wire n_11700;
wire n_7557;
wire n_3772;
wire n_7408;
wire n_12940;
wire n_12555;
wire n_14539;
wire n_2891;
wire n_7026;
wire n_4335;
wire n_3128;
wire n_10052;
wire n_13656;
wire n_11668;
wire n_6146;
wire n_13667;
wire n_5677;
wire n_13641;
wire n_4277;
wire n_12487;
wire n_4614;
wire n_4629;
wire n_7394;
wire n_11387;
wire n_9515;
wire n_10560;
wire n_9502;
wire n_13103;
wire n_4516;
wire n_5235;
wire n_13183;
wire n_13720;
wire n_13971;
wire n_11099;
wire n_7627;
wire n_6436;
wire n_12305;
wire n_7719;
wire n_2798;
wire n_10773;
wire n_7450;
wire n_9316;
wire n_3217;
wire n_11996;
wire n_8938;
wire n_6081;
wire n_13436;
wire n_14479;
wire n_10455;
wire n_14410;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_12526;
wire n_3201;
wire n_12622;
wire n_7462;
wire n_12456;
wire n_7780;
wire n_3503;
wire n_8523;
wire n_10391;
wire n_12857;
wire n_5979;
wire n_10476;
wire n_10630;
wire n_10559;
wire n_13797;
wire n_6027;
wire n_13321;
wire n_10911;
wire n_11547;
wire n_10121;
wire n_11064;
wire n_12439;
wire n_4467;
wire n_13809;
wire n_7582;
wire n_10540;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_13575;
wire n_11104;
wire n_9873;
wire n_10473;
wire n_12287;
wire n_10828;
wire n_12182;
wire n_13390;
wire n_8924;
wire n_2965;
wire n_12366;
wire n_4955;
wire n_7555;
wire n_11112;
wire n_10114;
wire n_5410;
wire n_2689;
wire n_6110;
wire n_12552;
wire n_14123;
wire n_10269;
wire n_14258;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_8380;
wire n_13371;
wire n_12777;
wire n_9978;
wire n_5241;
wire n_12492;
wire n_10418;
wire n_4248;
wire n_4645;
wire n_13231;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_3204;
wire n_10672;
wire n_7451;
wire n_9494;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_14601;
wire n_11850;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_12437;
wire n_6612;
wire n_10922;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_1536),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_763),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_1080),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_1864),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_1645),
.Y(n_2559)
);

CKINVDCx5p33_ASAP7_75t_R g2560 ( 
.A(n_1143),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_1528),
.Y(n_2561)
);

CKINVDCx5p33_ASAP7_75t_R g2562 ( 
.A(n_2013),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2469),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_2275),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_1746),
.Y(n_2565)
);

BUFx2_ASAP7_75t_L g2566 ( 
.A(n_2058),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2044),
.Y(n_2567)
);

BUFx10_ASAP7_75t_L g2568 ( 
.A(n_1161),
.Y(n_2568)
);

INVx2_ASAP7_75t_SL g2569 ( 
.A(n_882),
.Y(n_2569)
);

CKINVDCx5p33_ASAP7_75t_R g2570 ( 
.A(n_519),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_2504),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2323),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_1501),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_132),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_170),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_1144),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_701),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2203),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_781),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_311),
.Y(n_2580)
);

CKINVDCx5p33_ASAP7_75t_R g2581 ( 
.A(n_1607),
.Y(n_2581)
);

INVx1_ASAP7_75t_SL g2582 ( 
.A(n_440),
.Y(n_2582)
);

CKINVDCx20_ASAP7_75t_R g2583 ( 
.A(n_1289),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2400),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_1626),
.Y(n_2585)
);

CKINVDCx20_ASAP7_75t_R g2586 ( 
.A(n_1080),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_1402),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_1156),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_2288),
.Y(n_2589)
);

CKINVDCx20_ASAP7_75t_R g2590 ( 
.A(n_1536),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_829),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_843),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_1651),
.Y(n_2593)
);

CKINVDCx20_ASAP7_75t_R g2594 ( 
.A(n_1191),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_1973),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_486),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2422),
.Y(n_2597)
);

BUFx3_ASAP7_75t_L g2598 ( 
.A(n_2270),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_255),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_66),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_306),
.Y(n_2601)
);

CKINVDCx5p33_ASAP7_75t_R g2602 ( 
.A(n_2494),
.Y(n_2602)
);

CKINVDCx5p33_ASAP7_75t_R g2603 ( 
.A(n_2059),
.Y(n_2603)
);

BUFx5_ASAP7_75t_L g2604 ( 
.A(n_2374),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_1957),
.Y(n_2605)
);

BUFx2_ASAP7_75t_L g2606 ( 
.A(n_2042),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2318),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_490),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_1256),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_2011),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2029),
.Y(n_2611)
);

CKINVDCx5p33_ASAP7_75t_R g2612 ( 
.A(n_2033),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_2267),
.Y(n_2613)
);

BUFx5_ASAP7_75t_L g2614 ( 
.A(n_789),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_1228),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2218),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_1002),
.Y(n_2617)
);

BUFx3_ASAP7_75t_L g2618 ( 
.A(n_2342),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_796),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_1561),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_92),
.Y(n_2621)
);

CKINVDCx5p33_ASAP7_75t_R g2622 ( 
.A(n_1853),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_1032),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2415),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_1432),
.Y(n_2625)
);

CKINVDCx20_ASAP7_75t_R g2626 ( 
.A(n_1355),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_1394),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_893),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_634),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_385),
.Y(n_2630)
);

CKINVDCx5p33_ASAP7_75t_R g2631 ( 
.A(n_283),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_384),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_2549),
.Y(n_2633)
);

BUFx10_ASAP7_75t_L g2634 ( 
.A(n_1487),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_1179),
.Y(n_2635)
);

CKINVDCx5p33_ASAP7_75t_R g2636 ( 
.A(n_1571),
.Y(n_2636)
);

CKINVDCx5p33_ASAP7_75t_R g2637 ( 
.A(n_2221),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_1219),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_671),
.Y(n_2639)
);

CKINVDCx5p33_ASAP7_75t_R g2640 ( 
.A(n_584),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2472),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_1681),
.Y(n_2642)
);

CKINVDCx5p33_ASAP7_75t_R g2643 ( 
.A(n_1483),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_1009),
.Y(n_2644)
);

CKINVDCx5p33_ASAP7_75t_R g2645 ( 
.A(n_2304),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_2018),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_390),
.Y(n_2647)
);

CKINVDCx20_ASAP7_75t_R g2648 ( 
.A(n_286),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_210),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_557),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2190),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_1522),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_714),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_1470),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_532),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_2340),
.Y(n_2656)
);

BUFx10_ASAP7_75t_L g2657 ( 
.A(n_2435),
.Y(n_2657)
);

CKINVDCx20_ASAP7_75t_R g2658 ( 
.A(n_1089),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_518),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_887),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_1461),
.Y(n_2661)
);

INVx1_ASAP7_75t_SL g2662 ( 
.A(n_1221),
.Y(n_2662)
);

CKINVDCx20_ASAP7_75t_R g2663 ( 
.A(n_840),
.Y(n_2663)
);

CKINVDCx5p33_ASAP7_75t_R g2664 ( 
.A(n_1173),
.Y(n_2664)
);

CKINVDCx5p33_ASAP7_75t_R g2665 ( 
.A(n_1949),
.Y(n_2665)
);

CKINVDCx5p33_ASAP7_75t_R g2666 ( 
.A(n_14),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_1029),
.Y(n_2667)
);

CKINVDCx20_ASAP7_75t_R g2668 ( 
.A(n_639),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_20),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_1530),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_18),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_1261),
.Y(n_2672)
);

CKINVDCx5p33_ASAP7_75t_R g2673 ( 
.A(n_250),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_2002),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_1020),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_1878),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2440),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2295),
.Y(n_2678)
);

CKINVDCx20_ASAP7_75t_R g2679 ( 
.A(n_2369),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_375),
.Y(n_2680)
);

CKINVDCx5p33_ASAP7_75t_R g2681 ( 
.A(n_836),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_662),
.Y(n_2682)
);

INVx1_ASAP7_75t_SL g2683 ( 
.A(n_179),
.Y(n_2683)
);

CKINVDCx20_ASAP7_75t_R g2684 ( 
.A(n_431),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_1138),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_195),
.Y(n_2686)
);

CKINVDCx20_ASAP7_75t_R g2687 ( 
.A(n_2534),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_716),
.Y(n_2688)
);

CKINVDCx5p33_ASAP7_75t_R g2689 ( 
.A(n_878),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2301),
.Y(n_2690)
);

CKINVDCx5p33_ASAP7_75t_R g2691 ( 
.A(n_2309),
.Y(n_2691)
);

CKINVDCx5p33_ASAP7_75t_R g2692 ( 
.A(n_2387),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_440),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2281),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_373),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2170),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_1566),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_1738),
.Y(n_2698)
);

CKINVDCx5p33_ASAP7_75t_R g2699 ( 
.A(n_528),
.Y(n_2699)
);

BUFx6f_ASAP7_75t_L g2700 ( 
.A(n_1663),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_541),
.Y(n_2701)
);

BUFx6f_ASAP7_75t_L g2702 ( 
.A(n_2237),
.Y(n_2702)
);

CKINVDCx5p33_ASAP7_75t_R g2703 ( 
.A(n_226),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_1898),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2354),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_1326),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_685),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_632),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_1061),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_1810),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_1598),
.Y(n_2711)
);

BUFx6f_ASAP7_75t_L g2712 ( 
.A(n_1903),
.Y(n_2712)
);

BUFx3_ASAP7_75t_L g2713 ( 
.A(n_1095),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_257),
.Y(n_2714)
);

CKINVDCx5p33_ASAP7_75t_R g2715 ( 
.A(n_2389),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2409),
.Y(n_2716)
);

CKINVDCx5p33_ASAP7_75t_R g2717 ( 
.A(n_1631),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_208),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_166),
.Y(n_2719)
);

BUFx2_ASAP7_75t_L g2720 ( 
.A(n_1962),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_504),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_2551),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2357),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_587),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_1084),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_2308),
.Y(n_2726)
);

CKINVDCx20_ASAP7_75t_R g2727 ( 
.A(n_37),
.Y(n_2727)
);

CKINVDCx5p33_ASAP7_75t_R g2728 ( 
.A(n_790),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_240),
.Y(n_2729)
);

BUFx10_ASAP7_75t_L g2730 ( 
.A(n_1125),
.Y(n_2730)
);

BUFx6f_ASAP7_75t_L g2731 ( 
.A(n_2493),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_179),
.Y(n_2732)
);

INVx1_ASAP7_75t_SL g2733 ( 
.A(n_2192),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2522),
.Y(n_2734)
);

INVx1_ASAP7_75t_SL g2735 ( 
.A(n_1647),
.Y(n_2735)
);

CKINVDCx5p33_ASAP7_75t_R g2736 ( 
.A(n_1615),
.Y(n_2736)
);

BUFx6f_ASAP7_75t_L g2737 ( 
.A(n_465),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2292),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2099),
.Y(n_2739)
);

CKINVDCx20_ASAP7_75t_R g2740 ( 
.A(n_570),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_510),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2379),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_701),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_1802),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_193),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_873),
.Y(n_2746)
);

CKINVDCx20_ASAP7_75t_R g2747 ( 
.A(n_1656),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_1553),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_114),
.Y(n_2749)
);

BUFx2_ASAP7_75t_L g2750 ( 
.A(n_472),
.Y(n_2750)
);

INVx1_ASAP7_75t_SL g2751 ( 
.A(n_2267),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_1399),
.Y(n_2752)
);

INVx1_ASAP7_75t_SL g2753 ( 
.A(n_2348),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_2355),
.Y(n_2754)
);

CKINVDCx5p33_ASAP7_75t_R g2755 ( 
.A(n_1018),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_1453),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2204),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_994),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_153),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2360),
.Y(n_2760)
);

BUFx6f_ASAP7_75t_L g2761 ( 
.A(n_1249),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_1984),
.Y(n_2762)
);

BUFx10_ASAP7_75t_L g2763 ( 
.A(n_1605),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2160),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_53),
.Y(n_2765)
);

CKINVDCx5p33_ASAP7_75t_R g2766 ( 
.A(n_2367),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2466),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2176),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_282),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_2200),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_412),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_2275),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_401),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_1353),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_1481),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_549),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_894),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_1120),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_1786),
.Y(n_2779)
);

CKINVDCx5p33_ASAP7_75t_R g2780 ( 
.A(n_2373),
.Y(n_2780)
);

BUFx5_ASAP7_75t_L g2781 ( 
.A(n_1218),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_2503),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_1760),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_1955),
.Y(n_2784)
);

CKINVDCx5p33_ASAP7_75t_R g2785 ( 
.A(n_47),
.Y(n_2785)
);

CKINVDCx5p33_ASAP7_75t_R g2786 ( 
.A(n_767),
.Y(n_2786)
);

CKINVDCx5p33_ASAP7_75t_R g2787 ( 
.A(n_428),
.Y(n_2787)
);

CKINVDCx5p33_ASAP7_75t_R g2788 ( 
.A(n_484),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_1376),
.Y(n_2789)
);

CKINVDCx5p33_ASAP7_75t_R g2790 ( 
.A(n_1877),
.Y(n_2790)
);

BUFx6f_ASAP7_75t_L g2791 ( 
.A(n_205),
.Y(n_2791)
);

INVxp67_ASAP7_75t_L g2792 ( 
.A(n_2123),
.Y(n_2792)
);

CKINVDCx20_ASAP7_75t_R g2793 ( 
.A(n_1148),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_1800),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_995),
.Y(n_2795)
);

CKINVDCx5p33_ASAP7_75t_R g2796 ( 
.A(n_296),
.Y(n_2796)
);

CKINVDCx5p33_ASAP7_75t_R g2797 ( 
.A(n_1420),
.Y(n_2797)
);

INVx2_ASAP7_75t_SL g2798 ( 
.A(n_492),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2400),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_212),
.Y(n_2800)
);

CKINVDCx5p33_ASAP7_75t_R g2801 ( 
.A(n_2210),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_1938),
.Y(n_2802)
);

CKINVDCx5p33_ASAP7_75t_R g2803 ( 
.A(n_411),
.Y(n_2803)
);

CKINVDCx5p33_ASAP7_75t_R g2804 ( 
.A(n_274),
.Y(n_2804)
);

INVx2_ASAP7_75t_SL g2805 ( 
.A(n_2540),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_497),
.Y(n_2806)
);

CKINVDCx5p33_ASAP7_75t_R g2807 ( 
.A(n_2352),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_854),
.Y(n_2808)
);

CKINVDCx5p33_ASAP7_75t_R g2809 ( 
.A(n_1151),
.Y(n_2809)
);

CKINVDCx20_ASAP7_75t_R g2810 ( 
.A(n_2350),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_1267),
.Y(n_2811)
);

CKINVDCx5p33_ASAP7_75t_R g2812 ( 
.A(n_2332),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_1232),
.Y(n_2813)
);

CKINVDCx5p33_ASAP7_75t_R g2814 ( 
.A(n_939),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2274),
.Y(n_2815)
);

BUFx2_ASAP7_75t_L g2816 ( 
.A(n_143),
.Y(n_2816)
);

CKINVDCx5p33_ASAP7_75t_R g2817 ( 
.A(n_182),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2368),
.Y(n_2818)
);

BUFx3_ASAP7_75t_L g2819 ( 
.A(n_711),
.Y(n_2819)
);

CKINVDCx5p33_ASAP7_75t_R g2820 ( 
.A(n_2266),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_1392),
.Y(n_2821)
);

CKINVDCx5p33_ASAP7_75t_R g2822 ( 
.A(n_152),
.Y(n_2822)
);

BUFx10_ASAP7_75t_L g2823 ( 
.A(n_2356),
.Y(n_2823)
);

CKINVDCx5p33_ASAP7_75t_R g2824 ( 
.A(n_914),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_1588),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_1756),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_1027),
.Y(n_2827)
);

CKINVDCx5p33_ASAP7_75t_R g2828 ( 
.A(n_2333),
.Y(n_2828)
);

CKINVDCx5p33_ASAP7_75t_R g2829 ( 
.A(n_1813),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_755),
.Y(n_2830)
);

CKINVDCx5p33_ASAP7_75t_R g2831 ( 
.A(n_1911),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_2025),
.Y(n_2832)
);

CKINVDCx5p33_ASAP7_75t_R g2833 ( 
.A(n_1386),
.Y(n_2833)
);

CKINVDCx5p33_ASAP7_75t_R g2834 ( 
.A(n_1085),
.Y(n_2834)
);

BUFx2_ASAP7_75t_L g2835 ( 
.A(n_1222),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2196),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2341),
.Y(n_2837)
);

CKINVDCx5p33_ASAP7_75t_R g2838 ( 
.A(n_345),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_0),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_949),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2324),
.Y(n_2841)
);

CKINVDCx5p33_ASAP7_75t_R g2842 ( 
.A(n_1666),
.Y(n_2842)
);

CKINVDCx5p33_ASAP7_75t_R g2843 ( 
.A(n_2203),
.Y(n_2843)
);

CKINVDCx5p33_ASAP7_75t_R g2844 ( 
.A(n_2168),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_1908),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_1414),
.Y(n_2846)
);

CKINVDCx5p33_ASAP7_75t_R g2847 ( 
.A(n_2327),
.Y(n_2847)
);

CKINVDCx5p33_ASAP7_75t_R g2848 ( 
.A(n_1256),
.Y(n_2848)
);

CKINVDCx5p33_ASAP7_75t_R g2849 ( 
.A(n_2313),
.Y(n_2849)
);

BUFx2_ASAP7_75t_SL g2850 ( 
.A(n_1584),
.Y(n_2850)
);

CKINVDCx5p33_ASAP7_75t_R g2851 ( 
.A(n_1067),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2315),
.Y(n_2852)
);

CKINVDCx20_ASAP7_75t_R g2853 ( 
.A(n_1764),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2405),
.Y(n_2854)
);

CKINVDCx20_ASAP7_75t_R g2855 ( 
.A(n_2399),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_1374),
.Y(n_2856)
);

CKINVDCx5p33_ASAP7_75t_R g2857 ( 
.A(n_2175),
.Y(n_2857)
);

CKINVDCx5p33_ASAP7_75t_R g2858 ( 
.A(n_588),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_1555),
.Y(n_2859)
);

CKINVDCx5p33_ASAP7_75t_R g2860 ( 
.A(n_1124),
.Y(n_2860)
);

CKINVDCx20_ASAP7_75t_R g2861 ( 
.A(n_820),
.Y(n_2861)
);

CKINVDCx5p33_ASAP7_75t_R g2862 ( 
.A(n_1051),
.Y(n_2862)
);

BUFx3_ASAP7_75t_L g2863 ( 
.A(n_2048),
.Y(n_2863)
);

CKINVDCx5p33_ASAP7_75t_R g2864 ( 
.A(n_1630),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_1814),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_1069),
.Y(n_2866)
);

CKINVDCx5p33_ASAP7_75t_R g2867 ( 
.A(n_2282),
.Y(n_2867)
);

CKINVDCx5p33_ASAP7_75t_R g2868 ( 
.A(n_1880),
.Y(n_2868)
);

CKINVDCx5p33_ASAP7_75t_R g2869 ( 
.A(n_1591),
.Y(n_2869)
);

INVxp33_ASAP7_75t_SL g2870 ( 
.A(n_1341),
.Y(n_2870)
);

BUFx3_ASAP7_75t_L g2871 ( 
.A(n_45),
.Y(n_2871)
);

CKINVDCx5p33_ASAP7_75t_R g2872 ( 
.A(n_1521),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2351),
.Y(n_2873)
);

CKINVDCx5p33_ASAP7_75t_R g2874 ( 
.A(n_15),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2272),
.Y(n_2875)
);

CKINVDCx5p33_ASAP7_75t_R g2876 ( 
.A(n_22),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_636),
.Y(n_2877)
);

CKINVDCx5p33_ASAP7_75t_R g2878 ( 
.A(n_65),
.Y(n_2878)
);

CKINVDCx5p33_ASAP7_75t_R g2879 ( 
.A(n_2226),
.Y(n_2879)
);

BUFx10_ASAP7_75t_L g2880 ( 
.A(n_855),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_167),
.Y(n_2881)
);

CKINVDCx20_ASAP7_75t_R g2882 ( 
.A(n_1078),
.Y(n_2882)
);

CKINVDCx5p33_ASAP7_75t_R g2883 ( 
.A(n_840),
.Y(n_2883)
);

CKINVDCx5p33_ASAP7_75t_R g2884 ( 
.A(n_2386),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_530),
.Y(n_2885)
);

CKINVDCx5p33_ASAP7_75t_R g2886 ( 
.A(n_796),
.Y(n_2886)
);

CKINVDCx5p33_ASAP7_75t_R g2887 ( 
.A(n_1158),
.Y(n_2887)
);

CKINVDCx5p33_ASAP7_75t_R g2888 ( 
.A(n_2394),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_644),
.Y(n_2889)
);

INVx2_ASAP7_75t_SL g2890 ( 
.A(n_1283),
.Y(n_2890)
);

CKINVDCx5p33_ASAP7_75t_R g2891 ( 
.A(n_1186),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_1426),
.Y(n_2892)
);

CKINVDCx5p33_ASAP7_75t_R g2893 ( 
.A(n_1367),
.Y(n_2893)
);

CKINVDCx5p33_ASAP7_75t_R g2894 ( 
.A(n_2133),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_321),
.Y(n_2895)
);

CKINVDCx5p33_ASAP7_75t_R g2896 ( 
.A(n_1648),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_885),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_1572),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_430),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_894),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_193),
.Y(n_2901)
);

CKINVDCx5p33_ASAP7_75t_R g2902 ( 
.A(n_419),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2246),
.Y(n_2903)
);

INVx2_ASAP7_75t_SL g2904 ( 
.A(n_1516),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_1166),
.Y(n_2905)
);

CKINVDCx5p33_ASAP7_75t_R g2906 ( 
.A(n_1620),
.Y(n_2906)
);

CKINVDCx5p33_ASAP7_75t_R g2907 ( 
.A(n_777),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_1178),
.Y(n_2908)
);

CKINVDCx5p33_ASAP7_75t_R g2909 ( 
.A(n_2272),
.Y(n_2909)
);

CKINVDCx5p33_ASAP7_75t_R g2910 ( 
.A(n_411),
.Y(n_2910)
);

CKINVDCx5p33_ASAP7_75t_R g2911 ( 
.A(n_2529),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2297),
.Y(n_2912)
);

CKINVDCx5p33_ASAP7_75t_R g2913 ( 
.A(n_1905),
.Y(n_2913)
);

CKINVDCx5p33_ASAP7_75t_R g2914 ( 
.A(n_1362),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_1276),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2320),
.Y(n_2916)
);

CKINVDCx5p33_ASAP7_75t_R g2917 ( 
.A(n_1130),
.Y(n_2917)
);

BUFx2_ASAP7_75t_L g2918 ( 
.A(n_395),
.Y(n_2918)
);

HB1xp67_ASAP7_75t_L g2919 ( 
.A(n_2338),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_499),
.Y(n_2920)
);

INVx2_ASAP7_75t_SL g2921 ( 
.A(n_1268),
.Y(n_2921)
);

CKINVDCx5p33_ASAP7_75t_R g2922 ( 
.A(n_1269),
.Y(n_2922)
);

CKINVDCx14_ASAP7_75t_R g2923 ( 
.A(n_45),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_1089),
.Y(n_2924)
);

CKINVDCx5p33_ASAP7_75t_R g2925 ( 
.A(n_1452),
.Y(n_2925)
);

BUFx6f_ASAP7_75t_L g2926 ( 
.A(n_227),
.Y(n_2926)
);

CKINVDCx5p33_ASAP7_75t_R g2927 ( 
.A(n_1543),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2302),
.Y(n_2928)
);

CKINVDCx5p33_ASAP7_75t_R g2929 ( 
.A(n_729),
.Y(n_2929)
);

CKINVDCx20_ASAP7_75t_R g2930 ( 
.A(n_784),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_836),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_480),
.Y(n_2932)
);

CKINVDCx5p33_ASAP7_75t_R g2933 ( 
.A(n_182),
.Y(n_2933)
);

CKINVDCx5p33_ASAP7_75t_R g2934 ( 
.A(n_1195),
.Y(n_2934)
);

CKINVDCx5p33_ASAP7_75t_R g2935 ( 
.A(n_1195),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_1714),
.Y(n_2936)
);

CKINVDCx5p33_ASAP7_75t_R g2937 ( 
.A(n_1547),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_259),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2267),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_233),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_528),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_2542),
.Y(n_2942)
);

CKINVDCx5p33_ASAP7_75t_R g2943 ( 
.A(n_1407),
.Y(n_2943)
);

CKINVDCx5p33_ASAP7_75t_R g2944 ( 
.A(n_210),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_1503),
.Y(n_2945)
);

HB1xp67_ASAP7_75t_L g2946 ( 
.A(n_460),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_591),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_1399),
.Y(n_2948)
);

INVxp33_ASAP7_75t_SL g2949 ( 
.A(n_1413),
.Y(n_2949)
);

CKINVDCx5p33_ASAP7_75t_R g2950 ( 
.A(n_839),
.Y(n_2950)
);

CKINVDCx20_ASAP7_75t_R g2951 ( 
.A(n_905),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2076),
.Y(n_2952)
);

INVx2_ASAP7_75t_SL g2953 ( 
.A(n_1161),
.Y(n_2953)
);

BUFx10_ASAP7_75t_L g2954 ( 
.A(n_1750),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_114),
.Y(n_2955)
);

CKINVDCx20_ASAP7_75t_R g2956 ( 
.A(n_2336),
.Y(n_2956)
);

CKINVDCx5p33_ASAP7_75t_R g2957 ( 
.A(n_1274),
.Y(n_2957)
);

CKINVDCx5p33_ASAP7_75t_R g2958 ( 
.A(n_676),
.Y(n_2958)
);

CKINVDCx5p33_ASAP7_75t_R g2959 ( 
.A(n_2183),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_1477),
.Y(n_2960)
);

INVxp67_ASAP7_75t_SL g2961 ( 
.A(n_1840),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2271),
.Y(n_2962)
);

INVx1_ASAP7_75t_SL g2963 ( 
.A(n_230),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2439),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_590),
.Y(n_2965)
);

BUFx3_ASAP7_75t_L g2966 ( 
.A(n_902),
.Y(n_2966)
);

CKINVDCx5p33_ASAP7_75t_R g2967 ( 
.A(n_626),
.Y(n_2967)
);

BUFx3_ASAP7_75t_L g2968 ( 
.A(n_929),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_913),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2365),
.Y(n_2970)
);

CKINVDCx5p33_ASAP7_75t_R g2971 ( 
.A(n_1970),
.Y(n_2971)
);

INVx2_ASAP7_75t_SL g2972 ( 
.A(n_1327),
.Y(n_2972)
);

CKINVDCx5p33_ASAP7_75t_R g2973 ( 
.A(n_2113),
.Y(n_2973)
);

CKINVDCx5p33_ASAP7_75t_R g2974 ( 
.A(n_436),
.Y(n_2974)
);

CKINVDCx5p33_ASAP7_75t_R g2975 ( 
.A(n_346),
.Y(n_2975)
);

CKINVDCx5p33_ASAP7_75t_R g2976 ( 
.A(n_1674),
.Y(n_2976)
);

INVx1_ASAP7_75t_SL g2977 ( 
.A(n_1527),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2212),
.Y(n_2978)
);

BUFx3_ASAP7_75t_L g2979 ( 
.A(n_1268),
.Y(n_2979)
);

CKINVDCx20_ASAP7_75t_R g2980 ( 
.A(n_1517),
.Y(n_2980)
);

INVx1_ASAP7_75t_SL g2981 ( 
.A(n_512),
.Y(n_2981)
);

CKINVDCx5p33_ASAP7_75t_R g2982 ( 
.A(n_18),
.Y(n_2982)
);

INVx1_ASAP7_75t_SL g2983 ( 
.A(n_1169),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_988),
.Y(n_2984)
);

BUFx2_ASAP7_75t_L g2985 ( 
.A(n_714),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_1845),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_1461),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2161),
.Y(n_2988)
);

CKINVDCx5p33_ASAP7_75t_R g2989 ( 
.A(n_1854),
.Y(n_2989)
);

CKINVDCx5p33_ASAP7_75t_R g2990 ( 
.A(n_1780),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_1109),
.Y(n_2991)
);

CKINVDCx5p33_ASAP7_75t_R g2992 ( 
.A(n_614),
.Y(n_2992)
);

CKINVDCx5p33_ASAP7_75t_R g2993 ( 
.A(n_520),
.Y(n_2993)
);

CKINVDCx5p33_ASAP7_75t_R g2994 ( 
.A(n_1737),
.Y(n_2994)
);

CKINVDCx5p33_ASAP7_75t_R g2995 ( 
.A(n_327),
.Y(n_2995)
);

CKINVDCx5p33_ASAP7_75t_R g2996 ( 
.A(n_2241),
.Y(n_2996)
);

CKINVDCx5p33_ASAP7_75t_R g2997 ( 
.A(n_1515),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2499),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2353),
.Y(n_2999)
);

CKINVDCx16_ASAP7_75t_R g3000 ( 
.A(n_1225),
.Y(n_3000)
);

HB1xp67_ASAP7_75t_L g3001 ( 
.A(n_200),
.Y(n_3001)
);

BUFx3_ASAP7_75t_L g3002 ( 
.A(n_2254),
.Y(n_3002)
);

CKINVDCx5p33_ASAP7_75t_R g3003 ( 
.A(n_972),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2469),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_1353),
.Y(n_3005)
);

CKINVDCx5p33_ASAP7_75t_R g3006 ( 
.A(n_332),
.Y(n_3006)
);

CKINVDCx5p33_ASAP7_75t_R g3007 ( 
.A(n_215),
.Y(n_3007)
);

CKINVDCx5p33_ASAP7_75t_R g3008 ( 
.A(n_851),
.Y(n_3008)
);

CKINVDCx5p33_ASAP7_75t_R g3009 ( 
.A(n_927),
.Y(n_3009)
);

INVx2_ASAP7_75t_SL g3010 ( 
.A(n_1684),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_1372),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_1353),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2486),
.Y(n_3013)
);

BUFx3_ASAP7_75t_L g3014 ( 
.A(n_1858),
.Y(n_3014)
);

CKINVDCx5p33_ASAP7_75t_R g3015 ( 
.A(n_2291),
.Y(n_3015)
);

INVx1_ASAP7_75t_SL g3016 ( 
.A(n_2261),
.Y(n_3016)
);

BUFx6f_ASAP7_75t_L g3017 ( 
.A(n_76),
.Y(n_3017)
);

CKINVDCx5p33_ASAP7_75t_R g3018 ( 
.A(n_1032),
.Y(n_3018)
);

CKINVDCx5p33_ASAP7_75t_R g3019 ( 
.A(n_2111),
.Y(n_3019)
);

CKINVDCx5p33_ASAP7_75t_R g3020 ( 
.A(n_838),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_1033),
.Y(n_3021)
);

CKINVDCx5p33_ASAP7_75t_R g3022 ( 
.A(n_1307),
.Y(n_3022)
);

CKINVDCx5p33_ASAP7_75t_R g3023 ( 
.A(n_2541),
.Y(n_3023)
);

CKINVDCx5p33_ASAP7_75t_R g3024 ( 
.A(n_512),
.Y(n_3024)
);

CKINVDCx5p33_ASAP7_75t_R g3025 ( 
.A(n_1817),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_70),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_1147),
.Y(n_3027)
);

CKINVDCx5p33_ASAP7_75t_R g3028 ( 
.A(n_1013),
.Y(n_3028)
);

CKINVDCx16_ASAP7_75t_R g3029 ( 
.A(n_2228),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_434),
.Y(n_3030)
);

CKINVDCx5p33_ASAP7_75t_R g3031 ( 
.A(n_1786),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_778),
.Y(n_3032)
);

CKINVDCx5p33_ASAP7_75t_R g3033 ( 
.A(n_1243),
.Y(n_3033)
);

BUFx3_ASAP7_75t_L g3034 ( 
.A(n_1229),
.Y(n_3034)
);

CKINVDCx5p33_ASAP7_75t_R g3035 ( 
.A(n_959),
.Y(n_3035)
);

CKINVDCx20_ASAP7_75t_R g3036 ( 
.A(n_2347),
.Y(n_3036)
);

CKINVDCx5p33_ASAP7_75t_R g3037 ( 
.A(n_513),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2278),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_1204),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_1192),
.Y(n_3040)
);

CKINVDCx20_ASAP7_75t_R g3041 ( 
.A(n_42),
.Y(n_3041)
);

CKINVDCx5p33_ASAP7_75t_R g3042 ( 
.A(n_1396),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2264),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_425),
.Y(n_3044)
);

CKINVDCx5p33_ASAP7_75t_R g3045 ( 
.A(n_463),
.Y(n_3045)
);

CKINVDCx5p33_ASAP7_75t_R g3046 ( 
.A(n_2409),
.Y(n_3046)
);

CKINVDCx20_ASAP7_75t_R g3047 ( 
.A(n_276),
.Y(n_3047)
);

INVx1_ASAP7_75t_SL g3048 ( 
.A(n_2380),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_593),
.Y(n_3049)
);

CKINVDCx16_ASAP7_75t_R g3050 ( 
.A(n_1331),
.Y(n_3050)
);

CKINVDCx5p33_ASAP7_75t_R g3051 ( 
.A(n_862),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_653),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2299),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2481),
.Y(n_3054)
);

CKINVDCx5p33_ASAP7_75t_R g3055 ( 
.A(n_1202),
.Y(n_3055)
);

HB1xp67_ASAP7_75t_L g3056 ( 
.A(n_2379),
.Y(n_3056)
);

CKINVDCx5p33_ASAP7_75t_R g3057 ( 
.A(n_1311),
.Y(n_3057)
);

INVx1_ASAP7_75t_SL g3058 ( 
.A(n_2366),
.Y(n_3058)
);

CKINVDCx5p33_ASAP7_75t_R g3059 ( 
.A(n_1722),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_364),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_647),
.Y(n_3061)
);

CKINVDCx5p33_ASAP7_75t_R g3062 ( 
.A(n_1052),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2390),
.Y(n_3063)
);

CKINVDCx5p33_ASAP7_75t_R g3064 ( 
.A(n_921),
.Y(n_3064)
);

CKINVDCx5p33_ASAP7_75t_R g3065 ( 
.A(n_1552),
.Y(n_3065)
);

INVx1_ASAP7_75t_SL g3066 ( 
.A(n_2287),
.Y(n_3066)
);

CKINVDCx5p33_ASAP7_75t_R g3067 ( 
.A(n_2066),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_1081),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2409),
.Y(n_3069)
);

CKINVDCx5p33_ASAP7_75t_R g3070 ( 
.A(n_330),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_1265),
.Y(n_3071)
);

CKINVDCx5p33_ASAP7_75t_R g3072 ( 
.A(n_1698),
.Y(n_3072)
);

CKINVDCx20_ASAP7_75t_R g3073 ( 
.A(n_1682),
.Y(n_3073)
);

CKINVDCx5p33_ASAP7_75t_R g3074 ( 
.A(n_178),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_318),
.Y(n_3075)
);

CKINVDCx5p33_ASAP7_75t_R g3076 ( 
.A(n_193),
.Y(n_3076)
);

BUFx6f_ASAP7_75t_L g3077 ( 
.A(n_701),
.Y(n_3077)
);

CKINVDCx5p33_ASAP7_75t_R g3078 ( 
.A(n_855),
.Y(n_3078)
);

CKINVDCx5p33_ASAP7_75t_R g3079 ( 
.A(n_1103),
.Y(n_3079)
);

BUFx6f_ASAP7_75t_L g3080 ( 
.A(n_1751),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2296),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_53),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_13),
.Y(n_3083)
);

BUFx8_ASAP7_75t_SL g3084 ( 
.A(n_1285),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_1472),
.Y(n_3085)
);

CKINVDCx5p33_ASAP7_75t_R g3086 ( 
.A(n_284),
.Y(n_3086)
);

CKINVDCx5p33_ASAP7_75t_R g3087 ( 
.A(n_2010),
.Y(n_3087)
);

CKINVDCx5p33_ASAP7_75t_R g3088 ( 
.A(n_859),
.Y(n_3088)
);

CKINVDCx5p33_ASAP7_75t_R g3089 ( 
.A(n_2250),
.Y(n_3089)
);

CKINVDCx5p33_ASAP7_75t_R g3090 ( 
.A(n_2377),
.Y(n_3090)
);

CKINVDCx5p33_ASAP7_75t_R g3091 ( 
.A(n_573),
.Y(n_3091)
);

CKINVDCx5p33_ASAP7_75t_R g3092 ( 
.A(n_981),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2321),
.Y(n_3093)
);

CKINVDCx5p33_ASAP7_75t_R g3094 ( 
.A(n_1120),
.Y(n_3094)
);

CKINVDCx5p33_ASAP7_75t_R g3095 ( 
.A(n_1287),
.Y(n_3095)
);

CKINVDCx20_ASAP7_75t_R g3096 ( 
.A(n_1357),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2148),
.Y(n_3097)
);

CKINVDCx5p33_ASAP7_75t_R g3098 ( 
.A(n_1807),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_475),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_262),
.Y(n_3100)
);

CKINVDCx16_ASAP7_75t_R g3101 ( 
.A(n_680),
.Y(n_3101)
);

CKINVDCx5p33_ASAP7_75t_R g3102 ( 
.A(n_1528),
.Y(n_3102)
);

CKINVDCx5p33_ASAP7_75t_R g3103 ( 
.A(n_1806),
.Y(n_3103)
);

CKINVDCx5p33_ASAP7_75t_R g3104 ( 
.A(n_2337),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_439),
.Y(n_3105)
);

CKINVDCx5p33_ASAP7_75t_R g3106 ( 
.A(n_1684),
.Y(n_3106)
);

CKINVDCx16_ASAP7_75t_R g3107 ( 
.A(n_325),
.Y(n_3107)
);

CKINVDCx14_ASAP7_75t_R g3108 ( 
.A(n_165),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_214),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_1799),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_771),
.Y(n_3111)
);

CKINVDCx5p33_ASAP7_75t_R g3112 ( 
.A(n_1817),
.Y(n_3112)
);

CKINVDCx5p33_ASAP7_75t_R g3113 ( 
.A(n_2101),
.Y(n_3113)
);

BUFx10_ASAP7_75t_L g3114 ( 
.A(n_2199),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2349),
.Y(n_3115)
);

CKINVDCx5p33_ASAP7_75t_R g3116 ( 
.A(n_1284),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_1051),
.Y(n_3117)
);

HB1xp67_ASAP7_75t_L g3118 ( 
.A(n_2505),
.Y(n_3118)
);

CKINVDCx5p33_ASAP7_75t_R g3119 ( 
.A(n_1031),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_876),
.Y(n_3120)
);

CKINVDCx5p33_ASAP7_75t_R g3121 ( 
.A(n_2197),
.Y(n_3121)
);

CKINVDCx5p33_ASAP7_75t_R g3122 ( 
.A(n_508),
.Y(n_3122)
);

CKINVDCx5p33_ASAP7_75t_R g3123 ( 
.A(n_2385),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_1877),
.Y(n_3124)
);

CKINVDCx5p33_ASAP7_75t_R g3125 ( 
.A(n_2528),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_256),
.Y(n_3126)
);

CKINVDCx5p33_ASAP7_75t_R g3127 ( 
.A(n_1699),
.Y(n_3127)
);

INVxp33_ASAP7_75t_R g3128 ( 
.A(n_730),
.Y(n_3128)
);

CKINVDCx5p33_ASAP7_75t_R g3129 ( 
.A(n_40),
.Y(n_3129)
);

CKINVDCx5p33_ASAP7_75t_R g3130 ( 
.A(n_324),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2075),
.Y(n_3131)
);

CKINVDCx5p33_ASAP7_75t_R g3132 ( 
.A(n_1246),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_1994),
.Y(n_3133)
);

CKINVDCx5p33_ASAP7_75t_R g3134 ( 
.A(n_1478),
.Y(n_3134)
);

BUFx2_ASAP7_75t_SL g3135 ( 
.A(n_1503),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_481),
.Y(n_3136)
);

BUFx3_ASAP7_75t_L g3137 ( 
.A(n_1416),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_187),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_104),
.Y(n_3139)
);

CKINVDCx5p33_ASAP7_75t_R g3140 ( 
.A(n_215),
.Y(n_3140)
);

BUFx10_ASAP7_75t_L g3141 ( 
.A(n_1637),
.Y(n_3141)
);

CKINVDCx5p33_ASAP7_75t_R g3142 ( 
.A(n_1599),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_445),
.Y(n_3143)
);

CKINVDCx5p33_ASAP7_75t_R g3144 ( 
.A(n_2384),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_544),
.Y(n_3145)
);

CKINVDCx5p33_ASAP7_75t_R g3146 ( 
.A(n_2501),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2497),
.Y(n_3147)
);

BUFx10_ASAP7_75t_L g3148 ( 
.A(n_1203),
.Y(n_3148)
);

BUFx2_ASAP7_75t_L g3149 ( 
.A(n_1317),
.Y(n_3149)
);

CKINVDCx5p33_ASAP7_75t_R g3150 ( 
.A(n_2329),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_1081),
.Y(n_3151)
);

CKINVDCx5p33_ASAP7_75t_R g3152 ( 
.A(n_137),
.Y(n_3152)
);

BUFx10_ASAP7_75t_L g3153 ( 
.A(n_805),
.Y(n_3153)
);

BUFx6f_ASAP7_75t_L g3154 ( 
.A(n_767),
.Y(n_3154)
);

CKINVDCx5p33_ASAP7_75t_R g3155 ( 
.A(n_2148),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_734),
.Y(n_3156)
);

CKINVDCx5p33_ASAP7_75t_R g3157 ( 
.A(n_1841),
.Y(n_3157)
);

CKINVDCx5p33_ASAP7_75t_R g3158 ( 
.A(n_1831),
.Y(n_3158)
);

BUFx2_ASAP7_75t_SL g3159 ( 
.A(n_2410),
.Y(n_3159)
);

INVx2_ASAP7_75t_SL g3160 ( 
.A(n_358),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2134),
.Y(n_3161)
);

CKINVDCx5p33_ASAP7_75t_R g3162 ( 
.A(n_350),
.Y(n_3162)
);

CKINVDCx20_ASAP7_75t_R g3163 ( 
.A(n_1194),
.Y(n_3163)
);

INVx3_ASAP7_75t_L g3164 ( 
.A(n_1644),
.Y(n_3164)
);

BUFx3_ASAP7_75t_L g3165 ( 
.A(n_711),
.Y(n_3165)
);

BUFx3_ASAP7_75t_L g3166 ( 
.A(n_163),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_1089),
.Y(n_3167)
);

INVxp67_ASAP7_75t_SL g3168 ( 
.A(n_372),
.Y(n_3168)
);

INVxp67_ASAP7_75t_L g3169 ( 
.A(n_17),
.Y(n_3169)
);

CKINVDCx5p33_ASAP7_75t_R g3170 ( 
.A(n_848),
.Y(n_3170)
);

INVx1_ASAP7_75t_SL g3171 ( 
.A(n_311),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_1415),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_650),
.Y(n_3173)
);

CKINVDCx5p33_ASAP7_75t_R g3174 ( 
.A(n_677),
.Y(n_3174)
);

CKINVDCx5p33_ASAP7_75t_R g3175 ( 
.A(n_2418),
.Y(n_3175)
);

CKINVDCx5p33_ASAP7_75t_R g3176 ( 
.A(n_1306),
.Y(n_3176)
);

CKINVDCx20_ASAP7_75t_R g3177 ( 
.A(n_2022),
.Y(n_3177)
);

CKINVDCx20_ASAP7_75t_R g3178 ( 
.A(n_449),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_1499),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_577),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_1667),
.Y(n_3181)
);

CKINVDCx5p33_ASAP7_75t_R g3182 ( 
.A(n_2334),
.Y(n_3182)
);

CKINVDCx5p33_ASAP7_75t_R g3183 ( 
.A(n_69),
.Y(n_3183)
);

CKINVDCx5p33_ASAP7_75t_R g3184 ( 
.A(n_1574),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_1390),
.Y(n_3185)
);

CKINVDCx5p33_ASAP7_75t_R g3186 ( 
.A(n_347),
.Y(n_3186)
);

CKINVDCx5p33_ASAP7_75t_R g3187 ( 
.A(n_2376),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_774),
.Y(n_3188)
);

CKINVDCx5p33_ASAP7_75t_R g3189 ( 
.A(n_2393),
.Y(n_3189)
);

CKINVDCx5p33_ASAP7_75t_R g3190 ( 
.A(n_2327),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_1294),
.Y(n_3191)
);

CKINVDCx5p33_ASAP7_75t_R g3192 ( 
.A(n_2149),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_333),
.Y(n_3193)
);

CKINVDCx5p33_ASAP7_75t_R g3194 ( 
.A(n_443),
.Y(n_3194)
);

BUFx3_ASAP7_75t_L g3195 ( 
.A(n_867),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_486),
.Y(n_3196)
);

CKINVDCx5p33_ASAP7_75t_R g3197 ( 
.A(n_2170),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_1713),
.Y(n_3198)
);

BUFx2_ASAP7_75t_L g3199 ( 
.A(n_1834),
.Y(n_3199)
);

CKINVDCx5p33_ASAP7_75t_R g3200 ( 
.A(n_1125),
.Y(n_3200)
);

CKINVDCx5p33_ASAP7_75t_R g3201 ( 
.A(n_2228),
.Y(n_3201)
);

CKINVDCx5p33_ASAP7_75t_R g3202 ( 
.A(n_145),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2294),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_1442),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2295),
.Y(n_3205)
);

CKINVDCx5p33_ASAP7_75t_R g3206 ( 
.A(n_1469),
.Y(n_3206)
);

CKINVDCx5p33_ASAP7_75t_R g3207 ( 
.A(n_2475),
.Y(n_3207)
);

CKINVDCx5p33_ASAP7_75t_R g3208 ( 
.A(n_2359),
.Y(n_3208)
);

CKINVDCx5p33_ASAP7_75t_R g3209 ( 
.A(n_1748),
.Y(n_3209)
);

CKINVDCx5p33_ASAP7_75t_R g3210 ( 
.A(n_225),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_904),
.Y(n_3211)
);

CKINVDCx5p33_ASAP7_75t_R g3212 ( 
.A(n_539),
.Y(n_3212)
);

CKINVDCx5p33_ASAP7_75t_R g3213 ( 
.A(n_1237),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2006),
.Y(n_3214)
);

INVx1_ASAP7_75t_SL g3215 ( 
.A(n_644),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2247),
.Y(n_3216)
);

BUFx3_ASAP7_75t_L g3217 ( 
.A(n_685),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2195),
.Y(n_3218)
);

CKINVDCx5p33_ASAP7_75t_R g3219 ( 
.A(n_264),
.Y(n_3219)
);

CKINVDCx5p33_ASAP7_75t_R g3220 ( 
.A(n_1536),
.Y(n_3220)
);

BUFx2_ASAP7_75t_L g3221 ( 
.A(n_2172),
.Y(n_3221)
);

CKINVDCx5p33_ASAP7_75t_R g3222 ( 
.A(n_1122),
.Y(n_3222)
);

CKINVDCx5p33_ASAP7_75t_R g3223 ( 
.A(n_2175),
.Y(n_3223)
);

CKINVDCx5p33_ASAP7_75t_R g3224 ( 
.A(n_624),
.Y(n_3224)
);

CKINVDCx5p33_ASAP7_75t_R g3225 ( 
.A(n_1050),
.Y(n_3225)
);

CKINVDCx5p33_ASAP7_75t_R g3226 ( 
.A(n_2248),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_641),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_1194),
.Y(n_3228)
);

INVx2_ASAP7_75t_SL g3229 ( 
.A(n_1625),
.Y(n_3229)
);

CKINVDCx5p33_ASAP7_75t_R g3230 ( 
.A(n_2029),
.Y(n_3230)
);

CKINVDCx5p33_ASAP7_75t_R g3231 ( 
.A(n_1019),
.Y(n_3231)
);

CKINVDCx5p33_ASAP7_75t_R g3232 ( 
.A(n_2024),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_1699),
.Y(n_3233)
);

CKINVDCx5p33_ASAP7_75t_R g3234 ( 
.A(n_1775),
.Y(n_3234)
);

CKINVDCx20_ASAP7_75t_R g3235 ( 
.A(n_886),
.Y(n_3235)
);

CKINVDCx20_ASAP7_75t_R g3236 ( 
.A(n_431),
.Y(n_3236)
);

BUFx3_ASAP7_75t_L g3237 ( 
.A(n_220),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_577),
.Y(n_3238)
);

CKINVDCx5p33_ASAP7_75t_R g3239 ( 
.A(n_1785),
.Y(n_3239)
);

CKINVDCx5p33_ASAP7_75t_R g3240 ( 
.A(n_899),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_1100),
.Y(n_3241)
);

CKINVDCx5p33_ASAP7_75t_R g3242 ( 
.A(n_1054),
.Y(n_3242)
);

BUFx3_ASAP7_75t_L g3243 ( 
.A(n_1812),
.Y(n_3243)
);

BUFx3_ASAP7_75t_L g3244 ( 
.A(n_2316),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2419),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_1776),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_154),
.Y(n_3247)
);

BUFx5_ASAP7_75t_L g3248 ( 
.A(n_704),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2009),
.Y(n_3249)
);

CKINVDCx5p33_ASAP7_75t_R g3250 ( 
.A(n_1073),
.Y(n_3250)
);

BUFx6f_ASAP7_75t_L g3251 ( 
.A(n_1568),
.Y(n_3251)
);

CKINVDCx5p33_ASAP7_75t_R g3252 ( 
.A(n_1169),
.Y(n_3252)
);

HB1xp67_ASAP7_75t_L g3253 ( 
.A(n_1532),
.Y(n_3253)
);

HB1xp67_ASAP7_75t_L g3254 ( 
.A(n_249),
.Y(n_3254)
);

CKINVDCx5p33_ASAP7_75t_R g3255 ( 
.A(n_2295),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_46),
.Y(n_3256)
);

CKINVDCx20_ASAP7_75t_R g3257 ( 
.A(n_2169),
.Y(n_3257)
);

CKINVDCx5p33_ASAP7_75t_R g3258 ( 
.A(n_666),
.Y(n_3258)
);

CKINVDCx5p33_ASAP7_75t_R g3259 ( 
.A(n_686),
.Y(n_3259)
);

CKINVDCx5p33_ASAP7_75t_R g3260 ( 
.A(n_1719),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_2507),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2330),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_2332),
.Y(n_3263)
);

CKINVDCx5p33_ASAP7_75t_R g3264 ( 
.A(n_663),
.Y(n_3264)
);

CKINVDCx5p33_ASAP7_75t_R g3265 ( 
.A(n_1793),
.Y(n_3265)
);

CKINVDCx5p33_ASAP7_75t_R g3266 ( 
.A(n_1382),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_2305),
.Y(n_3267)
);

CKINVDCx5p33_ASAP7_75t_R g3268 ( 
.A(n_421),
.Y(n_3268)
);

BUFx10_ASAP7_75t_L g3269 ( 
.A(n_2026),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_2265),
.Y(n_3270)
);

CKINVDCx5p33_ASAP7_75t_R g3271 ( 
.A(n_112),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_563),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_1394),
.Y(n_3273)
);

CKINVDCx20_ASAP7_75t_R g3274 ( 
.A(n_561),
.Y(n_3274)
);

CKINVDCx5p33_ASAP7_75t_R g3275 ( 
.A(n_414),
.Y(n_3275)
);

BUFx10_ASAP7_75t_L g3276 ( 
.A(n_2053),
.Y(n_3276)
);

CKINVDCx5p33_ASAP7_75t_R g3277 ( 
.A(n_510),
.Y(n_3277)
);

CKINVDCx5p33_ASAP7_75t_R g3278 ( 
.A(n_2317),
.Y(n_3278)
);

INVxp67_ASAP7_75t_L g3279 ( 
.A(n_2427),
.Y(n_3279)
);

CKINVDCx5p33_ASAP7_75t_R g3280 ( 
.A(n_1575),
.Y(n_3280)
);

BUFx6f_ASAP7_75t_L g3281 ( 
.A(n_2530),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_1365),
.Y(n_3282)
);

BUFx10_ASAP7_75t_L g3283 ( 
.A(n_1500),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_430),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_365),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_362),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_1931),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_831),
.Y(n_3288)
);

CKINVDCx16_ASAP7_75t_R g3289 ( 
.A(n_659),
.Y(n_3289)
);

CKINVDCx20_ASAP7_75t_R g3290 ( 
.A(n_971),
.Y(n_3290)
);

INVx3_ASAP7_75t_L g3291 ( 
.A(n_716),
.Y(n_3291)
);

CKINVDCx5p33_ASAP7_75t_R g3292 ( 
.A(n_2258),
.Y(n_3292)
);

BUFx10_ASAP7_75t_L g3293 ( 
.A(n_1201),
.Y(n_3293)
);

CKINVDCx5p33_ASAP7_75t_R g3294 ( 
.A(n_1052),
.Y(n_3294)
);

CKINVDCx5p33_ASAP7_75t_R g3295 ( 
.A(n_1651),
.Y(n_3295)
);

CKINVDCx5p33_ASAP7_75t_R g3296 ( 
.A(n_2497),
.Y(n_3296)
);

CKINVDCx5p33_ASAP7_75t_R g3297 ( 
.A(n_2041),
.Y(n_3297)
);

CKINVDCx5p33_ASAP7_75t_R g3298 ( 
.A(n_195),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_1686),
.Y(n_3299)
);

BUFx6f_ASAP7_75t_L g3300 ( 
.A(n_2312),
.Y(n_3300)
);

CKINVDCx5p33_ASAP7_75t_R g3301 ( 
.A(n_2054),
.Y(n_3301)
);

CKINVDCx5p33_ASAP7_75t_R g3302 ( 
.A(n_479),
.Y(n_3302)
);

INVx1_ASAP7_75t_SL g3303 ( 
.A(n_1939),
.Y(n_3303)
);

INVx2_ASAP7_75t_SL g3304 ( 
.A(n_179),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_1903),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_84),
.Y(n_3306)
);

BUFx5_ASAP7_75t_L g3307 ( 
.A(n_2512),
.Y(n_3307)
);

CKINVDCx5p33_ASAP7_75t_R g3308 ( 
.A(n_2269),
.Y(n_3308)
);

CKINVDCx5p33_ASAP7_75t_R g3309 ( 
.A(n_615),
.Y(n_3309)
);

INVx3_ASAP7_75t_L g3310 ( 
.A(n_438),
.Y(n_3310)
);

BUFx10_ASAP7_75t_L g3311 ( 
.A(n_988),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_381),
.Y(n_3312)
);

BUFx3_ASAP7_75t_L g3313 ( 
.A(n_2239),
.Y(n_3313)
);

BUFx3_ASAP7_75t_L g3314 ( 
.A(n_22),
.Y(n_3314)
);

BUFx8_ASAP7_75t_SL g3315 ( 
.A(n_2219),
.Y(n_3315)
);

CKINVDCx5p33_ASAP7_75t_R g3316 ( 
.A(n_342),
.Y(n_3316)
);

CKINVDCx5p33_ASAP7_75t_R g3317 ( 
.A(n_1768),
.Y(n_3317)
);

CKINVDCx5p33_ASAP7_75t_R g3318 ( 
.A(n_1362),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_1642),
.Y(n_3319)
);

CKINVDCx5p33_ASAP7_75t_R g3320 ( 
.A(n_1316),
.Y(n_3320)
);

BUFx10_ASAP7_75t_L g3321 ( 
.A(n_782),
.Y(n_3321)
);

CKINVDCx5p33_ASAP7_75t_R g3322 ( 
.A(n_2300),
.Y(n_3322)
);

CKINVDCx5p33_ASAP7_75t_R g3323 ( 
.A(n_652),
.Y(n_3323)
);

CKINVDCx5p33_ASAP7_75t_R g3324 ( 
.A(n_2370),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_1070),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_2554),
.Y(n_3326)
);

CKINVDCx5p33_ASAP7_75t_R g3327 ( 
.A(n_607),
.Y(n_3327)
);

CKINVDCx5p33_ASAP7_75t_R g3328 ( 
.A(n_289),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_344),
.Y(n_3329)
);

CKINVDCx5p33_ASAP7_75t_R g3330 ( 
.A(n_1329),
.Y(n_3330)
);

CKINVDCx5p33_ASAP7_75t_R g3331 ( 
.A(n_709),
.Y(n_3331)
);

CKINVDCx5p33_ASAP7_75t_R g3332 ( 
.A(n_1582),
.Y(n_3332)
);

CKINVDCx5p33_ASAP7_75t_R g3333 ( 
.A(n_1103),
.Y(n_3333)
);

INVx2_ASAP7_75t_SL g3334 ( 
.A(n_1810),
.Y(n_3334)
);

CKINVDCx5p33_ASAP7_75t_R g3335 ( 
.A(n_166),
.Y(n_3335)
);

CKINVDCx5p33_ASAP7_75t_R g3336 ( 
.A(n_2285),
.Y(n_3336)
);

INVxp67_ASAP7_75t_L g3337 ( 
.A(n_1166),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_1233),
.Y(n_3338)
);

CKINVDCx14_ASAP7_75t_R g3339 ( 
.A(n_407),
.Y(n_3339)
);

BUFx3_ASAP7_75t_L g3340 ( 
.A(n_1046),
.Y(n_3340)
);

CKINVDCx5p33_ASAP7_75t_R g3341 ( 
.A(n_2251),
.Y(n_3341)
);

CKINVDCx5p33_ASAP7_75t_R g3342 ( 
.A(n_30),
.Y(n_3342)
);

CKINVDCx5p33_ASAP7_75t_R g3343 ( 
.A(n_1242),
.Y(n_3343)
);

CKINVDCx5p33_ASAP7_75t_R g3344 ( 
.A(n_1144),
.Y(n_3344)
);

CKINVDCx5p33_ASAP7_75t_R g3345 ( 
.A(n_1488),
.Y(n_3345)
);

CKINVDCx5p33_ASAP7_75t_R g3346 ( 
.A(n_789),
.Y(n_3346)
);

CKINVDCx5p33_ASAP7_75t_R g3347 ( 
.A(n_1667),
.Y(n_3347)
);

CKINVDCx5p33_ASAP7_75t_R g3348 ( 
.A(n_1115),
.Y(n_3348)
);

CKINVDCx5p33_ASAP7_75t_R g3349 ( 
.A(n_120),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_1995),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_1417),
.Y(n_3351)
);

INVx3_ASAP7_75t_L g3352 ( 
.A(n_165),
.Y(n_3352)
);

BUFx8_ASAP7_75t_SL g3353 ( 
.A(n_815),
.Y(n_3353)
);

CKINVDCx5p33_ASAP7_75t_R g3354 ( 
.A(n_2298),
.Y(n_3354)
);

HB1xp67_ASAP7_75t_L g3355 ( 
.A(n_434),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2170),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2322),
.Y(n_3357)
);

CKINVDCx5p33_ASAP7_75t_R g3358 ( 
.A(n_2156),
.Y(n_3358)
);

BUFx6f_ASAP7_75t_L g3359 ( 
.A(n_2015),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_2127),
.Y(n_3360)
);

CKINVDCx5p33_ASAP7_75t_R g3361 ( 
.A(n_1572),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_791),
.Y(n_3362)
);

CKINVDCx5p33_ASAP7_75t_R g3363 ( 
.A(n_30),
.Y(n_3363)
);

CKINVDCx5p33_ASAP7_75t_R g3364 ( 
.A(n_449),
.Y(n_3364)
);

CKINVDCx5p33_ASAP7_75t_R g3365 ( 
.A(n_2345),
.Y(n_3365)
);

CKINVDCx5p33_ASAP7_75t_R g3366 ( 
.A(n_2049),
.Y(n_3366)
);

CKINVDCx5p33_ASAP7_75t_R g3367 ( 
.A(n_614),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_661),
.Y(n_3368)
);

CKINVDCx5p33_ASAP7_75t_R g3369 ( 
.A(n_2396),
.Y(n_3369)
);

CKINVDCx5p33_ASAP7_75t_R g3370 ( 
.A(n_2514),
.Y(n_3370)
);

CKINVDCx5p33_ASAP7_75t_R g3371 ( 
.A(n_2163),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_864),
.Y(n_3372)
);

CKINVDCx5p33_ASAP7_75t_R g3373 ( 
.A(n_1770),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_1200),
.Y(n_3374)
);

BUFx3_ASAP7_75t_L g3375 ( 
.A(n_939),
.Y(n_3375)
);

CKINVDCx5p33_ASAP7_75t_R g3376 ( 
.A(n_2136),
.Y(n_3376)
);

CKINVDCx5p33_ASAP7_75t_R g3377 ( 
.A(n_2536),
.Y(n_3377)
);

CKINVDCx16_ASAP7_75t_R g3378 ( 
.A(n_850),
.Y(n_3378)
);

CKINVDCx20_ASAP7_75t_R g3379 ( 
.A(n_2037),
.Y(n_3379)
);

INVx2_ASAP7_75t_SL g3380 ( 
.A(n_1816),
.Y(n_3380)
);

BUFx8_ASAP7_75t_SL g3381 ( 
.A(n_863),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_1623),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2030),
.Y(n_3383)
);

BUFx6f_ASAP7_75t_L g3384 ( 
.A(n_1663),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_1779),
.Y(n_3385)
);

INVxp67_ASAP7_75t_L g3386 ( 
.A(n_660),
.Y(n_3386)
);

CKINVDCx5p33_ASAP7_75t_R g3387 ( 
.A(n_378),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_2164),
.Y(n_3388)
);

CKINVDCx5p33_ASAP7_75t_R g3389 ( 
.A(n_672),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_317),
.Y(n_3390)
);

CKINVDCx5p33_ASAP7_75t_R g3391 ( 
.A(n_329),
.Y(n_3391)
);

BUFx5_ASAP7_75t_L g3392 ( 
.A(n_2276),
.Y(n_3392)
);

CKINVDCx5p33_ASAP7_75t_R g3393 ( 
.A(n_160),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_876),
.Y(n_3394)
);

CKINVDCx5p33_ASAP7_75t_R g3395 ( 
.A(n_75),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_614),
.Y(n_3396)
);

CKINVDCx5p33_ASAP7_75t_R g3397 ( 
.A(n_915),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_1814),
.Y(n_3398)
);

CKINVDCx5p33_ASAP7_75t_R g3399 ( 
.A(n_1579),
.Y(n_3399)
);

CKINVDCx5p33_ASAP7_75t_R g3400 ( 
.A(n_319),
.Y(n_3400)
);

CKINVDCx5p33_ASAP7_75t_R g3401 ( 
.A(n_1893),
.Y(n_3401)
);

INVx2_ASAP7_75t_SL g3402 ( 
.A(n_1336),
.Y(n_3402)
);

CKINVDCx16_ASAP7_75t_R g3403 ( 
.A(n_108),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_2343),
.Y(n_3404)
);

CKINVDCx5p33_ASAP7_75t_R g3405 ( 
.A(n_2264),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_883),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_164),
.Y(n_3407)
);

CKINVDCx5p33_ASAP7_75t_R g3408 ( 
.A(n_1574),
.Y(n_3408)
);

CKINVDCx5p33_ASAP7_75t_R g3409 ( 
.A(n_246),
.Y(n_3409)
);

BUFx5_ASAP7_75t_L g3410 ( 
.A(n_771),
.Y(n_3410)
);

BUFx3_ASAP7_75t_L g3411 ( 
.A(n_877),
.Y(n_3411)
);

CKINVDCx5p33_ASAP7_75t_R g3412 ( 
.A(n_94),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_286),
.Y(n_3413)
);

CKINVDCx5p33_ASAP7_75t_R g3414 ( 
.A(n_1763),
.Y(n_3414)
);

CKINVDCx5p33_ASAP7_75t_R g3415 ( 
.A(n_1313),
.Y(n_3415)
);

CKINVDCx5p33_ASAP7_75t_R g3416 ( 
.A(n_1026),
.Y(n_3416)
);

INVx2_ASAP7_75t_SL g3417 ( 
.A(n_817),
.Y(n_3417)
);

CKINVDCx5p33_ASAP7_75t_R g3418 ( 
.A(n_282),
.Y(n_3418)
);

CKINVDCx20_ASAP7_75t_R g3419 ( 
.A(n_1507),
.Y(n_3419)
);

HB1xp67_ASAP7_75t_L g3420 ( 
.A(n_727),
.Y(n_3420)
);

CKINVDCx5p33_ASAP7_75t_R g3421 ( 
.A(n_2072),
.Y(n_3421)
);

CKINVDCx20_ASAP7_75t_R g3422 ( 
.A(n_2273),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_892),
.Y(n_3423)
);

CKINVDCx5p33_ASAP7_75t_R g3424 ( 
.A(n_980),
.Y(n_3424)
);

CKINVDCx5p33_ASAP7_75t_R g3425 ( 
.A(n_1285),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_2413),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_1472),
.Y(n_3427)
);

INVx1_ASAP7_75t_SL g3428 ( 
.A(n_1573),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2007),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_867),
.Y(n_3430)
);

CKINVDCx5p33_ASAP7_75t_R g3431 ( 
.A(n_824),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_452),
.Y(n_3432)
);

CKINVDCx5p33_ASAP7_75t_R g3433 ( 
.A(n_63),
.Y(n_3433)
);

CKINVDCx5p33_ASAP7_75t_R g3434 ( 
.A(n_2458),
.Y(n_3434)
);

CKINVDCx5p33_ASAP7_75t_R g3435 ( 
.A(n_497),
.Y(n_3435)
);

INVxp67_ASAP7_75t_L g3436 ( 
.A(n_939),
.Y(n_3436)
);

CKINVDCx5p33_ASAP7_75t_R g3437 ( 
.A(n_826),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_1860),
.Y(n_3438)
);

CKINVDCx5p33_ASAP7_75t_R g3439 ( 
.A(n_778),
.Y(n_3439)
);

BUFx2_ASAP7_75t_L g3440 ( 
.A(n_1551),
.Y(n_3440)
);

CKINVDCx16_ASAP7_75t_R g3441 ( 
.A(n_1301),
.Y(n_3441)
);

BUFx6f_ASAP7_75t_L g3442 ( 
.A(n_1505),
.Y(n_3442)
);

CKINVDCx5p33_ASAP7_75t_R g3443 ( 
.A(n_1821),
.Y(n_3443)
);

CKINVDCx20_ASAP7_75t_R g3444 ( 
.A(n_2446),
.Y(n_3444)
);

CKINVDCx5p33_ASAP7_75t_R g3445 ( 
.A(n_1525),
.Y(n_3445)
);

CKINVDCx5p33_ASAP7_75t_R g3446 ( 
.A(n_1098),
.Y(n_3446)
);

CKINVDCx5p33_ASAP7_75t_R g3447 ( 
.A(n_2323),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_2478),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_2489),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_1441),
.Y(n_3450)
);

CKINVDCx5p33_ASAP7_75t_R g3451 ( 
.A(n_1380),
.Y(n_3451)
);

CKINVDCx5p33_ASAP7_75t_R g3452 ( 
.A(n_197),
.Y(n_3452)
);

CKINVDCx5p33_ASAP7_75t_R g3453 ( 
.A(n_1403),
.Y(n_3453)
);

CKINVDCx20_ASAP7_75t_R g3454 ( 
.A(n_2395),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_737),
.Y(n_3455)
);

CKINVDCx20_ASAP7_75t_R g3456 ( 
.A(n_149),
.Y(n_3456)
);

CKINVDCx5p33_ASAP7_75t_R g3457 ( 
.A(n_822),
.Y(n_3457)
);

CKINVDCx5p33_ASAP7_75t_R g3458 ( 
.A(n_2262),
.Y(n_3458)
);

INVx1_ASAP7_75t_SL g3459 ( 
.A(n_243),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_1314),
.Y(n_3460)
);

CKINVDCx5p33_ASAP7_75t_R g3461 ( 
.A(n_478),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2018),
.Y(n_3462)
);

CKINVDCx5p33_ASAP7_75t_R g3463 ( 
.A(n_884),
.Y(n_3463)
);

CKINVDCx20_ASAP7_75t_R g3464 ( 
.A(n_86),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_163),
.Y(n_3465)
);

CKINVDCx5p33_ASAP7_75t_R g3466 ( 
.A(n_2346),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_1965),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_1305),
.Y(n_3468)
);

CKINVDCx5p33_ASAP7_75t_R g3469 ( 
.A(n_350),
.Y(n_3469)
);

CKINVDCx5p33_ASAP7_75t_R g3470 ( 
.A(n_1102),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_1254),
.Y(n_3471)
);

CKINVDCx5p33_ASAP7_75t_R g3472 ( 
.A(n_1878),
.Y(n_3472)
);

CKINVDCx5p33_ASAP7_75t_R g3473 ( 
.A(n_2388),
.Y(n_3473)
);

CKINVDCx5p33_ASAP7_75t_R g3474 ( 
.A(n_377),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_2383),
.Y(n_3475)
);

CKINVDCx5p33_ASAP7_75t_R g3476 ( 
.A(n_301),
.Y(n_3476)
);

CKINVDCx5p33_ASAP7_75t_R g3477 ( 
.A(n_1011),
.Y(n_3477)
);

CKINVDCx5p33_ASAP7_75t_R g3478 ( 
.A(n_1132),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_2362),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_1256),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_2406),
.Y(n_3481)
);

CKINVDCx5p33_ASAP7_75t_R g3482 ( 
.A(n_653),
.Y(n_3482)
);

CKINVDCx5p33_ASAP7_75t_R g3483 ( 
.A(n_2381),
.Y(n_3483)
);

CKINVDCx5p33_ASAP7_75t_R g3484 ( 
.A(n_2454),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_2539),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_52),
.Y(n_3486)
);

CKINVDCx5p33_ASAP7_75t_R g3487 ( 
.A(n_1814),
.Y(n_3487)
);

CKINVDCx5p33_ASAP7_75t_R g3488 ( 
.A(n_609),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_1717),
.Y(n_3489)
);

CKINVDCx5p33_ASAP7_75t_R g3490 ( 
.A(n_2485),
.Y(n_3490)
);

CKINVDCx5p33_ASAP7_75t_R g3491 ( 
.A(n_1119),
.Y(n_3491)
);

CKINVDCx5p33_ASAP7_75t_R g3492 ( 
.A(n_542),
.Y(n_3492)
);

CKINVDCx5p33_ASAP7_75t_R g3493 ( 
.A(n_908),
.Y(n_3493)
);

CKINVDCx5p33_ASAP7_75t_R g3494 ( 
.A(n_1163),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_464),
.Y(n_3495)
);

CKINVDCx5p33_ASAP7_75t_R g3496 ( 
.A(n_1075),
.Y(n_3496)
);

CKINVDCx5p33_ASAP7_75t_R g3497 ( 
.A(n_2479),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_860),
.Y(n_3498)
);

CKINVDCx5p33_ASAP7_75t_R g3499 ( 
.A(n_2526),
.Y(n_3499)
);

CKINVDCx20_ASAP7_75t_R g3500 ( 
.A(n_2183),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_2263),
.Y(n_3501)
);

CKINVDCx5p33_ASAP7_75t_R g3502 ( 
.A(n_159),
.Y(n_3502)
);

INVx4_ASAP7_75t_R g3503 ( 
.A(n_1561),
.Y(n_3503)
);

CKINVDCx5p33_ASAP7_75t_R g3504 ( 
.A(n_1073),
.Y(n_3504)
);

CKINVDCx5p33_ASAP7_75t_R g3505 ( 
.A(n_1088),
.Y(n_3505)
);

CKINVDCx5p33_ASAP7_75t_R g3506 ( 
.A(n_251),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_661),
.Y(n_3507)
);

CKINVDCx5p33_ASAP7_75t_R g3508 ( 
.A(n_911),
.Y(n_3508)
);

CKINVDCx5p33_ASAP7_75t_R g3509 ( 
.A(n_540),
.Y(n_3509)
);

CKINVDCx5p33_ASAP7_75t_R g3510 ( 
.A(n_1826),
.Y(n_3510)
);

CKINVDCx5p33_ASAP7_75t_R g3511 ( 
.A(n_1151),
.Y(n_3511)
);

CKINVDCx5p33_ASAP7_75t_R g3512 ( 
.A(n_1307),
.Y(n_3512)
);

CKINVDCx5p33_ASAP7_75t_R g3513 ( 
.A(n_1778),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_787),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_1363),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_1794),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_1893),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_2378),
.Y(n_3518)
);

CKINVDCx5p33_ASAP7_75t_R g3519 ( 
.A(n_58),
.Y(n_3519)
);

BUFx3_ASAP7_75t_L g3520 ( 
.A(n_2018),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_1844),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_2458),
.Y(n_3522)
);

CKINVDCx5p33_ASAP7_75t_R g3523 ( 
.A(n_1274),
.Y(n_3523)
);

CKINVDCx5p33_ASAP7_75t_R g3524 ( 
.A(n_1558),
.Y(n_3524)
);

CKINVDCx5p33_ASAP7_75t_R g3525 ( 
.A(n_116),
.Y(n_3525)
);

CKINVDCx20_ASAP7_75t_R g3526 ( 
.A(n_251),
.Y(n_3526)
);

CKINVDCx5p33_ASAP7_75t_R g3527 ( 
.A(n_2514),
.Y(n_3527)
);

CKINVDCx5p33_ASAP7_75t_R g3528 ( 
.A(n_1950),
.Y(n_3528)
);

CKINVDCx5p33_ASAP7_75t_R g3529 ( 
.A(n_2414),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_2306),
.Y(n_3530)
);

CKINVDCx5p33_ASAP7_75t_R g3531 ( 
.A(n_551),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_657),
.Y(n_3532)
);

CKINVDCx5p33_ASAP7_75t_R g3533 ( 
.A(n_1157),
.Y(n_3533)
);

CKINVDCx5p33_ASAP7_75t_R g3534 ( 
.A(n_405),
.Y(n_3534)
);

CKINVDCx5p33_ASAP7_75t_R g3535 ( 
.A(n_131),
.Y(n_3535)
);

CKINVDCx5p33_ASAP7_75t_R g3536 ( 
.A(n_22),
.Y(n_3536)
);

BUFx2_ASAP7_75t_L g3537 ( 
.A(n_1778),
.Y(n_3537)
);

INVx1_ASAP7_75t_SL g3538 ( 
.A(n_669),
.Y(n_3538)
);

HB1xp67_ASAP7_75t_L g3539 ( 
.A(n_580),
.Y(n_3539)
);

CKINVDCx5p33_ASAP7_75t_R g3540 ( 
.A(n_495),
.Y(n_3540)
);

BUFx5_ASAP7_75t_L g3541 ( 
.A(n_812),
.Y(n_3541)
);

CKINVDCx5p33_ASAP7_75t_R g3542 ( 
.A(n_89),
.Y(n_3542)
);

CKINVDCx5p33_ASAP7_75t_R g3543 ( 
.A(n_105),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_1772),
.Y(n_3544)
);

BUFx3_ASAP7_75t_L g3545 ( 
.A(n_1478),
.Y(n_3545)
);

CKINVDCx5p33_ASAP7_75t_R g3546 ( 
.A(n_1465),
.Y(n_3546)
);

CKINVDCx5p33_ASAP7_75t_R g3547 ( 
.A(n_1086),
.Y(n_3547)
);

CKINVDCx5p33_ASAP7_75t_R g3548 ( 
.A(n_72),
.Y(n_3548)
);

INVx1_ASAP7_75t_SL g3549 ( 
.A(n_513),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_2397),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_2252),
.Y(n_3551)
);

CKINVDCx5p33_ASAP7_75t_R g3552 ( 
.A(n_1564),
.Y(n_3552)
);

CKINVDCx5p33_ASAP7_75t_R g3553 ( 
.A(n_787),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_1017),
.Y(n_3554)
);

CKINVDCx20_ASAP7_75t_R g3555 ( 
.A(n_186),
.Y(n_3555)
);

CKINVDCx5p33_ASAP7_75t_R g3556 ( 
.A(n_2225),
.Y(n_3556)
);

BUFx3_ASAP7_75t_L g3557 ( 
.A(n_1801),
.Y(n_3557)
);

INVx2_ASAP7_75t_SL g3558 ( 
.A(n_932),
.Y(n_3558)
);

CKINVDCx5p33_ASAP7_75t_R g3559 ( 
.A(n_1447),
.Y(n_3559)
);

CKINVDCx5p33_ASAP7_75t_R g3560 ( 
.A(n_43),
.Y(n_3560)
);

CKINVDCx5p33_ASAP7_75t_R g3561 ( 
.A(n_1559),
.Y(n_3561)
);

INVxp67_ASAP7_75t_L g3562 ( 
.A(n_82),
.Y(n_3562)
);

CKINVDCx5p33_ASAP7_75t_R g3563 ( 
.A(n_888),
.Y(n_3563)
);

CKINVDCx5p33_ASAP7_75t_R g3564 ( 
.A(n_872),
.Y(n_3564)
);

INVx1_ASAP7_75t_SL g3565 ( 
.A(n_1481),
.Y(n_3565)
);

CKINVDCx5p33_ASAP7_75t_R g3566 ( 
.A(n_1754),
.Y(n_3566)
);

CKINVDCx16_ASAP7_75t_R g3567 ( 
.A(n_1275),
.Y(n_3567)
);

HB1xp67_ASAP7_75t_L g3568 ( 
.A(n_547),
.Y(n_3568)
);

CKINVDCx5p33_ASAP7_75t_R g3569 ( 
.A(n_419),
.Y(n_3569)
);

CKINVDCx5p33_ASAP7_75t_R g3570 ( 
.A(n_1396),
.Y(n_3570)
);

CKINVDCx5p33_ASAP7_75t_R g3571 ( 
.A(n_2431),
.Y(n_3571)
);

CKINVDCx5p33_ASAP7_75t_R g3572 ( 
.A(n_1574),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_1283),
.Y(n_3573)
);

CKINVDCx5p33_ASAP7_75t_R g3574 ( 
.A(n_1545),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_284),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_388),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_1280),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_1725),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_892),
.Y(n_3579)
);

BUFx10_ASAP7_75t_L g3580 ( 
.A(n_1553),
.Y(n_3580)
);

CKINVDCx5p33_ASAP7_75t_R g3581 ( 
.A(n_1198),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_110),
.Y(n_3582)
);

CKINVDCx5p33_ASAP7_75t_R g3583 ( 
.A(n_2033),
.Y(n_3583)
);

CKINVDCx5p33_ASAP7_75t_R g3584 ( 
.A(n_119),
.Y(n_3584)
);

CKINVDCx5p33_ASAP7_75t_R g3585 ( 
.A(n_2372),
.Y(n_3585)
);

BUFx2_ASAP7_75t_L g3586 ( 
.A(n_2353),
.Y(n_3586)
);

CKINVDCx5p33_ASAP7_75t_R g3587 ( 
.A(n_173),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_1977),
.Y(n_3588)
);

BUFx6f_ASAP7_75t_L g3589 ( 
.A(n_580),
.Y(n_3589)
);

BUFx2_ASAP7_75t_L g3590 ( 
.A(n_743),
.Y(n_3590)
);

BUFx6f_ASAP7_75t_L g3591 ( 
.A(n_376),
.Y(n_3591)
);

CKINVDCx5p33_ASAP7_75t_R g3592 ( 
.A(n_1266),
.Y(n_3592)
);

CKINVDCx5p33_ASAP7_75t_R g3593 ( 
.A(n_1664),
.Y(n_3593)
);

CKINVDCx5p33_ASAP7_75t_R g3594 ( 
.A(n_131),
.Y(n_3594)
);

CKINVDCx16_ASAP7_75t_R g3595 ( 
.A(n_2356),
.Y(n_3595)
);

INVx1_ASAP7_75t_SL g3596 ( 
.A(n_1644),
.Y(n_3596)
);

CKINVDCx20_ASAP7_75t_R g3597 ( 
.A(n_1699),
.Y(n_3597)
);

CKINVDCx5p33_ASAP7_75t_R g3598 ( 
.A(n_2481),
.Y(n_3598)
);

INVx2_ASAP7_75t_SL g3599 ( 
.A(n_475),
.Y(n_3599)
);

BUFx6f_ASAP7_75t_L g3600 ( 
.A(n_2173),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_1968),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_517),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_181),
.Y(n_3603)
);

CKINVDCx5p33_ASAP7_75t_R g3604 ( 
.A(n_1689),
.Y(n_3604)
);

CKINVDCx5p33_ASAP7_75t_R g3605 ( 
.A(n_240),
.Y(n_3605)
);

CKINVDCx5p33_ASAP7_75t_R g3606 ( 
.A(n_1760),
.Y(n_3606)
);

INVx2_ASAP7_75t_L g3607 ( 
.A(n_622),
.Y(n_3607)
);

CKINVDCx20_ASAP7_75t_R g3608 ( 
.A(n_2010),
.Y(n_3608)
);

CKINVDCx5p33_ASAP7_75t_R g3609 ( 
.A(n_633),
.Y(n_3609)
);

CKINVDCx5p33_ASAP7_75t_R g3610 ( 
.A(n_1937),
.Y(n_3610)
);

CKINVDCx5p33_ASAP7_75t_R g3611 ( 
.A(n_700),
.Y(n_3611)
);

CKINVDCx5p33_ASAP7_75t_R g3612 ( 
.A(n_2014),
.Y(n_3612)
);

CKINVDCx20_ASAP7_75t_R g3613 ( 
.A(n_2413),
.Y(n_3613)
);

CKINVDCx5p33_ASAP7_75t_R g3614 ( 
.A(n_2055),
.Y(n_3614)
);

CKINVDCx5p33_ASAP7_75t_R g3615 ( 
.A(n_1644),
.Y(n_3615)
);

CKINVDCx5p33_ASAP7_75t_R g3616 ( 
.A(n_1334),
.Y(n_3616)
);

INVx1_ASAP7_75t_SL g3617 ( 
.A(n_1712),
.Y(n_3617)
);

BUFx6f_ASAP7_75t_L g3618 ( 
.A(n_1031),
.Y(n_3618)
);

CKINVDCx5p33_ASAP7_75t_R g3619 ( 
.A(n_1637),
.Y(n_3619)
);

INVx2_ASAP7_75t_L g3620 ( 
.A(n_2310),
.Y(n_3620)
);

BUFx3_ASAP7_75t_L g3621 ( 
.A(n_2339),
.Y(n_3621)
);

CKINVDCx5p33_ASAP7_75t_R g3622 ( 
.A(n_1624),
.Y(n_3622)
);

CKINVDCx5p33_ASAP7_75t_R g3623 ( 
.A(n_87),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_2227),
.Y(n_3624)
);

CKINVDCx5p33_ASAP7_75t_R g3625 ( 
.A(n_2146),
.Y(n_3625)
);

CKINVDCx20_ASAP7_75t_R g3626 ( 
.A(n_1541),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_2382),
.Y(n_3627)
);

CKINVDCx5p33_ASAP7_75t_R g3628 ( 
.A(n_507),
.Y(n_3628)
);

CKINVDCx5p33_ASAP7_75t_R g3629 ( 
.A(n_866),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_2392),
.Y(n_3630)
);

INVx2_ASAP7_75t_SL g3631 ( 
.A(n_2256),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_1189),
.Y(n_3632)
);

CKINVDCx5p33_ASAP7_75t_R g3633 ( 
.A(n_136),
.Y(n_3633)
);

CKINVDCx5p33_ASAP7_75t_R g3634 ( 
.A(n_2459),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_2450),
.Y(n_3635)
);

INVx1_ASAP7_75t_SL g3636 ( 
.A(n_918),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_2314),
.Y(n_3637)
);

NOR2xp33_ASAP7_75t_L g3638 ( 
.A(n_715),
.B(n_1387),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_674),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_2265),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_37),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_1412),
.Y(n_3642)
);

CKINVDCx5p33_ASAP7_75t_R g3643 ( 
.A(n_1893),
.Y(n_3643)
);

CKINVDCx5p33_ASAP7_75t_R g3644 ( 
.A(n_427),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_655),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_1259),
.Y(n_3646)
);

CKINVDCx5p33_ASAP7_75t_R g3647 ( 
.A(n_2544),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_2268),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_L g3649 ( 
.A(n_2371),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_1383),
.Y(n_3650)
);

INVx1_ASAP7_75t_SL g3651 ( 
.A(n_2216),
.Y(n_3651)
);

CKINVDCx5p33_ASAP7_75t_R g3652 ( 
.A(n_791),
.Y(n_3652)
);

CKINVDCx5p33_ASAP7_75t_R g3653 ( 
.A(n_176),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_1965),
.Y(n_3654)
);

BUFx3_ASAP7_75t_L g3655 ( 
.A(n_2415),
.Y(n_3655)
);

CKINVDCx5p33_ASAP7_75t_R g3656 ( 
.A(n_508),
.Y(n_3656)
);

CKINVDCx5p33_ASAP7_75t_R g3657 ( 
.A(n_209),
.Y(n_3657)
);

CKINVDCx5p33_ASAP7_75t_R g3658 ( 
.A(n_2013),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_1509),
.Y(n_3659)
);

CKINVDCx5p33_ASAP7_75t_R g3660 ( 
.A(n_1899),
.Y(n_3660)
);

CKINVDCx5p33_ASAP7_75t_R g3661 ( 
.A(n_2330),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_82),
.Y(n_3662)
);

CKINVDCx5p33_ASAP7_75t_R g3663 ( 
.A(n_333),
.Y(n_3663)
);

CKINVDCx5p33_ASAP7_75t_R g3664 ( 
.A(n_1934),
.Y(n_3664)
);

CKINVDCx5p33_ASAP7_75t_R g3665 ( 
.A(n_391),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_906),
.Y(n_3666)
);

CKINVDCx5p33_ASAP7_75t_R g3667 ( 
.A(n_2528),
.Y(n_3667)
);

CKINVDCx5p33_ASAP7_75t_R g3668 ( 
.A(n_1037),
.Y(n_3668)
);

CKINVDCx5p33_ASAP7_75t_R g3669 ( 
.A(n_13),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_2363),
.Y(n_3670)
);

CKINVDCx5p33_ASAP7_75t_R g3671 ( 
.A(n_491),
.Y(n_3671)
);

CKINVDCx5p33_ASAP7_75t_R g3672 ( 
.A(n_265),
.Y(n_3672)
);

CKINVDCx5p33_ASAP7_75t_R g3673 ( 
.A(n_254),
.Y(n_3673)
);

CKINVDCx5p33_ASAP7_75t_R g3674 ( 
.A(n_2523),
.Y(n_3674)
);

CKINVDCx5p33_ASAP7_75t_R g3675 ( 
.A(n_1802),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_1420),
.Y(n_3676)
);

INVx1_ASAP7_75t_SL g3677 ( 
.A(n_679),
.Y(n_3677)
);

CKINVDCx5p33_ASAP7_75t_R g3678 ( 
.A(n_1440),
.Y(n_3678)
);

CKINVDCx5p33_ASAP7_75t_R g3679 ( 
.A(n_1413),
.Y(n_3679)
);

CKINVDCx5p33_ASAP7_75t_R g3680 ( 
.A(n_2011),
.Y(n_3680)
);

CKINVDCx5p33_ASAP7_75t_R g3681 ( 
.A(n_552),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_1569),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_177),
.Y(n_3683)
);

CKINVDCx5p33_ASAP7_75t_R g3684 ( 
.A(n_781),
.Y(n_3684)
);

CKINVDCx5p33_ASAP7_75t_R g3685 ( 
.A(n_562),
.Y(n_3685)
);

CKINVDCx5p33_ASAP7_75t_R g3686 ( 
.A(n_2325),
.Y(n_3686)
);

CKINVDCx5p33_ASAP7_75t_R g3687 ( 
.A(n_431),
.Y(n_3687)
);

CKINVDCx5p33_ASAP7_75t_R g3688 ( 
.A(n_1399),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_1066),
.Y(n_3689)
);

CKINVDCx20_ASAP7_75t_R g3690 ( 
.A(n_2086),
.Y(n_3690)
);

BUFx3_ASAP7_75t_L g3691 ( 
.A(n_1824),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_1621),
.Y(n_3692)
);

CKINVDCx5p33_ASAP7_75t_R g3693 ( 
.A(n_1584),
.Y(n_3693)
);

CKINVDCx5p33_ASAP7_75t_R g3694 ( 
.A(n_1629),
.Y(n_3694)
);

BUFx2_ASAP7_75t_R g3695 ( 
.A(n_2486),
.Y(n_3695)
);

BUFx3_ASAP7_75t_L g3696 ( 
.A(n_2005),
.Y(n_3696)
);

CKINVDCx5p33_ASAP7_75t_R g3697 ( 
.A(n_1858),
.Y(n_3697)
);

CKINVDCx5p33_ASAP7_75t_R g3698 ( 
.A(n_2260),
.Y(n_3698)
);

CKINVDCx5p33_ASAP7_75t_R g3699 ( 
.A(n_811),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_360),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_2311),
.Y(n_3701)
);

CKINVDCx5p33_ASAP7_75t_R g3702 ( 
.A(n_2085),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_2107),
.Y(n_3703)
);

CKINVDCx5p33_ASAP7_75t_R g3704 ( 
.A(n_2084),
.Y(n_3704)
);

CKINVDCx5p33_ASAP7_75t_R g3705 ( 
.A(n_1065),
.Y(n_3705)
);

CKINVDCx5p33_ASAP7_75t_R g3706 ( 
.A(n_912),
.Y(n_3706)
);

BUFx10_ASAP7_75t_L g3707 ( 
.A(n_2331),
.Y(n_3707)
);

CKINVDCx5p33_ASAP7_75t_R g3708 ( 
.A(n_746),
.Y(n_3708)
);

BUFx2_ASAP7_75t_L g3709 ( 
.A(n_498),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_2241),
.Y(n_3710)
);

CKINVDCx5p33_ASAP7_75t_R g3711 ( 
.A(n_952),
.Y(n_3711)
);

CKINVDCx5p33_ASAP7_75t_R g3712 ( 
.A(n_718),
.Y(n_3712)
);

CKINVDCx5p33_ASAP7_75t_R g3713 ( 
.A(n_2482),
.Y(n_3713)
);

CKINVDCx5p33_ASAP7_75t_R g3714 ( 
.A(n_949),
.Y(n_3714)
);

CKINVDCx5p33_ASAP7_75t_R g3715 ( 
.A(n_587),
.Y(n_3715)
);

CKINVDCx5p33_ASAP7_75t_R g3716 ( 
.A(n_1034),
.Y(n_3716)
);

CKINVDCx5p33_ASAP7_75t_R g3717 ( 
.A(n_1065),
.Y(n_3717)
);

CKINVDCx5p33_ASAP7_75t_R g3718 ( 
.A(n_2358),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_1718),
.Y(n_3719)
);

CKINVDCx5p33_ASAP7_75t_R g3720 ( 
.A(n_2087),
.Y(n_3720)
);

CKINVDCx5p33_ASAP7_75t_R g3721 ( 
.A(n_2320),
.Y(n_3721)
);

INVx2_ASAP7_75t_SL g3722 ( 
.A(n_2285),
.Y(n_3722)
);

CKINVDCx14_ASAP7_75t_R g3723 ( 
.A(n_526),
.Y(n_3723)
);

CKINVDCx5p33_ASAP7_75t_R g3724 ( 
.A(n_1747),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_1357),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_197),
.Y(n_3726)
);

CKINVDCx5p33_ASAP7_75t_R g3727 ( 
.A(n_737),
.Y(n_3727)
);

CKINVDCx5p33_ASAP7_75t_R g3728 ( 
.A(n_1580),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_1199),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_1235),
.Y(n_3730)
);

BUFx8_ASAP7_75t_SL g3731 ( 
.A(n_598),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_1876),
.Y(n_3732)
);

CKINVDCx5p33_ASAP7_75t_R g3733 ( 
.A(n_315),
.Y(n_3733)
);

INVx1_ASAP7_75t_SL g3734 ( 
.A(n_1556),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_2520),
.Y(n_3735)
);

HB1xp67_ASAP7_75t_L g3736 ( 
.A(n_1858),
.Y(n_3736)
);

CKINVDCx5p33_ASAP7_75t_R g3737 ( 
.A(n_760),
.Y(n_3737)
);

CKINVDCx5p33_ASAP7_75t_R g3738 ( 
.A(n_1870),
.Y(n_3738)
);

CKINVDCx5p33_ASAP7_75t_R g3739 ( 
.A(n_1038),
.Y(n_3739)
);

CKINVDCx5p33_ASAP7_75t_R g3740 ( 
.A(n_1953),
.Y(n_3740)
);

CKINVDCx20_ASAP7_75t_R g3741 ( 
.A(n_1749),
.Y(n_3741)
);

CKINVDCx5p33_ASAP7_75t_R g3742 ( 
.A(n_517),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_1843),
.Y(n_3743)
);

INVx3_ASAP7_75t_L g3744 ( 
.A(n_2424),
.Y(n_3744)
);

CKINVDCx5p33_ASAP7_75t_R g3745 ( 
.A(n_2190),
.Y(n_3745)
);

BUFx10_ASAP7_75t_L g3746 ( 
.A(n_1577),
.Y(n_3746)
);

CKINVDCx5p33_ASAP7_75t_R g3747 ( 
.A(n_1703),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_1539),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_318),
.Y(n_3749)
);

CKINVDCx5p33_ASAP7_75t_R g3750 ( 
.A(n_825),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_2280),
.Y(n_3751)
);

CKINVDCx5p33_ASAP7_75t_R g3752 ( 
.A(n_1904),
.Y(n_3752)
);

CKINVDCx5p33_ASAP7_75t_R g3753 ( 
.A(n_2521),
.Y(n_3753)
);

CKINVDCx5p33_ASAP7_75t_R g3754 ( 
.A(n_1267),
.Y(n_3754)
);

CKINVDCx5p33_ASAP7_75t_R g3755 ( 
.A(n_853),
.Y(n_3755)
);

CKINVDCx5p33_ASAP7_75t_R g3756 ( 
.A(n_2122),
.Y(n_3756)
);

CKINVDCx5p33_ASAP7_75t_R g3757 ( 
.A(n_1479),
.Y(n_3757)
);

CKINVDCx5p33_ASAP7_75t_R g3758 ( 
.A(n_1555),
.Y(n_3758)
);

INVxp67_ASAP7_75t_SL g3759 ( 
.A(n_1166),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_1455),
.Y(n_3760)
);

CKINVDCx5p33_ASAP7_75t_R g3761 ( 
.A(n_671),
.Y(n_3761)
);

CKINVDCx5p33_ASAP7_75t_R g3762 ( 
.A(n_1562),
.Y(n_3762)
);

CKINVDCx5p33_ASAP7_75t_R g3763 ( 
.A(n_2319),
.Y(n_3763)
);

CKINVDCx5p33_ASAP7_75t_R g3764 ( 
.A(n_1626),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_1303),
.Y(n_3765)
);

INVxp33_ASAP7_75t_L g3766 ( 
.A(n_2249),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_656),
.Y(n_3767)
);

CKINVDCx5p33_ASAP7_75t_R g3768 ( 
.A(n_2144),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_2065),
.Y(n_3769)
);

CKINVDCx5p33_ASAP7_75t_R g3770 ( 
.A(n_2521),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_1942),
.Y(n_3771)
);

CKINVDCx5p33_ASAP7_75t_R g3772 ( 
.A(n_390),
.Y(n_3772)
);

CKINVDCx5p33_ASAP7_75t_R g3773 ( 
.A(n_1242),
.Y(n_3773)
);

CKINVDCx20_ASAP7_75t_R g3774 ( 
.A(n_2362),
.Y(n_3774)
);

CKINVDCx20_ASAP7_75t_R g3775 ( 
.A(n_1568),
.Y(n_3775)
);

CKINVDCx5p33_ASAP7_75t_R g3776 ( 
.A(n_846),
.Y(n_3776)
);

CKINVDCx5p33_ASAP7_75t_R g3777 ( 
.A(n_555),
.Y(n_3777)
);

CKINVDCx5p33_ASAP7_75t_R g3778 ( 
.A(n_2446),
.Y(n_3778)
);

CKINVDCx5p33_ASAP7_75t_R g3779 ( 
.A(n_2306),
.Y(n_3779)
);

CKINVDCx5p33_ASAP7_75t_R g3780 ( 
.A(n_1074),
.Y(n_3780)
);

CKINVDCx5p33_ASAP7_75t_R g3781 ( 
.A(n_735),
.Y(n_3781)
);

CKINVDCx5p33_ASAP7_75t_R g3782 ( 
.A(n_2326),
.Y(n_3782)
);

CKINVDCx5p33_ASAP7_75t_R g3783 ( 
.A(n_608),
.Y(n_3783)
);

CKINVDCx5p33_ASAP7_75t_R g3784 ( 
.A(n_1982),
.Y(n_3784)
);

CKINVDCx5p33_ASAP7_75t_R g3785 ( 
.A(n_1848),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_2375),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_2440),
.Y(n_3787)
);

CKINVDCx5p33_ASAP7_75t_R g3788 ( 
.A(n_1312),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_1633),
.Y(n_3789)
);

CKINVDCx5p33_ASAP7_75t_R g3790 ( 
.A(n_2335),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_1125),
.Y(n_3791)
);

BUFx2_ASAP7_75t_SL g3792 ( 
.A(n_2178),
.Y(n_3792)
);

CKINVDCx5p33_ASAP7_75t_R g3793 ( 
.A(n_998),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_227),
.Y(n_3794)
);

CKINVDCx5p33_ASAP7_75t_R g3795 ( 
.A(n_1269),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_2135),
.Y(n_3796)
);

CKINVDCx5p33_ASAP7_75t_R g3797 ( 
.A(n_587),
.Y(n_3797)
);

BUFx6f_ASAP7_75t_L g3798 ( 
.A(n_216),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_962),
.Y(n_3799)
);

BUFx6f_ASAP7_75t_L g3800 ( 
.A(n_592),
.Y(n_3800)
);

CKINVDCx16_ASAP7_75t_R g3801 ( 
.A(n_2179),
.Y(n_3801)
);

CKINVDCx5p33_ASAP7_75t_R g3802 ( 
.A(n_1694),
.Y(n_3802)
);

CKINVDCx5p33_ASAP7_75t_R g3803 ( 
.A(n_878),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_2512),
.Y(n_3804)
);

HB1xp67_ASAP7_75t_L g3805 ( 
.A(n_2320),
.Y(n_3805)
);

CKINVDCx5p33_ASAP7_75t_R g3806 ( 
.A(n_1969),
.Y(n_3806)
);

CKINVDCx5p33_ASAP7_75t_R g3807 ( 
.A(n_1631),
.Y(n_3807)
);

CKINVDCx14_ASAP7_75t_R g3808 ( 
.A(n_2286),
.Y(n_3808)
);

CKINVDCx5p33_ASAP7_75t_R g3809 ( 
.A(n_2109),
.Y(n_3809)
);

CKINVDCx5p33_ASAP7_75t_R g3810 ( 
.A(n_584),
.Y(n_3810)
);

CKINVDCx5p33_ASAP7_75t_R g3811 ( 
.A(n_314),
.Y(n_3811)
);

BUFx6f_ASAP7_75t_L g3812 ( 
.A(n_2028),
.Y(n_3812)
);

CKINVDCx5p33_ASAP7_75t_R g3813 ( 
.A(n_2544),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_319),
.Y(n_3814)
);

INVx1_ASAP7_75t_SL g3815 ( 
.A(n_515),
.Y(n_3815)
);

CKINVDCx5p33_ASAP7_75t_R g3816 ( 
.A(n_1116),
.Y(n_3816)
);

INVxp67_ASAP7_75t_L g3817 ( 
.A(n_1379),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_1602),
.Y(n_3818)
);

CKINVDCx5p33_ASAP7_75t_R g3819 ( 
.A(n_2279),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_2192),
.Y(n_3820)
);

BUFx6f_ASAP7_75t_L g3821 ( 
.A(n_31),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_2505),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_514),
.Y(n_3823)
);

CKINVDCx20_ASAP7_75t_R g3824 ( 
.A(n_1555),
.Y(n_3824)
);

INVx1_ASAP7_75t_SL g3825 ( 
.A(n_1671),
.Y(n_3825)
);

CKINVDCx5p33_ASAP7_75t_R g3826 ( 
.A(n_662),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_1277),
.Y(n_3827)
);

CKINVDCx5p33_ASAP7_75t_R g3828 ( 
.A(n_1217),
.Y(n_3828)
);

CKINVDCx5p33_ASAP7_75t_R g3829 ( 
.A(n_1283),
.Y(n_3829)
);

CKINVDCx5p33_ASAP7_75t_R g3830 ( 
.A(n_1046),
.Y(n_3830)
);

CKINVDCx5p33_ASAP7_75t_R g3831 ( 
.A(n_2361),
.Y(n_3831)
);

CKINVDCx5p33_ASAP7_75t_R g3832 ( 
.A(n_2285),
.Y(n_3832)
);

INVx1_ASAP7_75t_SL g3833 ( 
.A(n_1874),
.Y(n_3833)
);

CKINVDCx5p33_ASAP7_75t_R g3834 ( 
.A(n_1230),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_2146),
.Y(n_3835)
);

CKINVDCx5p33_ASAP7_75t_R g3836 ( 
.A(n_1905),
.Y(n_3836)
);

BUFx2_ASAP7_75t_L g3837 ( 
.A(n_2132),
.Y(n_3837)
);

CKINVDCx5p33_ASAP7_75t_R g3838 ( 
.A(n_70),
.Y(n_3838)
);

CKINVDCx5p33_ASAP7_75t_R g3839 ( 
.A(n_2283),
.Y(n_3839)
);

CKINVDCx5p33_ASAP7_75t_R g3840 ( 
.A(n_2483),
.Y(n_3840)
);

CKINVDCx5p33_ASAP7_75t_R g3841 ( 
.A(n_1338),
.Y(n_3841)
);

CKINVDCx5p33_ASAP7_75t_R g3842 ( 
.A(n_558),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_1477),
.Y(n_3843)
);

BUFx10_ASAP7_75t_L g3844 ( 
.A(n_1222),
.Y(n_3844)
);

CKINVDCx5p33_ASAP7_75t_R g3845 ( 
.A(n_2530),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_776),
.Y(n_3846)
);

CKINVDCx5p33_ASAP7_75t_R g3847 ( 
.A(n_725),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_2220),
.Y(n_3848)
);

CKINVDCx16_ASAP7_75t_R g3849 ( 
.A(n_75),
.Y(n_3849)
);

CKINVDCx5p33_ASAP7_75t_R g3850 ( 
.A(n_2336),
.Y(n_3850)
);

CKINVDCx5p33_ASAP7_75t_R g3851 ( 
.A(n_829),
.Y(n_3851)
);

CKINVDCx5p33_ASAP7_75t_R g3852 ( 
.A(n_1983),
.Y(n_3852)
);

CKINVDCx5p33_ASAP7_75t_R g3853 ( 
.A(n_2448),
.Y(n_3853)
);

CKINVDCx5p33_ASAP7_75t_R g3854 ( 
.A(n_1105),
.Y(n_3854)
);

CKINVDCx5p33_ASAP7_75t_R g3855 ( 
.A(n_795),
.Y(n_3855)
);

CKINVDCx5p33_ASAP7_75t_R g3856 ( 
.A(n_319),
.Y(n_3856)
);

CKINVDCx5p33_ASAP7_75t_R g3857 ( 
.A(n_641),
.Y(n_3857)
);

CKINVDCx20_ASAP7_75t_R g3858 ( 
.A(n_203),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_2418),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_2290),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_261),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_2403),
.Y(n_3862)
);

CKINVDCx5p33_ASAP7_75t_R g3863 ( 
.A(n_2034),
.Y(n_3863)
);

CKINVDCx5p33_ASAP7_75t_R g3864 ( 
.A(n_1732),
.Y(n_3864)
);

CKINVDCx16_ASAP7_75t_R g3865 ( 
.A(n_1834),
.Y(n_3865)
);

BUFx5_ASAP7_75t_L g3866 ( 
.A(n_1289),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_2241),
.Y(n_3867)
);

CKINVDCx5p33_ASAP7_75t_R g3868 ( 
.A(n_1860),
.Y(n_3868)
);

CKINVDCx5p33_ASAP7_75t_R g3869 ( 
.A(n_1861),
.Y(n_3869)
);

CKINVDCx20_ASAP7_75t_R g3870 ( 
.A(n_872),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_2370),
.Y(n_3871)
);

CKINVDCx5p33_ASAP7_75t_R g3872 ( 
.A(n_1445),
.Y(n_3872)
);

CKINVDCx16_ASAP7_75t_R g3873 ( 
.A(n_917),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_223),
.Y(n_3874)
);

CKINVDCx5p33_ASAP7_75t_R g3875 ( 
.A(n_1475),
.Y(n_3875)
);

CKINVDCx5p33_ASAP7_75t_R g3876 ( 
.A(n_32),
.Y(n_3876)
);

CKINVDCx5p33_ASAP7_75t_R g3877 ( 
.A(n_1378),
.Y(n_3877)
);

CKINVDCx5p33_ASAP7_75t_R g3878 ( 
.A(n_2303),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_1844),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_2103),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_428),
.Y(n_3881)
);

CKINVDCx5p33_ASAP7_75t_R g3882 ( 
.A(n_2542),
.Y(n_3882)
);

HB1xp67_ASAP7_75t_L g3883 ( 
.A(n_972),
.Y(n_3883)
);

BUFx10_ASAP7_75t_L g3884 ( 
.A(n_2158),
.Y(n_3884)
);

CKINVDCx5p33_ASAP7_75t_R g3885 ( 
.A(n_544),
.Y(n_3885)
);

CKINVDCx5p33_ASAP7_75t_R g3886 ( 
.A(n_1433),
.Y(n_3886)
);

CKINVDCx5p33_ASAP7_75t_R g3887 ( 
.A(n_2229),
.Y(n_3887)
);

CKINVDCx5p33_ASAP7_75t_R g3888 ( 
.A(n_1924),
.Y(n_3888)
);

CKINVDCx5p33_ASAP7_75t_R g3889 ( 
.A(n_640),
.Y(n_3889)
);

CKINVDCx5p33_ASAP7_75t_R g3890 ( 
.A(n_1390),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_1437),
.Y(n_3891)
);

CKINVDCx5p33_ASAP7_75t_R g3892 ( 
.A(n_988),
.Y(n_3892)
);

CKINVDCx5p33_ASAP7_75t_R g3893 ( 
.A(n_1225),
.Y(n_3893)
);

CKINVDCx5p33_ASAP7_75t_R g3894 ( 
.A(n_2515),
.Y(n_3894)
);

CKINVDCx5p33_ASAP7_75t_R g3895 ( 
.A(n_2177),
.Y(n_3895)
);

CKINVDCx5p33_ASAP7_75t_R g3896 ( 
.A(n_1471),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_176),
.Y(n_3897)
);

CKINVDCx5p33_ASAP7_75t_R g3898 ( 
.A(n_2289),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_467),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_250),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_2259),
.Y(n_3901)
);

CKINVDCx5p33_ASAP7_75t_R g3902 ( 
.A(n_1960),
.Y(n_3902)
);

CKINVDCx20_ASAP7_75t_R g3903 ( 
.A(n_1933),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_280),
.Y(n_3904)
);

CKINVDCx5p33_ASAP7_75t_R g3905 ( 
.A(n_2266),
.Y(n_3905)
);

CKINVDCx5p33_ASAP7_75t_R g3906 ( 
.A(n_2498),
.Y(n_3906)
);

INVxp33_ASAP7_75t_L g3907 ( 
.A(n_1319),
.Y(n_3907)
);

CKINVDCx5p33_ASAP7_75t_R g3908 ( 
.A(n_2277),
.Y(n_3908)
);

CKINVDCx5p33_ASAP7_75t_R g3909 ( 
.A(n_290),
.Y(n_3909)
);

CKINVDCx5p33_ASAP7_75t_R g3910 ( 
.A(n_922),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_1045),
.Y(n_3911)
);

CKINVDCx5p33_ASAP7_75t_R g3912 ( 
.A(n_1151),
.Y(n_3912)
);

CKINVDCx5p33_ASAP7_75t_R g3913 ( 
.A(n_2309),
.Y(n_3913)
);

CKINVDCx5p33_ASAP7_75t_R g3914 ( 
.A(n_2141),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_112),
.Y(n_3915)
);

CKINVDCx20_ASAP7_75t_R g3916 ( 
.A(n_1938),
.Y(n_3916)
);

CKINVDCx5p33_ASAP7_75t_R g3917 ( 
.A(n_1345),
.Y(n_3917)
);

CKINVDCx5p33_ASAP7_75t_R g3918 ( 
.A(n_677),
.Y(n_3918)
);

CKINVDCx5p33_ASAP7_75t_R g3919 ( 
.A(n_1676),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_320),
.Y(n_3920)
);

CKINVDCx5p33_ASAP7_75t_R g3921 ( 
.A(n_417),
.Y(n_3921)
);

CKINVDCx5p33_ASAP7_75t_R g3922 ( 
.A(n_1231),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_972),
.Y(n_3923)
);

CKINVDCx5p33_ASAP7_75t_R g3924 ( 
.A(n_365),
.Y(n_3924)
);

CKINVDCx5p33_ASAP7_75t_R g3925 ( 
.A(n_2255),
.Y(n_3925)
);

BUFx2_ASAP7_75t_L g3926 ( 
.A(n_2307),
.Y(n_3926)
);

CKINVDCx20_ASAP7_75t_R g3927 ( 
.A(n_2554),
.Y(n_3927)
);

CKINVDCx5p33_ASAP7_75t_R g3928 ( 
.A(n_1153),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_1080),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_1216),
.Y(n_3930)
);

CKINVDCx5p33_ASAP7_75t_R g3931 ( 
.A(n_1165),
.Y(n_3931)
);

CKINVDCx5p33_ASAP7_75t_R g3932 ( 
.A(n_1707),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_1210),
.Y(n_3933)
);

CKINVDCx5p33_ASAP7_75t_R g3934 ( 
.A(n_2335),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_878),
.Y(n_3935)
);

CKINVDCx5p33_ASAP7_75t_R g3936 ( 
.A(n_928),
.Y(n_3936)
);

CKINVDCx5p33_ASAP7_75t_R g3937 ( 
.A(n_1733),
.Y(n_3937)
);

CKINVDCx20_ASAP7_75t_R g3938 ( 
.A(n_1761),
.Y(n_3938)
);

CKINVDCx5p33_ASAP7_75t_R g3939 ( 
.A(n_1230),
.Y(n_3939)
);

CKINVDCx5p33_ASAP7_75t_R g3940 ( 
.A(n_135),
.Y(n_3940)
);

CKINVDCx14_ASAP7_75t_R g3941 ( 
.A(n_165),
.Y(n_3941)
);

CKINVDCx5p33_ASAP7_75t_R g3942 ( 
.A(n_135),
.Y(n_3942)
);

CKINVDCx5p33_ASAP7_75t_R g3943 ( 
.A(n_369),
.Y(n_3943)
);

CKINVDCx5p33_ASAP7_75t_R g3944 ( 
.A(n_1958),
.Y(n_3944)
);

BUFx10_ASAP7_75t_L g3945 ( 
.A(n_617),
.Y(n_3945)
);

CKINVDCx5p33_ASAP7_75t_R g3946 ( 
.A(n_1162),
.Y(n_3946)
);

CKINVDCx5p33_ASAP7_75t_R g3947 ( 
.A(n_33),
.Y(n_3947)
);

CKINVDCx5p33_ASAP7_75t_R g3948 ( 
.A(n_422),
.Y(n_3948)
);

CKINVDCx5p33_ASAP7_75t_R g3949 ( 
.A(n_1083),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_2257),
.Y(n_3950)
);

CKINVDCx5p33_ASAP7_75t_R g3951 ( 
.A(n_1809),
.Y(n_3951)
);

CKINVDCx5p33_ASAP7_75t_R g3952 ( 
.A(n_1470),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_1308),
.Y(n_3953)
);

CKINVDCx5p33_ASAP7_75t_R g3954 ( 
.A(n_2065),
.Y(n_3954)
);

CKINVDCx20_ASAP7_75t_R g3955 ( 
.A(n_2380),
.Y(n_3955)
);

CKINVDCx5p33_ASAP7_75t_R g3956 ( 
.A(n_1383),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_2523),
.Y(n_3957)
);

CKINVDCx5p33_ASAP7_75t_R g3958 ( 
.A(n_1847),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_191),
.Y(n_3959)
);

CKINVDCx5p33_ASAP7_75t_R g3960 ( 
.A(n_2288),
.Y(n_3960)
);

CKINVDCx5p33_ASAP7_75t_R g3961 ( 
.A(n_2008),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_1196),
.Y(n_3962)
);

CKINVDCx5p33_ASAP7_75t_R g3963 ( 
.A(n_1112),
.Y(n_3963)
);

INVxp67_ASAP7_75t_L g3964 ( 
.A(n_785),
.Y(n_3964)
);

BUFx2_ASAP7_75t_L g3965 ( 
.A(n_1158),
.Y(n_3965)
);

INVx2_ASAP7_75t_SL g3966 ( 
.A(n_2368),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_2344),
.Y(n_3967)
);

INVx2_ASAP7_75t_SL g3968 ( 
.A(n_1511),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_1903),
.Y(n_3969)
);

CKINVDCx5p33_ASAP7_75t_R g3970 ( 
.A(n_961),
.Y(n_3970)
);

CKINVDCx5p33_ASAP7_75t_R g3971 ( 
.A(n_1877),
.Y(n_3971)
);

BUFx2_ASAP7_75t_L g3972 ( 
.A(n_267),
.Y(n_3972)
);

CKINVDCx5p33_ASAP7_75t_R g3973 ( 
.A(n_1679),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_2532),
.Y(n_3974)
);

CKINVDCx20_ASAP7_75t_R g3975 ( 
.A(n_2092),
.Y(n_3975)
);

CKINVDCx5p33_ASAP7_75t_R g3976 ( 
.A(n_830),
.Y(n_3976)
);

INVx2_ASAP7_75t_SL g3977 ( 
.A(n_1692),
.Y(n_3977)
);

CKINVDCx5p33_ASAP7_75t_R g3978 ( 
.A(n_1292),
.Y(n_3978)
);

INVx2_ASAP7_75t_L g3979 ( 
.A(n_947),
.Y(n_3979)
);

BUFx10_ASAP7_75t_L g3980 ( 
.A(n_113),
.Y(n_3980)
);

CKINVDCx20_ASAP7_75t_R g3981 ( 
.A(n_1241),
.Y(n_3981)
);

CKINVDCx5p33_ASAP7_75t_R g3982 ( 
.A(n_1898),
.Y(n_3982)
);

INVxp67_ASAP7_75t_L g3983 ( 
.A(n_1809),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_2172),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_1956),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_862),
.Y(n_3986)
);

CKINVDCx5p33_ASAP7_75t_R g3987 ( 
.A(n_2042),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_2253),
.Y(n_3988)
);

BUFx6f_ASAP7_75t_L g3989 ( 
.A(n_425),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_2082),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_2546),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_1177),
.Y(n_3992)
);

CKINVDCx5p33_ASAP7_75t_R g3993 ( 
.A(n_1771),
.Y(n_3993)
);

CKINVDCx5p33_ASAP7_75t_R g3994 ( 
.A(n_1274),
.Y(n_3994)
);

CKINVDCx5p33_ASAP7_75t_R g3995 ( 
.A(n_681),
.Y(n_3995)
);

CKINVDCx20_ASAP7_75t_R g3996 ( 
.A(n_157),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_49),
.Y(n_3997)
);

INVx1_ASAP7_75t_SL g3998 ( 
.A(n_1762),
.Y(n_3998)
);

CKINVDCx20_ASAP7_75t_R g3999 ( 
.A(n_682),
.Y(n_3999)
);

CKINVDCx5p33_ASAP7_75t_R g4000 ( 
.A(n_161),
.Y(n_4000)
);

BUFx3_ASAP7_75t_L g4001 ( 
.A(n_1464),
.Y(n_4001)
);

CKINVDCx20_ASAP7_75t_R g4002 ( 
.A(n_1510),
.Y(n_4002)
);

CKINVDCx5p33_ASAP7_75t_R g4003 ( 
.A(n_2401),
.Y(n_4003)
);

CKINVDCx5p33_ASAP7_75t_R g4004 ( 
.A(n_2328),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_303),
.Y(n_4005)
);

CKINVDCx5p33_ASAP7_75t_R g4006 ( 
.A(n_1073),
.Y(n_4006)
);

CKINVDCx5p33_ASAP7_75t_R g4007 ( 
.A(n_611),
.Y(n_4007)
);

CKINVDCx20_ASAP7_75t_R g4008 ( 
.A(n_1106),
.Y(n_4008)
);

BUFx10_ASAP7_75t_L g4009 ( 
.A(n_2284),
.Y(n_4009)
);

BUFx5_ASAP7_75t_L g4010 ( 
.A(n_622),
.Y(n_4010)
);

CKINVDCx5p33_ASAP7_75t_R g4011 ( 
.A(n_1525),
.Y(n_4011)
);

BUFx3_ASAP7_75t_L g4012 ( 
.A(n_429),
.Y(n_4012)
);

CKINVDCx5p33_ASAP7_75t_R g4013 ( 
.A(n_2040),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_2365),
.Y(n_4014)
);

BUFx3_ASAP7_75t_L g4015 ( 
.A(n_733),
.Y(n_4015)
);

CKINVDCx5p33_ASAP7_75t_R g4016 ( 
.A(n_2205),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_1512),
.Y(n_4017)
);

CKINVDCx5p33_ASAP7_75t_R g4018 ( 
.A(n_749),
.Y(n_4018)
);

CKINVDCx20_ASAP7_75t_R g4019 ( 
.A(n_1993),
.Y(n_4019)
);

CKINVDCx5p33_ASAP7_75t_R g4020 ( 
.A(n_2433),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_2437),
.Y(n_4021)
);

CKINVDCx5p33_ASAP7_75t_R g4022 ( 
.A(n_2311),
.Y(n_4022)
);

CKINVDCx5p33_ASAP7_75t_R g4023 ( 
.A(n_2293),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_1408),
.Y(n_4024)
);

CKINVDCx5p33_ASAP7_75t_R g4025 ( 
.A(n_740),
.Y(n_4025)
);

CKINVDCx5p33_ASAP7_75t_R g4026 ( 
.A(n_834),
.Y(n_4026)
);

BUFx6f_ASAP7_75t_L g4027 ( 
.A(n_899),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_605),
.Y(n_4028)
);

CKINVDCx5p33_ASAP7_75t_R g4029 ( 
.A(n_173),
.Y(n_4029)
);

CKINVDCx5p33_ASAP7_75t_R g4030 ( 
.A(n_1841),
.Y(n_4030)
);

BUFx2_ASAP7_75t_L g4031 ( 
.A(n_1404),
.Y(n_4031)
);

CKINVDCx5p33_ASAP7_75t_R g4032 ( 
.A(n_2364),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_2391),
.Y(n_4033)
);

BUFx2_ASAP7_75t_L g4034 ( 
.A(n_350),
.Y(n_4034)
);

CKINVDCx5p33_ASAP7_75t_R g4035 ( 
.A(n_925),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_1718),
.Y(n_4036)
);

CKINVDCx5p33_ASAP7_75t_R g4037 ( 
.A(n_865),
.Y(n_4037)
);

BUFx2_ASAP7_75t_L g4038 ( 
.A(n_2137),
.Y(n_4038)
);

CKINVDCx5p33_ASAP7_75t_R g4039 ( 
.A(n_2300),
.Y(n_4039)
);

CKINVDCx5p33_ASAP7_75t_R g4040 ( 
.A(n_1112),
.Y(n_4040)
);

CKINVDCx5p33_ASAP7_75t_R g4041 ( 
.A(n_1137),
.Y(n_4041)
);

CKINVDCx5p33_ASAP7_75t_R g4042 ( 
.A(n_647),
.Y(n_4042)
);

CKINVDCx5p33_ASAP7_75t_R g4043 ( 
.A(n_1210),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_881),
.Y(n_4044)
);

CKINVDCx16_ASAP7_75t_R g4045 ( 
.A(n_2214),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_2129),
.Y(n_4046)
);

CKINVDCx5p33_ASAP7_75t_R g4047 ( 
.A(n_635),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_2405),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_2529),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_1953),
.Y(n_4050)
);

CKINVDCx5p33_ASAP7_75t_R g4051 ( 
.A(n_2055),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_897),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_264),
.Y(n_4053)
);

CKINVDCx5p33_ASAP7_75t_R g4054 ( 
.A(n_924),
.Y(n_4054)
);

INVxp67_ASAP7_75t_L g4055 ( 
.A(n_2566),
.Y(n_4055)
);

BUFx3_ASAP7_75t_L g4056 ( 
.A(n_3164),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3164),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3291),
.Y(n_4058)
);

CKINVDCx5p33_ASAP7_75t_R g4059 ( 
.A(n_3084),
.Y(n_4059)
);

CKINVDCx5p33_ASAP7_75t_R g4060 ( 
.A(n_3315),
.Y(n_4060)
);

INVxp67_ASAP7_75t_L g4061 ( 
.A(n_2606),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3291),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3310),
.Y(n_4063)
);

BUFx5_ASAP7_75t_L g4064 ( 
.A(n_2558),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3310),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3352),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3352),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3744),
.Y(n_4068)
);

INVxp33_ASAP7_75t_L g4069 ( 
.A(n_3353),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3744),
.Y(n_4070)
);

INVxp33_ASAP7_75t_SL g4071 ( 
.A(n_2919),
.Y(n_4071)
);

CKINVDCx16_ASAP7_75t_R g4072 ( 
.A(n_2923),
.Y(n_4072)
);

CKINVDCx5p33_ASAP7_75t_R g4073 ( 
.A(n_3381),
.Y(n_4073)
);

CKINVDCx16_ASAP7_75t_R g4074 ( 
.A(n_3108),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_2604),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_2604),
.Y(n_4076)
);

INVx2_ASAP7_75t_L g4077 ( 
.A(n_2604),
.Y(n_4077)
);

CKINVDCx5p33_ASAP7_75t_R g4078 ( 
.A(n_3731),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_2604),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_2604),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_2614),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_2614),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_2614),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_2614),
.Y(n_4084)
);

BUFx6f_ASAP7_75t_L g4085 ( 
.A(n_2700),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_2614),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_2781),
.Y(n_4087)
);

CKINVDCx5p33_ASAP7_75t_R g4088 ( 
.A(n_3339),
.Y(n_4088)
);

BUFx6f_ASAP7_75t_L g4089 ( 
.A(n_2700),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_2781),
.Y(n_4090)
);

BUFx6f_ASAP7_75t_L g4091 ( 
.A(n_2700),
.Y(n_4091)
);

CKINVDCx5p33_ASAP7_75t_R g4092 ( 
.A(n_3723),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_2781),
.Y(n_4093)
);

INVx2_ASAP7_75t_L g4094 ( 
.A(n_2781),
.Y(n_4094)
);

BUFx3_ASAP7_75t_L g4095 ( 
.A(n_2556),
.Y(n_4095)
);

INVxp67_ASAP7_75t_SL g4096 ( 
.A(n_2702),
.Y(n_4096)
);

BUFx2_ASAP7_75t_L g4097 ( 
.A(n_3808),
.Y(n_4097)
);

CKINVDCx16_ASAP7_75t_R g4098 ( 
.A(n_3941),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_2781),
.Y(n_4099)
);

NOR2xp33_ASAP7_75t_L g4100 ( 
.A(n_2870),
.B(n_0),
.Y(n_4100)
);

BUFx2_ASAP7_75t_SL g4101 ( 
.A(n_3307),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3248),
.Y(n_4102)
);

CKINVDCx5p33_ASAP7_75t_R g4103 ( 
.A(n_2571),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3248),
.Y(n_4104)
);

CKINVDCx20_ASAP7_75t_R g4105 ( 
.A(n_2687),
.Y(n_4105)
);

CKINVDCx5p33_ASAP7_75t_R g4106 ( 
.A(n_2602),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_3248),
.Y(n_4107)
);

CKINVDCx5p33_ASAP7_75t_R g4108 ( 
.A(n_2633),
.Y(n_4108)
);

CKINVDCx5p33_ASAP7_75t_R g4109 ( 
.A(n_2722),
.Y(n_4109)
);

CKINVDCx5p33_ASAP7_75t_R g4110 ( 
.A(n_2782),
.Y(n_4110)
);

CKINVDCx16_ASAP7_75t_R g4111 ( 
.A(n_3000),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3248),
.Y(n_4112)
);

CKINVDCx5p33_ASAP7_75t_R g4113 ( 
.A(n_2911),
.Y(n_4113)
);

CKINVDCx5p33_ASAP7_75t_R g4114 ( 
.A(n_2942),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3248),
.Y(n_4115)
);

CKINVDCx5p33_ASAP7_75t_R g4116 ( 
.A(n_3023),
.Y(n_4116)
);

CKINVDCx5p33_ASAP7_75t_R g4117 ( 
.A(n_3125),
.Y(n_4117)
);

CKINVDCx16_ASAP7_75t_R g4118 ( 
.A(n_3029),
.Y(n_4118)
);

CKINVDCx5p33_ASAP7_75t_R g4119 ( 
.A(n_3146),
.Y(n_4119)
);

BUFx2_ASAP7_75t_L g4120 ( 
.A(n_3050),
.Y(n_4120)
);

CKINVDCx5p33_ASAP7_75t_R g4121 ( 
.A(n_3207),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3392),
.Y(n_4122)
);

CKINVDCx5p33_ASAP7_75t_R g4123 ( 
.A(n_3296),
.Y(n_4123)
);

CKINVDCx5p33_ASAP7_75t_R g4124 ( 
.A(n_3370),
.Y(n_4124)
);

CKINVDCx5p33_ASAP7_75t_R g4125 ( 
.A(n_3377),
.Y(n_4125)
);

NOR2xp33_ASAP7_75t_L g4126 ( 
.A(n_2949),
.B(n_0),
.Y(n_4126)
);

CKINVDCx5p33_ASAP7_75t_R g4127 ( 
.A(n_3434),
.Y(n_4127)
);

CKINVDCx5p33_ASAP7_75t_R g4128 ( 
.A(n_3484),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3392),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3392),
.Y(n_4130)
);

INVx2_ASAP7_75t_SL g4131 ( 
.A(n_2568),
.Y(n_4131)
);

CKINVDCx5p33_ASAP7_75t_R g4132 ( 
.A(n_3490),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3392),
.Y(n_4133)
);

BUFx2_ASAP7_75t_L g4134 ( 
.A(n_3101),
.Y(n_4134)
);

CKINVDCx20_ASAP7_75t_R g4135 ( 
.A(n_3927),
.Y(n_4135)
);

CKINVDCx5p33_ASAP7_75t_R g4136 ( 
.A(n_3497),
.Y(n_4136)
);

CKINVDCx5p33_ASAP7_75t_R g4137 ( 
.A(n_3499),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_3392),
.Y(n_4138)
);

INVx1_ASAP7_75t_SL g4139 ( 
.A(n_3695),
.Y(n_4139)
);

INVxp67_ASAP7_75t_SL g4140 ( 
.A(n_2702),
.Y(n_4140)
);

BUFx3_ASAP7_75t_L g4141 ( 
.A(n_2598),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_3410),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3410),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3410),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3410),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3410),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_3541),
.Y(n_4147)
);

HB1xp67_ASAP7_75t_L g4148 ( 
.A(n_3107),
.Y(n_4148)
);

CKINVDCx20_ASAP7_75t_R g4149 ( 
.A(n_2583),
.Y(n_4149)
);

CKINVDCx20_ASAP7_75t_R g4150 ( 
.A(n_2586),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_3541),
.Y(n_4151)
);

CKINVDCx5p33_ASAP7_75t_R g4152 ( 
.A(n_3527),
.Y(n_4152)
);

CKINVDCx5p33_ASAP7_75t_R g4153 ( 
.A(n_3598),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3541),
.Y(n_4154)
);

CKINVDCx5p33_ASAP7_75t_R g4155 ( 
.A(n_3634),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3541),
.Y(n_4156)
);

INVxp67_ASAP7_75t_L g4157 ( 
.A(n_2720),
.Y(n_4157)
);

CKINVDCx5p33_ASAP7_75t_R g4158 ( 
.A(n_3647),
.Y(n_4158)
);

BUFx6f_ASAP7_75t_L g4159 ( 
.A(n_2702),
.Y(n_4159)
);

BUFx3_ASAP7_75t_L g4160 ( 
.A(n_2618),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3541),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_3866),
.Y(n_4162)
);

CKINVDCx5p33_ASAP7_75t_R g4163 ( 
.A(n_3667),
.Y(n_4163)
);

CKINVDCx5p33_ASAP7_75t_R g4164 ( 
.A(n_3674),
.Y(n_4164)
);

CKINVDCx5p33_ASAP7_75t_R g4165 ( 
.A(n_3713),
.Y(n_4165)
);

BUFx6f_ASAP7_75t_L g4166 ( 
.A(n_2712),
.Y(n_4166)
);

BUFx6f_ASAP7_75t_L g4167 ( 
.A(n_2712),
.Y(n_4167)
);

CKINVDCx5p33_ASAP7_75t_R g4168 ( 
.A(n_3753),
.Y(n_4168)
);

XOR2x2_ASAP7_75t_L g4169 ( 
.A(n_3128),
.B(n_1),
.Y(n_4169)
);

BUFx2_ASAP7_75t_L g4170 ( 
.A(n_3289),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3866),
.Y(n_4171)
);

CKINVDCx5p33_ASAP7_75t_R g4172 ( 
.A(n_3770),
.Y(n_4172)
);

INVx2_ASAP7_75t_SL g4173 ( 
.A(n_2568),
.Y(n_4173)
);

BUFx2_ASAP7_75t_L g4174 ( 
.A(n_3378),
.Y(n_4174)
);

CKINVDCx5p33_ASAP7_75t_R g4175 ( 
.A(n_3813),
.Y(n_4175)
);

INVx1_ASAP7_75t_SL g4176 ( 
.A(n_3403),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3866),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3866),
.Y(n_4178)
);

CKINVDCx5p33_ASAP7_75t_R g4179 ( 
.A(n_3840),
.Y(n_4179)
);

CKINVDCx5p33_ASAP7_75t_R g4180 ( 
.A(n_3845),
.Y(n_4180)
);

CKINVDCx20_ASAP7_75t_R g4181 ( 
.A(n_2590),
.Y(n_4181)
);

CKINVDCx5p33_ASAP7_75t_R g4182 ( 
.A(n_3882),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3866),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_4010),
.Y(n_4184)
);

INVx1_ASAP7_75t_SL g4185 ( 
.A(n_3441),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_4010),
.Y(n_4186)
);

INVx2_ASAP7_75t_L g4187 ( 
.A(n_4010),
.Y(n_4187)
);

CKINVDCx20_ASAP7_75t_R g4188 ( 
.A(n_2594),
.Y(n_4188)
);

CKINVDCx5p33_ASAP7_75t_R g4189 ( 
.A(n_3894),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4010),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4010),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_3307),
.Y(n_4192)
);

CKINVDCx5p33_ASAP7_75t_R g4193 ( 
.A(n_3906),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_2712),
.Y(n_4194)
);

CKINVDCx5p33_ASAP7_75t_R g4195 ( 
.A(n_2555),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_2737),
.Y(n_4196)
);

CKINVDCx16_ASAP7_75t_R g4197 ( 
.A(n_3567),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_2737),
.Y(n_4198)
);

CKINVDCx5p33_ASAP7_75t_R g4199 ( 
.A(n_2557),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_2737),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_2761),
.Y(n_4201)
);

HB1xp67_ASAP7_75t_L g4202 ( 
.A(n_3595),
.Y(n_4202)
);

CKINVDCx20_ASAP7_75t_R g4203 ( 
.A(n_2626),
.Y(n_4203)
);

CKINVDCx14_ASAP7_75t_R g4204 ( 
.A(n_2634),
.Y(n_4204)
);

CKINVDCx5p33_ASAP7_75t_R g4205 ( 
.A(n_2559),
.Y(n_4205)
);

INVx2_ASAP7_75t_SL g4206 ( 
.A(n_2634),
.Y(n_4206)
);

CKINVDCx5p33_ASAP7_75t_R g4207 ( 
.A(n_2560),
.Y(n_4207)
);

CKINVDCx5p33_ASAP7_75t_R g4208 ( 
.A(n_2562),
.Y(n_4208)
);

CKINVDCx5p33_ASAP7_75t_R g4209 ( 
.A(n_2564),
.Y(n_4209)
);

CKINVDCx5p33_ASAP7_75t_R g4210 ( 
.A(n_2565),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_2761),
.Y(n_4211)
);

CKINVDCx5p33_ASAP7_75t_R g4212 ( 
.A(n_2567),
.Y(n_4212)
);

INVxp67_ASAP7_75t_SL g4213 ( 
.A(n_2761),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_2791),
.Y(n_4214)
);

CKINVDCx5p33_ASAP7_75t_R g4215 ( 
.A(n_2570),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_2791),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_2791),
.Y(n_4217)
);

INVx1_ASAP7_75t_SL g4218 ( 
.A(n_3801),
.Y(n_4218)
);

BUFx5_ASAP7_75t_L g4219 ( 
.A(n_2561),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_2926),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_3307),
.Y(n_4221)
);

BUFx2_ASAP7_75t_L g4222 ( 
.A(n_3849),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_2926),
.Y(n_4223)
);

BUFx6f_ASAP7_75t_L g4224 ( 
.A(n_2926),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3017),
.Y(n_4225)
);

CKINVDCx5p33_ASAP7_75t_R g4226 ( 
.A(n_2572),
.Y(n_4226)
);

CKINVDCx20_ASAP7_75t_R g4227 ( 
.A(n_2648),
.Y(n_4227)
);

CKINVDCx5p33_ASAP7_75t_R g4228 ( 
.A(n_2573),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3017),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3017),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3077),
.Y(n_4231)
);

CKINVDCx20_ASAP7_75t_R g4232 ( 
.A(n_2658),
.Y(n_4232)
);

BUFx2_ASAP7_75t_L g4233 ( 
.A(n_3865),
.Y(n_4233)
);

CKINVDCx5p33_ASAP7_75t_R g4234 ( 
.A(n_2575),
.Y(n_4234)
);

CKINVDCx5p33_ASAP7_75t_R g4235 ( 
.A(n_2576),
.Y(n_4235)
);

CKINVDCx5p33_ASAP7_75t_R g4236 ( 
.A(n_2577),
.Y(n_4236)
);

CKINVDCx20_ASAP7_75t_R g4237 ( 
.A(n_2663),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3077),
.Y(n_4238)
);

CKINVDCx5p33_ASAP7_75t_R g4239 ( 
.A(n_2579),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_3077),
.Y(n_4240)
);

INVx1_ASAP7_75t_SL g4241 ( 
.A(n_3873),
.Y(n_4241)
);

CKINVDCx5p33_ASAP7_75t_R g4242 ( 
.A(n_2580),
.Y(n_4242)
);

BUFx3_ASAP7_75t_L g4243 ( 
.A(n_2713),
.Y(n_4243)
);

NOR2xp67_ASAP7_75t_L g4244 ( 
.A(n_3638),
.B(n_1),
.Y(n_4244)
);

NOR2xp67_ASAP7_75t_L g4245 ( 
.A(n_3118),
.B(n_1),
.Y(n_4245)
);

BUFx3_ASAP7_75t_L g4246 ( 
.A(n_2819),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_3080),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_3080),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_3080),
.Y(n_4249)
);

HB1xp67_ASAP7_75t_L g4250 ( 
.A(n_4045),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_3154),
.Y(n_4251)
);

HB1xp67_ASAP7_75t_L g4252 ( 
.A(n_2750),
.Y(n_4252)
);

CKINVDCx5p33_ASAP7_75t_R g4253 ( 
.A(n_2581),
.Y(n_4253)
);

CKINVDCx20_ASAP7_75t_R g4254 ( 
.A(n_2668),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_3307),
.Y(n_4255)
);

CKINVDCx5p33_ASAP7_75t_R g4256 ( 
.A(n_2585),
.Y(n_4256)
);

HB1xp67_ASAP7_75t_L g4257 ( 
.A(n_2816),
.Y(n_4257)
);

CKINVDCx5p33_ASAP7_75t_R g4258 ( 
.A(n_2587),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_3154),
.Y(n_4259)
);

CKINVDCx5p33_ASAP7_75t_R g4260 ( 
.A(n_2588),
.Y(n_4260)
);

CKINVDCx5p33_ASAP7_75t_R g4261 ( 
.A(n_2589),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_3154),
.Y(n_4262)
);

CKINVDCx20_ASAP7_75t_R g4263 ( 
.A(n_2679),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3251),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3251),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_3307),
.Y(n_4266)
);

BUFx2_ASAP7_75t_R g4267 ( 
.A(n_2591),
.Y(n_4267)
);

CKINVDCx5p33_ASAP7_75t_R g4268 ( 
.A(n_2593),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_3251),
.Y(n_4269)
);

BUFx3_ASAP7_75t_L g4270 ( 
.A(n_2863),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_3300),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_3300),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_3300),
.Y(n_4273)
);

CKINVDCx5p33_ASAP7_75t_R g4274 ( 
.A(n_2595),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_3359),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3359),
.Y(n_4276)
);

CKINVDCx5p33_ASAP7_75t_R g4277 ( 
.A(n_2597),
.Y(n_4277)
);

CKINVDCx5p33_ASAP7_75t_R g4278 ( 
.A(n_2600),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_3359),
.Y(n_4279)
);

CKINVDCx5p33_ASAP7_75t_R g4280 ( 
.A(n_2601),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_3384),
.Y(n_4281)
);

CKINVDCx20_ASAP7_75t_R g4282 ( 
.A(n_2684),
.Y(n_4282)
);

CKINVDCx5p33_ASAP7_75t_R g4283 ( 
.A(n_2603),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3384),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_3384),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_3442),
.Y(n_4286)
);

CKINVDCx20_ASAP7_75t_R g4287 ( 
.A(n_2727),
.Y(n_4287)
);

CKINVDCx5p33_ASAP7_75t_R g4288 ( 
.A(n_2608),
.Y(n_4288)
);

INVx2_ASAP7_75t_L g4289 ( 
.A(n_3442),
.Y(n_4289)
);

BUFx2_ASAP7_75t_L g4290 ( 
.A(n_2835),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_3442),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_3589),
.Y(n_4292)
);

CKINVDCx5p33_ASAP7_75t_R g4293 ( 
.A(n_2609),
.Y(n_4293)
);

BUFx6f_ASAP7_75t_L g4294 ( 
.A(n_3589),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_3589),
.Y(n_4295)
);

CKINVDCx20_ASAP7_75t_R g4296 ( 
.A(n_2740),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_3591),
.Y(n_4297)
);

CKINVDCx20_ASAP7_75t_R g4298 ( 
.A(n_2747),
.Y(n_4298)
);

CKINVDCx5p33_ASAP7_75t_R g4299 ( 
.A(n_2610),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_3591),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_3591),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_3600),
.Y(n_4302)
);

CKINVDCx5p33_ASAP7_75t_R g4303 ( 
.A(n_2612),
.Y(n_4303)
);

CKINVDCx5p33_ASAP7_75t_R g4304 ( 
.A(n_2613),
.Y(n_4304)
);

INVx2_ASAP7_75t_L g4305 ( 
.A(n_3600),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3600),
.Y(n_4306)
);

INVx1_ASAP7_75t_SL g4307 ( 
.A(n_2582),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_3618),
.Y(n_4308)
);

CKINVDCx5p33_ASAP7_75t_R g4309 ( 
.A(n_2615),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_3618),
.Y(n_4310)
);

CKINVDCx14_ASAP7_75t_R g4311 ( 
.A(n_2657),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3618),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_3649),
.Y(n_4313)
);

BUFx2_ASAP7_75t_L g4314 ( 
.A(n_2918),
.Y(n_4314)
);

CKINVDCx5p33_ASAP7_75t_R g4315 ( 
.A(n_2617),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_3649),
.Y(n_4316)
);

INVxp67_ASAP7_75t_L g4317 ( 
.A(n_2985),
.Y(n_4317)
);

CKINVDCx20_ASAP7_75t_R g4318 ( 
.A(n_2793),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_3649),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_3798),
.Y(n_4320)
);

BUFx6f_ASAP7_75t_L g4321 ( 
.A(n_3798),
.Y(n_4321)
);

CKINVDCx5p33_ASAP7_75t_R g4322 ( 
.A(n_2620),
.Y(n_4322)
);

CKINVDCx5p33_ASAP7_75t_R g4323 ( 
.A(n_2621),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_3798),
.Y(n_4324)
);

CKINVDCx5p33_ASAP7_75t_R g4325 ( 
.A(n_2622),
.Y(n_4325)
);

CKINVDCx16_ASAP7_75t_R g4326 ( 
.A(n_2657),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_3800),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_3800),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_3800),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3812),
.Y(n_4330)
);

CKINVDCx5p33_ASAP7_75t_R g4331 ( 
.A(n_2624),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_3812),
.Y(n_4332)
);

CKINVDCx5p33_ASAP7_75t_R g4333 ( 
.A(n_2625),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_3812),
.Y(n_4334)
);

CKINVDCx5p33_ASAP7_75t_R g4335 ( 
.A(n_2627),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_3821),
.Y(n_4336)
);

CKINVDCx5p33_ASAP7_75t_R g4337 ( 
.A(n_2628),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_3821),
.Y(n_4338)
);

CKINVDCx5p33_ASAP7_75t_R g4339 ( 
.A(n_2630),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_3821),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_3766),
.B(n_2),
.Y(n_4341)
);

CKINVDCx5p33_ASAP7_75t_R g4342 ( 
.A(n_2631),
.Y(n_4342)
);

CKINVDCx5p33_ASAP7_75t_R g4343 ( 
.A(n_2636),
.Y(n_4343)
);

CKINVDCx5p33_ASAP7_75t_R g4344 ( 
.A(n_2637),
.Y(n_4344)
);

CKINVDCx20_ASAP7_75t_R g4345 ( 
.A(n_2810),
.Y(n_4345)
);

BUFx6f_ASAP7_75t_L g4346 ( 
.A(n_3989),
.Y(n_4346)
);

INVxp67_ASAP7_75t_SL g4347 ( 
.A(n_3989),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_3989),
.Y(n_4348)
);

CKINVDCx5p33_ASAP7_75t_R g4349 ( 
.A(n_2640),
.Y(n_4349)
);

INVx3_ASAP7_75t_L g4350 ( 
.A(n_2731),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4027),
.Y(n_4351)
);

BUFx3_ASAP7_75t_L g4352 ( 
.A(n_2871),
.Y(n_4352)
);

BUFx3_ASAP7_75t_L g4353 ( 
.A(n_2966),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4027),
.Y(n_4354)
);

NOR2xp33_ASAP7_75t_L g4355 ( 
.A(n_3907),
.B(n_2),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_4027),
.Y(n_4356)
);

CKINVDCx5p33_ASAP7_75t_R g4357 ( 
.A(n_2643),
.Y(n_4357)
);

BUFx3_ASAP7_75t_L g4358 ( 
.A(n_2968),
.Y(n_4358)
);

CKINVDCx5p33_ASAP7_75t_R g4359 ( 
.A(n_2644),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_2979),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_3002),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_3014),
.Y(n_4362)
);

HB1xp67_ASAP7_75t_L g4363 ( 
.A(n_3149),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_3034),
.Y(n_4364)
);

BUFx3_ASAP7_75t_L g4365 ( 
.A(n_3137),
.Y(n_4365)
);

INVx2_ASAP7_75t_SL g4366 ( 
.A(n_2730),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_3165),
.Y(n_4367)
);

BUFx3_ASAP7_75t_L g4368 ( 
.A(n_3166),
.Y(n_4368)
);

CKINVDCx5p33_ASAP7_75t_R g4369 ( 
.A(n_2645),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_3195),
.Y(n_4370)
);

CKINVDCx5p33_ASAP7_75t_R g4371 ( 
.A(n_2646),
.Y(n_4371)
);

CKINVDCx5p33_ASAP7_75t_R g4372 ( 
.A(n_2649),
.Y(n_4372)
);

INVx1_ASAP7_75t_SL g4373 ( 
.A(n_2639),
.Y(n_4373)
);

CKINVDCx16_ASAP7_75t_R g4374 ( 
.A(n_2730),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_3217),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_3237),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_3243),
.Y(n_4377)
);

NOR2xp67_ASAP7_75t_L g4378 ( 
.A(n_2569),
.B(n_2),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_3244),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_3313),
.Y(n_4380)
);

CKINVDCx5p33_ASAP7_75t_R g4381 ( 
.A(n_2650),
.Y(n_4381)
);

CKINVDCx5p33_ASAP7_75t_R g4382 ( 
.A(n_2651),
.Y(n_4382)
);

INVx2_ASAP7_75t_SL g4383 ( 
.A(n_2763),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_3314),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_3340),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_3375),
.Y(n_4386)
);

BUFx6f_ASAP7_75t_L g4387 ( 
.A(n_2731),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_3411),
.Y(n_4388)
);

CKINVDCx5p33_ASAP7_75t_R g4389 ( 
.A(n_2652),
.Y(n_4389)
);

CKINVDCx20_ASAP7_75t_R g4390 ( 
.A(n_2853),
.Y(n_4390)
);

INVx2_ASAP7_75t_SL g4391 ( 
.A(n_2763),
.Y(n_4391)
);

CKINVDCx5p33_ASAP7_75t_R g4392 ( 
.A(n_2653),
.Y(n_4392)
);

CKINVDCx5p33_ASAP7_75t_R g4393 ( 
.A(n_2654),
.Y(n_4393)
);

CKINVDCx5p33_ASAP7_75t_R g4394 ( 
.A(n_2656),
.Y(n_4394)
);

CKINVDCx5p33_ASAP7_75t_R g4395 ( 
.A(n_2661),
.Y(n_4395)
);

CKINVDCx5p33_ASAP7_75t_R g4396 ( 
.A(n_2664),
.Y(n_4396)
);

CKINVDCx16_ASAP7_75t_R g4397 ( 
.A(n_2823),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_3520),
.Y(n_4398)
);

BUFx2_ASAP7_75t_L g4399 ( 
.A(n_3199),
.Y(n_4399)
);

CKINVDCx5p33_ASAP7_75t_R g4400 ( 
.A(n_2665),
.Y(n_4400)
);

BUFx3_ASAP7_75t_L g4401 ( 
.A(n_3545),
.Y(n_4401)
);

CKINVDCx5p33_ASAP7_75t_R g4402 ( 
.A(n_2666),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_3557),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_3621),
.Y(n_4404)
);

CKINVDCx20_ASAP7_75t_R g4405 ( 
.A(n_2855),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_3655),
.Y(n_4406)
);

CKINVDCx20_ASAP7_75t_R g4407 ( 
.A(n_2861),
.Y(n_4407)
);

CKINVDCx5p33_ASAP7_75t_R g4408 ( 
.A(n_2670),
.Y(n_4408)
);

CKINVDCx5p33_ASAP7_75t_R g4409 ( 
.A(n_2672),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_3691),
.Y(n_4410)
);

CKINVDCx5p33_ASAP7_75t_R g4411 ( 
.A(n_2673),
.Y(n_4411)
);

CKINVDCx20_ASAP7_75t_R g4412 ( 
.A(n_2882),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_3696),
.Y(n_4413)
);

INVx2_ASAP7_75t_SL g4414 ( 
.A(n_2823),
.Y(n_4414)
);

CKINVDCx5p33_ASAP7_75t_R g4415 ( 
.A(n_2674),
.Y(n_4415)
);

CKINVDCx5p33_ASAP7_75t_R g4416 ( 
.A(n_2680),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4001),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4012),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4015),
.Y(n_4419)
);

INVx2_ASAP7_75t_L g4420 ( 
.A(n_2574),
.Y(n_4420)
);

CKINVDCx5p33_ASAP7_75t_R g4421 ( 
.A(n_2681),
.Y(n_4421)
);

HB1xp67_ASAP7_75t_L g4422 ( 
.A(n_3221),
.Y(n_4422)
);

CKINVDCx5p33_ASAP7_75t_R g4423 ( 
.A(n_2682),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_2946),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_3001),
.Y(n_4425)
);

CKINVDCx5p33_ASAP7_75t_R g4426 ( 
.A(n_2686),
.Y(n_4426)
);

CKINVDCx5p33_ASAP7_75t_R g4427 ( 
.A(n_2689),
.Y(n_4427)
);

INVx2_ASAP7_75t_L g4428 ( 
.A(n_2578),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_2584),
.Y(n_4429)
);

CKINVDCx20_ASAP7_75t_R g4430 ( 
.A(n_2930),
.Y(n_4430)
);

BUFx6f_ASAP7_75t_L g4431 ( 
.A(n_2731),
.Y(n_4431)
);

CKINVDCx5p33_ASAP7_75t_R g4432 ( 
.A(n_2691),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_3056),
.Y(n_4433)
);

CKINVDCx5p33_ASAP7_75t_R g4434 ( 
.A(n_2692),
.Y(n_4434)
);

CKINVDCx5p33_ASAP7_75t_R g4435 ( 
.A(n_2693),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_3253),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_3254),
.Y(n_4437)
);

CKINVDCx5p33_ASAP7_75t_R g4438 ( 
.A(n_2695),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_3355),
.Y(n_4439)
);

CKINVDCx5p33_ASAP7_75t_R g4440 ( 
.A(n_2696),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_3420),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_3539),
.Y(n_4442)
);

CKINVDCx5p33_ASAP7_75t_R g4443 ( 
.A(n_2697),
.Y(n_4443)
);

CKINVDCx5p33_ASAP7_75t_R g4444 ( 
.A(n_2698),
.Y(n_4444)
);

CKINVDCx5p33_ASAP7_75t_R g4445 ( 
.A(n_2699),
.Y(n_4445)
);

CKINVDCx5p33_ASAP7_75t_R g4446 ( 
.A(n_2701),
.Y(n_4446)
);

CKINVDCx5p33_ASAP7_75t_R g4447 ( 
.A(n_2703),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_3568),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_3736),
.Y(n_4449)
);

INVxp67_ASAP7_75t_L g4450 ( 
.A(n_3440),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_3805),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_3883),
.Y(n_4452)
);

BUFx6f_ASAP7_75t_L g4453 ( 
.A(n_3281),
.Y(n_4453)
);

BUFx10_ASAP7_75t_L g4454 ( 
.A(n_3281),
.Y(n_4454)
);

CKINVDCx5p33_ASAP7_75t_R g4455 ( 
.A(n_2706),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_3537),
.Y(n_4456)
);

INVxp33_ASAP7_75t_L g4457 ( 
.A(n_3586),
.Y(n_4457)
);

CKINVDCx5p33_ASAP7_75t_R g4458 ( 
.A(n_2707),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_3590),
.Y(n_4459)
);

INVx2_ASAP7_75t_SL g4460 ( 
.A(n_2880),
.Y(n_4460)
);

CKINVDCx14_ASAP7_75t_R g4461 ( 
.A(n_2880),
.Y(n_4461)
);

CKINVDCx16_ASAP7_75t_R g4462 ( 
.A(n_2954),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_3709),
.Y(n_4463)
);

CKINVDCx20_ASAP7_75t_R g4464 ( 
.A(n_2951),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_3837),
.Y(n_4465)
);

CKINVDCx5p33_ASAP7_75t_R g4466 ( 
.A(n_2709),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_2592),
.Y(n_4467)
);

CKINVDCx5p33_ASAP7_75t_R g4468 ( 
.A(n_2711),
.Y(n_4468)
);

INVx1_ASAP7_75t_L g4469 ( 
.A(n_3926),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_3965),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_3972),
.Y(n_4471)
);

BUFx6f_ASAP7_75t_L g4472 ( 
.A(n_3281),
.Y(n_4472)
);

BUFx2_ASAP7_75t_L g4473 ( 
.A(n_4031),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_2596),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4034),
.Y(n_4475)
);

CKINVDCx5p33_ASAP7_75t_R g4476 ( 
.A(n_2714),
.Y(n_4476)
);

BUFx8_ASAP7_75t_SL g4477 ( 
.A(n_4038),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_2599),
.Y(n_4478)
);

CKINVDCx16_ASAP7_75t_R g4479 ( 
.A(n_2954),
.Y(n_4479)
);

CKINVDCx5p33_ASAP7_75t_R g4480 ( 
.A(n_2715),
.Y(n_4480)
);

CKINVDCx5p33_ASAP7_75t_R g4481 ( 
.A(n_2717),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_2605),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4044),
.Y(n_4483)
);

CKINVDCx5p33_ASAP7_75t_R g4484 ( 
.A(n_2718),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4046),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_2619),
.Y(n_4486)
);

INVxp33_ASAP7_75t_SL g4487 ( 
.A(n_2850),
.Y(n_4487)
);

INVxp67_ASAP7_75t_SL g4488 ( 
.A(n_2623),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4048),
.Y(n_4489)
);

CKINVDCx16_ASAP7_75t_R g4490 ( 
.A(n_3114),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4050),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4052),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4053),
.Y(n_4493)
);

CKINVDCx16_ASAP7_75t_R g4494 ( 
.A(n_3114),
.Y(n_4494)
);

BUFx2_ASAP7_75t_L g4495 ( 
.A(n_2956),
.Y(n_4495)
);

CKINVDCx5p33_ASAP7_75t_R g4496 ( 
.A(n_2725),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_2629),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_2632),
.Y(n_4498)
);

CKINVDCx5p33_ASAP7_75t_R g4499 ( 
.A(n_2726),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4033),
.Y(n_4500)
);

OR2x2_ASAP7_75t_L g4501 ( 
.A(n_2635),
.B(n_3),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4036),
.Y(n_4502)
);

CKINVDCx20_ASAP7_75t_R g4503 ( 
.A(n_2980),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_2642),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_2655),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_2659),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_2660),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_2667),
.Y(n_4508)
);

INVx2_ASAP7_75t_SL g4509 ( 
.A(n_3141),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_2669),
.Y(n_4510)
);

INVx1_ASAP7_75t_L g4511 ( 
.A(n_2675),
.Y(n_4511)
);

CKINVDCx5p33_ASAP7_75t_R g4512 ( 
.A(n_2728),
.Y(n_4512)
);

CKINVDCx5p33_ASAP7_75t_R g4513 ( 
.A(n_2736),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_2676),
.Y(n_4514)
);

NOR2xp33_ASAP7_75t_L g4515 ( 
.A(n_2798),
.B(n_3),
.Y(n_4515)
);

INVx2_ASAP7_75t_L g4516 ( 
.A(n_2677),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_2678),
.Y(n_4517)
);

CKINVDCx5p33_ASAP7_75t_R g4518 ( 
.A(n_2738),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_2685),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_2688),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_2690),
.Y(n_4521)
);

CKINVDCx5p33_ASAP7_75t_R g4522 ( 
.A(n_2745),
.Y(n_4522)
);

CKINVDCx5p33_ASAP7_75t_R g4523 ( 
.A(n_2749),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_2694),
.Y(n_4524)
);

CKINVDCx5p33_ASAP7_75t_R g4525 ( 
.A(n_2754),
.Y(n_4525)
);

CKINVDCx5p33_ASAP7_75t_R g4526 ( 
.A(n_2755),
.Y(n_4526)
);

CKINVDCx5p33_ASAP7_75t_R g4527 ( 
.A(n_2765),
.Y(n_4527)
);

INVx2_ASAP7_75t_SL g4528 ( 
.A(n_3141),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_2704),
.Y(n_4529)
);

INVx2_ASAP7_75t_L g4530 ( 
.A(n_2705),
.Y(n_4530)
);

CKINVDCx5p33_ASAP7_75t_R g4531 ( 
.A(n_2766),
.Y(n_4531)
);

CKINVDCx5p33_ASAP7_75t_R g4532 ( 
.A(n_2768),
.Y(n_4532)
);

INVxp67_ASAP7_75t_L g4533 ( 
.A(n_3148),
.Y(n_4533)
);

CKINVDCx5p33_ASAP7_75t_R g4534 ( 
.A(n_2770),
.Y(n_4534)
);

BUFx3_ASAP7_75t_L g4535 ( 
.A(n_2708),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_2710),
.Y(n_4536)
);

INVx1_ASAP7_75t_SL g4537 ( 
.A(n_2662),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_2716),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_2719),
.Y(n_4539)
);

CKINVDCx5p33_ASAP7_75t_R g4540 ( 
.A(n_2772),
.Y(n_4540)
);

CKINVDCx5p33_ASAP7_75t_R g4541 ( 
.A(n_2773),
.Y(n_4541)
);

BUFx6f_ASAP7_75t_L g4542 ( 
.A(n_2607),
.Y(n_4542)
);

CKINVDCx5p33_ASAP7_75t_R g4543 ( 
.A(n_2775),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_2721),
.Y(n_4544)
);

INVx1_ASAP7_75t_L g4545 ( 
.A(n_2723),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_2724),
.Y(n_4546)
);

BUFx2_ASAP7_75t_L g4547 ( 
.A(n_3036),
.Y(n_4547)
);

CKINVDCx5p33_ASAP7_75t_R g4548 ( 
.A(n_2776),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_2732),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_2739),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_2741),
.Y(n_4551)
);

CKINVDCx5p33_ASAP7_75t_R g4552 ( 
.A(n_2777),
.Y(n_4552)
);

NOR2xp33_ASAP7_75t_R g4553 ( 
.A(n_4032),
.B(n_2779),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_2742),
.Y(n_4554)
);

CKINVDCx5p33_ASAP7_75t_R g4555 ( 
.A(n_2780),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_2743),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_2744),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_2746),
.Y(n_4558)
);

CKINVDCx6p67_ASAP7_75t_R g4559 ( 
.A(n_3148),
.Y(n_4559)
);

CKINVDCx5p33_ASAP7_75t_R g4560 ( 
.A(n_2783),
.Y(n_4560)
);

BUFx2_ASAP7_75t_L g4561 ( 
.A(n_3041),
.Y(n_4561)
);

CKINVDCx5p33_ASAP7_75t_R g4562 ( 
.A(n_2785),
.Y(n_4562)
);

BUFx2_ASAP7_75t_L g4563 ( 
.A(n_3047),
.Y(n_4563)
);

CKINVDCx5p33_ASAP7_75t_R g4564 ( 
.A(n_2786),
.Y(n_4564)
);

CKINVDCx5p33_ASAP7_75t_R g4565 ( 
.A(n_2787),
.Y(n_4565)
);

CKINVDCx5p33_ASAP7_75t_R g4566 ( 
.A(n_2788),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_2748),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_2752),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_2757),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_2758),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_2759),
.Y(n_4571)
);

CKINVDCx5p33_ASAP7_75t_R g4572 ( 
.A(n_2790),
.Y(n_4572)
);

CKINVDCx5p33_ASAP7_75t_R g4573 ( 
.A(n_2796),
.Y(n_4573)
);

BUFx3_ASAP7_75t_L g4574 ( 
.A(n_2760),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_2762),
.Y(n_4575)
);

CKINVDCx5p33_ASAP7_75t_R g4576 ( 
.A(n_2797),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_2764),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_2771),
.Y(n_4578)
);

CKINVDCx16_ASAP7_75t_R g4579 ( 
.A(n_3153),
.Y(n_4579)
);

CKINVDCx16_ASAP7_75t_R g4580 ( 
.A(n_3153),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_2774),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_2778),
.Y(n_4582)
);

CKINVDCx5p33_ASAP7_75t_R g4583 ( 
.A(n_2801),
.Y(n_4583)
);

INVx2_ASAP7_75t_L g4584 ( 
.A(n_2784),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_2789),
.Y(n_4585)
);

CKINVDCx5p33_ASAP7_75t_R g4586 ( 
.A(n_2803),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_2794),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_2795),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_2799),
.Y(n_4589)
);

CKINVDCx5p33_ASAP7_75t_R g4590 ( 
.A(n_2804),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_2800),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_2802),
.Y(n_4592)
);

BUFx3_ASAP7_75t_L g4593 ( 
.A(n_2806),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_2808),
.Y(n_4594)
);

INVx2_ASAP7_75t_L g4595 ( 
.A(n_2813),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_2815),
.Y(n_4596)
);

CKINVDCx5p33_ASAP7_75t_R g4597 ( 
.A(n_2807),
.Y(n_4597)
);

CKINVDCx20_ASAP7_75t_R g4598 ( 
.A(n_3073),
.Y(n_4598)
);

OR2x2_ASAP7_75t_L g4599 ( 
.A(n_2818),
.B(n_3),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_2821),
.Y(n_4600)
);

CKINVDCx20_ASAP7_75t_R g4601 ( 
.A(n_3096),
.Y(n_4601)
);

CKINVDCx5p33_ASAP7_75t_R g4602 ( 
.A(n_2809),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_2826),
.Y(n_4603)
);

CKINVDCx5p33_ASAP7_75t_R g4604 ( 
.A(n_2811),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_2827),
.Y(n_4605)
);

CKINVDCx20_ASAP7_75t_R g4606 ( 
.A(n_3163),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_2830),
.Y(n_4607)
);

CKINVDCx5p33_ASAP7_75t_R g4608 ( 
.A(n_2812),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_2836),
.Y(n_4609)
);

CKINVDCx5p33_ASAP7_75t_R g4610 ( 
.A(n_2814),
.Y(n_4610)
);

CKINVDCx5p33_ASAP7_75t_R g4611 ( 
.A(n_2817),
.Y(n_4611)
);

INVx2_ASAP7_75t_SL g4612 ( 
.A(n_3269),
.Y(n_4612)
);

CKINVDCx5p33_ASAP7_75t_R g4613 ( 
.A(n_2820),
.Y(n_4613)
);

CKINVDCx5p33_ASAP7_75t_R g4614 ( 
.A(n_2822),
.Y(n_4614)
);

INVx1_ASAP7_75t_SL g4615 ( 
.A(n_2683),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_2837),
.Y(n_4616)
);

BUFx10_ASAP7_75t_L g4617 ( 
.A(n_2890),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_2846),
.Y(n_4618)
);

CKINVDCx5p33_ASAP7_75t_R g4619 ( 
.A(n_2824),
.Y(n_4619)
);

HB1xp67_ASAP7_75t_L g4620 ( 
.A(n_2825),
.Y(n_4620)
);

CKINVDCx5p33_ASAP7_75t_R g4621 ( 
.A(n_2828),
.Y(n_4621)
);

OR2x2_ASAP7_75t_L g4622 ( 
.A(n_2852),
.B(n_4),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_2856),
.Y(n_4623)
);

CKINVDCx5p33_ASAP7_75t_R g4624 ( 
.A(n_2829),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_2865),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_2875),
.Y(n_4626)
);

CKINVDCx5p33_ASAP7_75t_R g4627 ( 
.A(n_2831),
.Y(n_4627)
);

BUFx6f_ASAP7_75t_L g4628 ( 
.A(n_2611),
.Y(n_4628)
);

CKINVDCx5p33_ASAP7_75t_R g4629 ( 
.A(n_2832),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_2877),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_2885),
.Y(n_4631)
);

INVxp67_ASAP7_75t_L g4632 ( 
.A(n_3269),
.Y(n_4632)
);

CKINVDCx20_ASAP7_75t_R g4633 ( 
.A(n_3177),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_2889),
.Y(n_4634)
);

BUFx2_ASAP7_75t_L g4635 ( 
.A(n_3178),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_2892),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_2895),
.Y(n_4637)
);

CKINVDCx5p33_ASAP7_75t_R g4638 ( 
.A(n_2833),
.Y(n_4638)
);

CKINVDCx5p33_ASAP7_75t_R g4639 ( 
.A(n_2834),
.Y(n_4639)
);

CKINVDCx5p33_ASAP7_75t_R g4640 ( 
.A(n_2838),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_2897),
.Y(n_4641)
);

INVxp33_ASAP7_75t_L g4642 ( 
.A(n_2616),
.Y(n_4642)
);

INVx1_ASAP7_75t_SL g4643 ( 
.A(n_2733),
.Y(n_4643)
);

INVx1_ASAP7_75t_SL g4644 ( 
.A(n_2735),
.Y(n_4644)
);

BUFx6f_ASAP7_75t_L g4645 ( 
.A(n_2638),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_2898),
.Y(n_4646)
);

CKINVDCx5p33_ASAP7_75t_R g4647 ( 
.A(n_2839),
.Y(n_4647)
);

XNOR2xp5_ASAP7_75t_L g4648 ( 
.A(n_3235),
.B(n_4),
.Y(n_4648)
);

CKINVDCx5p33_ASAP7_75t_R g4649 ( 
.A(n_2840),
.Y(n_4649)
);

CKINVDCx20_ASAP7_75t_R g4650 ( 
.A(n_3236),
.Y(n_4650)
);

BUFx5_ASAP7_75t_L g4651 ( 
.A(n_2899),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_2900),
.Y(n_4652)
);

CKINVDCx5p33_ASAP7_75t_R g4653 ( 
.A(n_2842),
.Y(n_4653)
);

CKINVDCx5p33_ASAP7_75t_R g4654 ( 
.A(n_2843),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_2901),
.Y(n_4655)
);

CKINVDCx5p33_ASAP7_75t_R g4656 ( 
.A(n_2844),
.Y(n_4656)
);

CKINVDCx5p33_ASAP7_75t_R g4657 ( 
.A(n_2845),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_2903),
.Y(n_4658)
);

CKINVDCx5p33_ASAP7_75t_R g4659 ( 
.A(n_2847),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_2905),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_2916),
.Y(n_4661)
);

CKINVDCx5p33_ASAP7_75t_R g4662 ( 
.A(n_2848),
.Y(n_4662)
);

CKINVDCx5p33_ASAP7_75t_R g4663 ( 
.A(n_2849),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_2924),
.Y(n_4664)
);

CKINVDCx5p33_ASAP7_75t_R g4665 ( 
.A(n_2851),
.Y(n_4665)
);

CKINVDCx5p33_ASAP7_75t_R g4666 ( 
.A(n_2854),
.Y(n_4666)
);

CKINVDCx5p33_ASAP7_75t_R g4667 ( 
.A(n_2857),
.Y(n_4667)
);

CKINVDCx5p33_ASAP7_75t_R g4668 ( 
.A(n_2858),
.Y(n_4668)
);

CKINVDCx5p33_ASAP7_75t_R g4669 ( 
.A(n_2859),
.Y(n_4669)
);

INVxp67_ASAP7_75t_L g4670 ( 
.A(n_3276),
.Y(n_4670)
);

INVx1_ASAP7_75t_SL g4671 ( 
.A(n_2751),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_2928),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_2932),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_2938),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_2940),
.Y(n_4675)
);

INVxp33_ASAP7_75t_L g4676 ( 
.A(n_2647),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_2941),
.Y(n_4677)
);

CKINVDCx5p33_ASAP7_75t_R g4678 ( 
.A(n_2860),
.Y(n_4678)
);

INVxp67_ASAP7_75t_L g4679 ( 
.A(n_3276),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_2945),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_2948),
.Y(n_4681)
);

BUFx3_ASAP7_75t_L g4682 ( 
.A(n_2952),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_2955),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_2960),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_2962),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_2964),
.Y(n_4686)
);

BUFx3_ASAP7_75t_L g4687 ( 
.A(n_2965),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_2969),
.Y(n_4688)
);

HB1xp67_ASAP7_75t_L g4689 ( 
.A(n_2862),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_2970),
.Y(n_4690)
);

INVx1_ASAP7_75t_SL g4691 ( 
.A(n_2753),
.Y(n_4691)
);

CKINVDCx5p33_ASAP7_75t_R g4692 ( 
.A(n_2864),
.Y(n_4692)
);

INVx1_ASAP7_75t_SL g4693 ( 
.A(n_2963),
.Y(n_4693)
);

BUFx10_ASAP7_75t_L g4694 ( 
.A(n_2904),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_2978),
.Y(n_4695)
);

CKINVDCx5p33_ASAP7_75t_R g4696 ( 
.A(n_2866),
.Y(n_4696)
);

CKINVDCx5p33_ASAP7_75t_R g4697 ( 
.A(n_2867),
.Y(n_4697)
);

CKINVDCx16_ASAP7_75t_R g4698 ( 
.A(n_3283),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_2988),
.Y(n_4699)
);

BUFx3_ASAP7_75t_L g4700 ( 
.A(n_2991),
.Y(n_4700)
);

INVx1_ASAP7_75t_SL g4701 ( 
.A(n_2977),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_2999),
.Y(n_4702)
);

BUFx6f_ASAP7_75t_L g4703 ( 
.A(n_2671),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_3005),
.Y(n_4704)
);

CKINVDCx5p33_ASAP7_75t_R g4705 ( 
.A(n_2868),
.Y(n_4705)
);

CKINVDCx20_ASAP7_75t_R g4706 ( 
.A(n_3257),
.Y(n_4706)
);

BUFx3_ASAP7_75t_L g4707 ( 
.A(n_3012),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_3021),
.Y(n_4708)
);

INVxp67_ASAP7_75t_SL g4709 ( 
.A(n_3026),
.Y(n_4709)
);

INVx1_ASAP7_75t_SL g4710 ( 
.A(n_2981),
.Y(n_4710)
);

CKINVDCx5p33_ASAP7_75t_R g4711 ( 
.A(n_2869),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_3027),
.Y(n_4712)
);

CKINVDCx5p33_ASAP7_75t_R g4713 ( 
.A(n_2872),
.Y(n_4713)
);

CKINVDCx5p33_ASAP7_75t_R g4714 ( 
.A(n_2874),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_3030),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4096),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4140),
.Y(n_4717)
);

INVx1_ASAP7_75t_SL g4718 ( 
.A(n_4537),
.Y(n_4718)
);

CKINVDCx20_ASAP7_75t_R g4719 ( 
.A(n_4105),
.Y(n_4719)
);

CKINVDCx5p33_ASAP7_75t_R g4720 ( 
.A(n_4059),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4213),
.Y(n_4721)
);

INVxp67_ASAP7_75t_L g4722 ( 
.A(n_4307),
.Y(n_4722)
);

INVxp67_ASAP7_75t_SL g4723 ( 
.A(n_4347),
.Y(n_4723)
);

CKINVDCx5p33_ASAP7_75t_R g4724 ( 
.A(n_4060),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4075),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_4073),
.Y(n_4726)
);

CKINVDCx5p33_ASAP7_75t_R g4727 ( 
.A(n_4078),
.Y(n_4727)
);

CKINVDCx20_ASAP7_75t_R g4728 ( 
.A(n_4135),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4076),
.Y(n_4729)
);

CKINVDCx20_ASAP7_75t_R g4730 ( 
.A(n_4149),
.Y(n_4730)
);

CKINVDCx20_ASAP7_75t_R g4731 ( 
.A(n_4150),
.Y(n_4731)
);

INVxp67_ASAP7_75t_SL g4732 ( 
.A(n_4056),
.Y(n_4732)
);

INVxp67_ASAP7_75t_SL g4733 ( 
.A(n_4095),
.Y(n_4733)
);

INVx2_ASAP7_75t_L g4734 ( 
.A(n_4085),
.Y(n_4734)
);

CKINVDCx20_ASAP7_75t_R g4735 ( 
.A(n_4181),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4079),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4080),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4081),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4082),
.Y(n_4739)
);

CKINVDCx20_ASAP7_75t_R g4740 ( 
.A(n_4188),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4083),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4084),
.Y(n_4742)
);

CKINVDCx16_ASAP7_75t_R g4743 ( 
.A(n_4072),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4086),
.Y(n_4744)
);

CKINVDCx5p33_ASAP7_75t_R g4745 ( 
.A(n_4103),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4087),
.Y(n_4746)
);

CKINVDCx20_ASAP7_75t_R g4747 ( 
.A(n_4203),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4090),
.Y(n_4748)
);

BUFx6f_ASAP7_75t_L g4749 ( 
.A(n_4085),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4093),
.Y(n_4750)
);

CKINVDCx20_ASAP7_75t_R g4751 ( 
.A(n_4227),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4099),
.Y(n_4752)
);

CKINVDCx5p33_ASAP7_75t_R g4753 ( 
.A(n_4106),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4102),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4104),
.Y(n_4755)
);

CKINVDCx20_ASAP7_75t_R g4756 ( 
.A(n_4232),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_4085),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4112),
.Y(n_4758)
);

CKINVDCx16_ASAP7_75t_R g4759 ( 
.A(n_4074),
.Y(n_4759)
);

CKINVDCx20_ASAP7_75t_R g4760 ( 
.A(n_4237),
.Y(n_4760)
);

CKINVDCx5p33_ASAP7_75t_R g4761 ( 
.A(n_4108),
.Y(n_4761)
);

CKINVDCx20_ASAP7_75t_R g4762 ( 
.A(n_4254),
.Y(n_4762)
);

INVxp33_ASAP7_75t_L g4763 ( 
.A(n_4148),
.Y(n_4763)
);

CKINVDCx20_ASAP7_75t_R g4764 ( 
.A(n_4263),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4115),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4122),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4129),
.Y(n_4767)
);

INVxp67_ASAP7_75t_SL g4768 ( 
.A(n_4141),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4130),
.Y(n_4769)
);

INVxp33_ASAP7_75t_SL g4770 ( 
.A(n_4088),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4133),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4138),
.Y(n_4772)
);

CKINVDCx20_ASAP7_75t_R g4773 ( 
.A(n_4282),
.Y(n_4773)
);

CKINVDCx20_ASAP7_75t_R g4774 ( 
.A(n_4287),
.Y(n_4774)
);

INVxp67_ASAP7_75t_L g4775 ( 
.A(n_4373),
.Y(n_4775)
);

HB1xp67_ASAP7_75t_L g4776 ( 
.A(n_4176),
.Y(n_4776)
);

CKINVDCx5p33_ASAP7_75t_R g4777 ( 
.A(n_4109),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4142),
.Y(n_4778)
);

CKINVDCx16_ASAP7_75t_R g4779 ( 
.A(n_4098),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4143),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4144),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4145),
.Y(n_4782)
);

CKINVDCx5p33_ASAP7_75t_R g4783 ( 
.A(n_4110),
.Y(n_4783)
);

INVxp33_ASAP7_75t_L g4784 ( 
.A(n_4202),
.Y(n_4784)
);

CKINVDCx5p33_ASAP7_75t_R g4785 ( 
.A(n_4113),
.Y(n_4785)
);

INVxp33_ASAP7_75t_L g4786 ( 
.A(n_4250),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4146),
.Y(n_4787)
);

CKINVDCx16_ASAP7_75t_R g4788 ( 
.A(n_4111),
.Y(n_4788)
);

INVxp67_ASAP7_75t_L g4789 ( 
.A(n_4615),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4147),
.Y(n_4790)
);

CKINVDCx5p33_ASAP7_75t_R g4791 ( 
.A(n_4114),
.Y(n_4791)
);

CKINVDCx20_ASAP7_75t_R g4792 ( 
.A(n_4296),
.Y(n_4792)
);

CKINVDCx20_ASAP7_75t_R g4793 ( 
.A(n_4298),
.Y(n_4793)
);

INVx1_ASAP7_75t_SL g4794 ( 
.A(n_4643),
.Y(n_4794)
);

CKINVDCx5p33_ASAP7_75t_R g4795 ( 
.A(n_4116),
.Y(n_4795)
);

INVx2_ASAP7_75t_L g4796 ( 
.A(n_4089),
.Y(n_4796)
);

INVxp33_ASAP7_75t_L g4797 ( 
.A(n_4553),
.Y(n_4797)
);

CKINVDCx14_ASAP7_75t_R g4798 ( 
.A(n_4204),
.Y(n_4798)
);

INVxp67_ASAP7_75t_L g4799 ( 
.A(n_4644),
.Y(n_4799)
);

CKINVDCx16_ASAP7_75t_R g4800 ( 
.A(n_4118),
.Y(n_4800)
);

INVx2_ASAP7_75t_L g4801 ( 
.A(n_4089),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4089),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4151),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4091),
.Y(n_4804)
);

CKINVDCx5p33_ASAP7_75t_R g4805 ( 
.A(n_4117),
.Y(n_4805)
);

CKINVDCx5p33_ASAP7_75t_R g4806 ( 
.A(n_4119),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4154),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4156),
.Y(n_4808)
);

CKINVDCx5p33_ASAP7_75t_R g4809 ( 
.A(n_4121),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_4161),
.Y(n_4810)
);

CKINVDCx5p33_ASAP7_75t_R g4811 ( 
.A(n_4123),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4162),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4171),
.Y(n_4813)
);

CKINVDCx5p33_ASAP7_75t_R g4814 ( 
.A(n_4124),
.Y(n_4814)
);

INVxp33_ASAP7_75t_SL g4815 ( 
.A(n_4092),
.Y(n_4815)
);

INVxp33_ASAP7_75t_SL g4816 ( 
.A(n_4125),
.Y(n_4816)
);

INVx1_ASAP7_75t_SL g4817 ( 
.A(n_4671),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4177),
.Y(n_4818)
);

INVxp67_ASAP7_75t_L g4819 ( 
.A(n_4691),
.Y(n_4819)
);

CKINVDCx5p33_ASAP7_75t_R g4820 ( 
.A(n_4127),
.Y(n_4820)
);

CKINVDCx5p33_ASAP7_75t_R g4821 ( 
.A(n_4128),
.Y(n_4821)
);

HB1xp67_ASAP7_75t_L g4822 ( 
.A(n_4185),
.Y(n_4822)
);

CKINVDCx16_ASAP7_75t_R g4823 ( 
.A(n_4197),
.Y(n_4823)
);

INVxp67_ASAP7_75t_SL g4824 ( 
.A(n_4160),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4178),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4183),
.Y(n_4826)
);

INVxp67_ASAP7_75t_L g4827 ( 
.A(n_4693),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4190),
.Y(n_4828)
);

INVxp33_ASAP7_75t_SL g4829 ( 
.A(n_4132),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4191),
.Y(n_4830)
);

INVx2_ASAP7_75t_L g4831 ( 
.A(n_4091),
.Y(n_4831)
);

CKINVDCx20_ASAP7_75t_R g4832 ( 
.A(n_4318),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4057),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4058),
.Y(n_4834)
);

BUFx6f_ASAP7_75t_SL g4835 ( 
.A(n_4617),
.Y(n_4835)
);

CKINVDCx5p33_ASAP7_75t_R g4836 ( 
.A(n_4136),
.Y(n_4836)
);

INVxp67_ASAP7_75t_SL g4837 ( 
.A(n_4243),
.Y(n_4837)
);

BUFx6f_ASAP7_75t_SL g4838 ( 
.A(n_4617),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4062),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4063),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4065),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4066),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4067),
.Y(n_4843)
);

CKINVDCx20_ASAP7_75t_R g4844 ( 
.A(n_4345),
.Y(n_4844)
);

CKINVDCx5p33_ASAP7_75t_R g4845 ( 
.A(n_4137),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4068),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4070),
.Y(n_4847)
);

CKINVDCx5p33_ASAP7_75t_R g4848 ( 
.A(n_4152),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4192),
.Y(n_4849)
);

INVx2_ASAP7_75t_L g4850 ( 
.A(n_4091),
.Y(n_4850)
);

INVxp67_ASAP7_75t_L g4851 ( 
.A(n_4701),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4221),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4255),
.Y(n_4853)
);

CKINVDCx20_ASAP7_75t_R g4854 ( 
.A(n_4390),
.Y(n_4854)
);

CKINVDCx16_ASAP7_75t_R g4855 ( 
.A(n_4326),
.Y(n_4855)
);

CKINVDCx5p33_ASAP7_75t_R g4856 ( 
.A(n_4153),
.Y(n_4856)
);

BUFx3_ASAP7_75t_L g4857 ( 
.A(n_4454),
.Y(n_4857)
);

HB1xp67_ASAP7_75t_L g4858 ( 
.A(n_4218),
.Y(n_4858)
);

CKINVDCx16_ASAP7_75t_R g4859 ( 
.A(n_4374),
.Y(n_4859)
);

CKINVDCx5p33_ASAP7_75t_R g4860 ( 
.A(n_4155),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4266),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4077),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4094),
.Y(n_4863)
);

CKINVDCx5p33_ASAP7_75t_R g4864 ( 
.A(n_4158),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4107),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4184),
.Y(n_4866)
);

CKINVDCx5p33_ASAP7_75t_R g4867 ( 
.A(n_4163),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_4186),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4187),
.Y(n_4869)
);

INVxp67_ASAP7_75t_L g4870 ( 
.A(n_4710),
.Y(n_4870)
);

INVx1_ASAP7_75t_L g4871 ( 
.A(n_4482),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4483),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4485),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4489),
.Y(n_4874)
);

CKINVDCx20_ASAP7_75t_R g4875 ( 
.A(n_4405),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4491),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4492),
.Y(n_4877)
);

CKINVDCx16_ASAP7_75t_R g4878 ( 
.A(n_4397),
.Y(n_4878)
);

CKINVDCx5p33_ASAP7_75t_R g4879 ( 
.A(n_4164),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4159),
.Y(n_4880)
);

CKINVDCx20_ASAP7_75t_R g4881 ( 
.A(n_4407),
.Y(n_4881)
);

INVxp33_ASAP7_75t_L g4882 ( 
.A(n_4120),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4493),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4497),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4498),
.Y(n_4885)
);

INVxp33_ASAP7_75t_L g4886 ( 
.A(n_4134),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4500),
.Y(n_4887)
);

CKINVDCx20_ASAP7_75t_R g4888 ( 
.A(n_4412),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4502),
.Y(n_4889)
);

CKINVDCx5p33_ASAP7_75t_R g4890 ( 
.A(n_4165),
.Y(n_4890)
);

BUFx6f_ASAP7_75t_L g4891 ( 
.A(n_4159),
.Y(n_4891)
);

BUFx3_ASAP7_75t_L g4892 ( 
.A(n_4454),
.Y(n_4892)
);

CKINVDCx20_ASAP7_75t_R g4893 ( 
.A(n_4430),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4505),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4506),
.Y(n_4895)
);

CKINVDCx5p33_ASAP7_75t_R g4896 ( 
.A(n_4168),
.Y(n_4896)
);

INVxp33_ASAP7_75t_L g4897 ( 
.A(n_4170),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4507),
.Y(n_4898)
);

CKINVDCx20_ASAP7_75t_R g4899 ( 
.A(n_4464),
.Y(n_4899)
);

CKINVDCx5p33_ASAP7_75t_R g4900 ( 
.A(n_4172),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4508),
.Y(n_4901)
);

CKINVDCx16_ASAP7_75t_R g4902 ( 
.A(n_4462),
.Y(n_4902)
);

CKINVDCx5p33_ASAP7_75t_R g4903 ( 
.A(n_4175),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4510),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4511),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4514),
.Y(n_4906)
);

BUFx6f_ASAP7_75t_L g4907 ( 
.A(n_4159),
.Y(n_4907)
);

CKINVDCx5p33_ASAP7_75t_R g4908 ( 
.A(n_4179),
.Y(n_4908)
);

INVx2_ASAP7_75t_L g4909 ( 
.A(n_4166),
.Y(n_4909)
);

CKINVDCx5p33_ASAP7_75t_R g4910 ( 
.A(n_4180),
.Y(n_4910)
);

HB1xp67_ASAP7_75t_L g4911 ( 
.A(n_4241),
.Y(n_4911)
);

INVxp67_ASAP7_75t_SL g4912 ( 
.A(n_4246),
.Y(n_4912)
);

CKINVDCx20_ASAP7_75t_R g4913 ( 
.A(n_4503),
.Y(n_4913)
);

CKINVDCx20_ASAP7_75t_R g4914 ( 
.A(n_4598),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4517),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4519),
.Y(n_4916)
);

CKINVDCx20_ASAP7_75t_R g4917 ( 
.A(n_4601),
.Y(n_4917)
);

BUFx3_ASAP7_75t_L g4918 ( 
.A(n_4270),
.Y(n_4918)
);

CKINVDCx20_ASAP7_75t_R g4919 ( 
.A(n_4606),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4520),
.Y(n_4920)
);

INVxp33_ASAP7_75t_SL g4921 ( 
.A(n_4182),
.Y(n_4921)
);

INVxp33_ASAP7_75t_SL g4922 ( 
.A(n_4189),
.Y(n_4922)
);

CKINVDCx14_ASAP7_75t_R g4923 ( 
.A(n_4311),
.Y(n_4923)
);

INVxp67_ASAP7_75t_SL g4924 ( 
.A(n_4352),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4521),
.Y(n_4925)
);

CKINVDCx20_ASAP7_75t_R g4926 ( 
.A(n_4633),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4524),
.Y(n_4927)
);

INVxp67_ASAP7_75t_SL g4928 ( 
.A(n_4353),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4529),
.Y(n_4929)
);

HB1xp67_ASAP7_75t_L g4930 ( 
.A(n_4174),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4536),
.Y(n_4931)
);

CKINVDCx20_ASAP7_75t_R g4932 ( 
.A(n_4650),
.Y(n_4932)
);

INVxp67_ASAP7_75t_SL g4933 ( 
.A(n_4358),
.Y(n_4933)
);

CKINVDCx5p33_ASAP7_75t_R g4934 ( 
.A(n_4193),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4538),
.Y(n_4935)
);

INVxp67_ASAP7_75t_L g4936 ( 
.A(n_4620),
.Y(n_4936)
);

INVx1_ASAP7_75t_L g4937 ( 
.A(n_4544),
.Y(n_4937)
);

INVxp67_ASAP7_75t_SL g4938 ( 
.A(n_4365),
.Y(n_4938)
);

CKINVDCx20_ASAP7_75t_R g4939 ( 
.A(n_4706),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4545),
.Y(n_4940)
);

INVxp33_ASAP7_75t_SL g4941 ( 
.A(n_4195),
.Y(n_4941)
);

BUFx3_ASAP7_75t_L g4942 ( 
.A(n_4368),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_4546),
.Y(n_4943)
);

CKINVDCx14_ASAP7_75t_R g4944 ( 
.A(n_4461),
.Y(n_4944)
);

CKINVDCx5p33_ASAP7_75t_R g4945 ( 
.A(n_4199),
.Y(n_4945)
);

CKINVDCx5p33_ASAP7_75t_R g4946 ( 
.A(n_4205),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4549),
.Y(n_4947)
);

CKINVDCx20_ASAP7_75t_R g4948 ( 
.A(n_4479),
.Y(n_4948)
);

INVx2_ASAP7_75t_L g4949 ( 
.A(n_4166),
.Y(n_4949)
);

CKINVDCx5p33_ASAP7_75t_R g4950 ( 
.A(n_4207),
.Y(n_4950)
);

INVxp67_ASAP7_75t_SL g4951 ( 
.A(n_4401),
.Y(n_4951)
);

CKINVDCx16_ASAP7_75t_R g4952 ( 
.A(n_4490),
.Y(n_4952)
);

CKINVDCx20_ASAP7_75t_R g4953 ( 
.A(n_4494),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4550),
.Y(n_4954)
);

INVx1_ASAP7_75t_L g4955 ( 
.A(n_4551),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4554),
.Y(n_4956)
);

CKINVDCx5p33_ASAP7_75t_R g4957 ( 
.A(n_4208),
.Y(n_4957)
);

HB1xp67_ASAP7_75t_L g4958 ( 
.A(n_4222),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4556),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4557),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4558),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4567),
.Y(n_4962)
);

INVxp67_ASAP7_75t_L g4963 ( 
.A(n_4689),
.Y(n_4963)
);

CKINVDCx5p33_ASAP7_75t_R g4964 ( 
.A(n_4209),
.Y(n_4964)
);

CKINVDCx5p33_ASAP7_75t_R g4965 ( 
.A(n_4210),
.Y(n_4965)
);

HB1xp67_ASAP7_75t_L g4966 ( 
.A(n_4233),
.Y(n_4966)
);

CKINVDCx20_ASAP7_75t_R g4967 ( 
.A(n_4579),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4568),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4569),
.Y(n_4969)
);

INVxp67_ASAP7_75t_SL g4970 ( 
.A(n_4642),
.Y(n_4970)
);

INVx2_ASAP7_75t_L g4971 ( 
.A(n_4166),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4570),
.Y(n_4972)
);

CKINVDCx5p33_ASAP7_75t_R g4973 ( 
.A(n_4212),
.Y(n_4973)
);

CKINVDCx14_ASAP7_75t_R g4974 ( 
.A(n_4097),
.Y(n_4974)
);

INVx1_ASAP7_75t_SL g4975 ( 
.A(n_4215),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4571),
.Y(n_4976)
);

CKINVDCx20_ASAP7_75t_R g4977 ( 
.A(n_4580),
.Y(n_4977)
);

CKINVDCx5p33_ASAP7_75t_R g4978 ( 
.A(n_4226),
.Y(n_4978)
);

INVx1_ASAP7_75t_L g4979 ( 
.A(n_4575),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4577),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4578),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4581),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4582),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_4585),
.Y(n_4984)
);

CKINVDCx16_ASAP7_75t_R g4985 ( 
.A(n_4698),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4587),
.Y(n_4986)
);

CKINVDCx20_ASAP7_75t_R g4987 ( 
.A(n_4559),
.Y(n_4987)
);

CKINVDCx16_ASAP7_75t_R g4988 ( 
.A(n_4694),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4588),
.Y(n_4989)
);

CKINVDCx5p33_ASAP7_75t_R g4990 ( 
.A(n_4228),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4589),
.Y(n_4991)
);

CKINVDCx20_ASAP7_75t_R g4992 ( 
.A(n_4234),
.Y(n_4992)
);

BUFx3_ASAP7_75t_L g4993 ( 
.A(n_4384),
.Y(n_4993)
);

CKINVDCx16_ASAP7_75t_R g4994 ( 
.A(n_4694),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4592),
.Y(n_4995)
);

CKINVDCx16_ASAP7_75t_R g4996 ( 
.A(n_4495),
.Y(n_4996)
);

CKINVDCx5p33_ASAP7_75t_R g4997 ( 
.A(n_4235),
.Y(n_4997)
);

INVx2_ASAP7_75t_L g4998 ( 
.A(n_4167),
.Y(n_4998)
);

CKINVDCx5p33_ASAP7_75t_R g4999 ( 
.A(n_4236),
.Y(n_4999)
);

INVx2_ASAP7_75t_L g5000 ( 
.A(n_4167),
.Y(n_5000)
);

BUFx3_ASAP7_75t_L g5001 ( 
.A(n_4413),
.Y(n_5001)
);

INVx2_ASAP7_75t_L g5002 ( 
.A(n_4167),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4594),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_4596),
.Y(n_5004)
);

INVxp33_ASAP7_75t_L g5005 ( 
.A(n_4477),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4600),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4603),
.Y(n_5007)
);

CKINVDCx16_ASAP7_75t_R g5008 ( 
.A(n_4547),
.Y(n_5008)
);

CKINVDCx5p33_ASAP7_75t_R g5009 ( 
.A(n_4239),
.Y(n_5009)
);

HB1xp67_ASAP7_75t_L g5010 ( 
.A(n_4242),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4605),
.Y(n_5011)
);

INVxp33_ASAP7_75t_SL g5012 ( 
.A(n_4253),
.Y(n_5012)
);

INVx2_ASAP7_75t_L g5013 ( 
.A(n_4224),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4607),
.Y(n_5014)
);

CKINVDCx20_ASAP7_75t_R g5015 ( 
.A(n_4256),
.Y(n_5015)
);

INVxp33_ASAP7_75t_L g5016 ( 
.A(n_4561),
.Y(n_5016)
);

CKINVDCx20_ASAP7_75t_R g5017 ( 
.A(n_4258),
.Y(n_5017)
);

INVx2_ASAP7_75t_L g5018 ( 
.A(n_4224),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4609),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_4616),
.Y(n_5020)
);

INVxp33_ASAP7_75t_SL g5021 ( 
.A(n_4260),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4618),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4623),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4625),
.Y(n_5024)
);

INVx3_ASAP7_75t_L g5025 ( 
.A(n_4224),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4626),
.Y(n_5026)
);

INVx1_ASAP7_75t_SL g5027 ( 
.A(n_4261),
.Y(n_5027)
);

CKINVDCx5p33_ASAP7_75t_R g5028 ( 
.A(n_4268),
.Y(n_5028)
);

BUFx6f_ASAP7_75t_SL g5029 ( 
.A(n_4131),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4630),
.Y(n_5030)
);

CKINVDCx5p33_ASAP7_75t_R g5031 ( 
.A(n_4274),
.Y(n_5031)
);

CKINVDCx5p33_ASAP7_75t_R g5032 ( 
.A(n_4277),
.Y(n_5032)
);

INVx1_ASAP7_75t_L g5033 ( 
.A(n_4631),
.Y(n_5033)
);

CKINVDCx5p33_ASAP7_75t_R g5034 ( 
.A(n_4278),
.Y(n_5034)
);

BUFx2_ASAP7_75t_SL g5035 ( 
.A(n_4173),
.Y(n_5035)
);

HB1xp67_ASAP7_75t_L g5036 ( 
.A(n_4280),
.Y(n_5036)
);

INVx1_ASAP7_75t_L g5037 ( 
.A(n_4634),
.Y(n_5037)
);

INVxp67_ASAP7_75t_SL g5038 ( 
.A(n_4676),
.Y(n_5038)
);

INVx3_ASAP7_75t_L g5039 ( 
.A(n_4294),
.Y(n_5039)
);

HB1xp67_ASAP7_75t_L g5040 ( 
.A(n_4283),
.Y(n_5040)
);

CKINVDCx20_ASAP7_75t_R g5041 ( 
.A(n_4288),
.Y(n_5041)
);

INVx2_ASAP7_75t_L g5042 ( 
.A(n_4294),
.Y(n_5042)
);

CKINVDCx5p33_ASAP7_75t_R g5043 ( 
.A(n_4293),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4636),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4637),
.Y(n_5045)
);

CKINVDCx20_ASAP7_75t_R g5046 ( 
.A(n_4299),
.Y(n_5046)
);

CKINVDCx20_ASAP7_75t_R g5047 ( 
.A(n_4303),
.Y(n_5047)
);

BUFx2_ASAP7_75t_L g5048 ( 
.A(n_4304),
.Y(n_5048)
);

CKINVDCx20_ASAP7_75t_R g5049 ( 
.A(n_4309),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_4646),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4652),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_4655),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4658),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4660),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4661),
.Y(n_5055)
);

CKINVDCx5p33_ASAP7_75t_R g5056 ( 
.A(n_4315),
.Y(n_5056)
);

CKINVDCx20_ASAP7_75t_R g5057 ( 
.A(n_4322),
.Y(n_5057)
);

BUFx2_ASAP7_75t_L g5058 ( 
.A(n_4323),
.Y(n_5058)
);

INVxp67_ASAP7_75t_SL g5059 ( 
.A(n_4487),
.Y(n_5059)
);

INVx2_ASAP7_75t_L g5060 ( 
.A(n_4294),
.Y(n_5060)
);

INVx2_ASAP7_75t_L g5061 ( 
.A(n_4321),
.Y(n_5061)
);

CKINVDCx5p33_ASAP7_75t_R g5062 ( 
.A(n_4325),
.Y(n_5062)
);

INVx1_ASAP7_75t_L g5063 ( 
.A(n_4664),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4672),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4673),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4674),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_4675),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_4677),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_4681),
.Y(n_5069)
);

INVx1_ASAP7_75t_L g5070 ( 
.A(n_4683),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4684),
.Y(n_5071)
);

BUFx3_ASAP7_75t_L g5072 ( 
.A(n_4360),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_4686),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4688),
.Y(n_5074)
);

CKINVDCx20_ASAP7_75t_R g5075 ( 
.A(n_4331),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4690),
.Y(n_5076)
);

CKINVDCx20_ASAP7_75t_R g5077 ( 
.A(n_4333),
.Y(n_5077)
);

CKINVDCx5p33_ASAP7_75t_R g5078 ( 
.A(n_4335),
.Y(n_5078)
);

HB1xp67_ASAP7_75t_L g5079 ( 
.A(n_4337),
.Y(n_5079)
);

INVxp67_ASAP7_75t_L g5080 ( 
.A(n_4339),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_4695),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_4699),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_4702),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4704),
.Y(n_5084)
);

INVx1_ASAP7_75t_L g5085 ( 
.A(n_4708),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4712),
.Y(n_5086)
);

CKINVDCx5p33_ASAP7_75t_R g5087 ( 
.A(n_4342),
.Y(n_5087)
);

CKINVDCx5p33_ASAP7_75t_R g5088 ( 
.A(n_4343),
.Y(n_5088)
);

INVxp67_ASAP7_75t_SL g5089 ( 
.A(n_4321),
.Y(n_5089)
);

CKINVDCx5p33_ASAP7_75t_R g5090 ( 
.A(n_4344),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_4715),
.Y(n_5091)
);

BUFx6f_ASAP7_75t_L g5092 ( 
.A(n_4321),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4101),
.Y(n_5093)
);

CKINVDCx5p33_ASAP7_75t_R g5094 ( 
.A(n_4349),
.Y(n_5094)
);

CKINVDCx20_ASAP7_75t_R g5095 ( 
.A(n_4357),
.Y(n_5095)
);

HB1xp67_ASAP7_75t_L g5096 ( 
.A(n_4359),
.Y(n_5096)
);

BUFx2_ASAP7_75t_SL g5097 ( 
.A(n_4206),
.Y(n_5097)
);

INVxp67_ASAP7_75t_SL g5098 ( 
.A(n_4346),
.Y(n_5098)
);

CKINVDCx20_ASAP7_75t_R g5099 ( 
.A(n_4369),
.Y(n_5099)
);

INVxp67_ASAP7_75t_SL g5100 ( 
.A(n_4346),
.Y(n_5100)
);

CKINVDCx5p33_ASAP7_75t_R g5101 ( 
.A(n_4371),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_4488),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_4709),
.Y(n_5103)
);

CKINVDCx5p33_ASAP7_75t_R g5104 ( 
.A(n_4372),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_4064),
.Y(n_5105)
);

CKINVDCx16_ASAP7_75t_R g5106 ( 
.A(n_4563),
.Y(n_5106)
);

HB1xp67_ASAP7_75t_L g5107 ( 
.A(n_4381),
.Y(n_5107)
);

INVxp67_ASAP7_75t_SL g5108 ( 
.A(n_4346),
.Y(n_5108)
);

HB1xp67_ASAP7_75t_L g5109 ( 
.A(n_4382),
.Y(n_5109)
);

BUFx2_ASAP7_75t_L g5110 ( 
.A(n_4389),
.Y(n_5110)
);

CKINVDCx16_ASAP7_75t_R g5111 ( 
.A(n_4635),
.Y(n_5111)
);

CKINVDCx20_ASAP7_75t_R g5112 ( 
.A(n_4392),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4064),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_4064),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4064),
.Y(n_5115)
);

CKINVDCx5p33_ASAP7_75t_R g5116 ( 
.A(n_4393),
.Y(n_5116)
);

INVx1_ASAP7_75t_L g5117 ( 
.A(n_4064),
.Y(n_5117)
);

INVx1_ASAP7_75t_SL g5118 ( 
.A(n_4394),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4219),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_4219),
.Y(n_5120)
);

HB1xp67_ASAP7_75t_L g5121 ( 
.A(n_4395),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4219),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_4219),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_4219),
.Y(n_5124)
);

CKINVDCx5p33_ASAP7_75t_R g5125 ( 
.A(n_4396),
.Y(n_5125)
);

CKINVDCx5p33_ASAP7_75t_R g5126 ( 
.A(n_4400),
.Y(n_5126)
);

CKINVDCx5p33_ASAP7_75t_R g5127 ( 
.A(n_4402),
.Y(n_5127)
);

CKINVDCx5p33_ASAP7_75t_R g5128 ( 
.A(n_4408),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_4651),
.Y(n_5129)
);

INVxp67_ASAP7_75t_SL g5130 ( 
.A(n_4361),
.Y(n_5130)
);

INVxp67_ASAP7_75t_SL g5131 ( 
.A(n_4362),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_4651),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_4651),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_4651),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4651),
.Y(n_5135)
);

CKINVDCx5p33_ASAP7_75t_R g5136 ( 
.A(n_4409),
.Y(n_5136)
);

CKINVDCx5p33_ASAP7_75t_R g5137 ( 
.A(n_4411),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4364),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_4367),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_4370),
.Y(n_5140)
);

CKINVDCx16_ASAP7_75t_R g5141 ( 
.A(n_4252),
.Y(n_5141)
);

CKINVDCx20_ASAP7_75t_R g5142 ( 
.A(n_4415),
.Y(n_5142)
);

CKINVDCx5p33_ASAP7_75t_R g5143 ( 
.A(n_4416),
.Y(n_5143)
);

INVxp67_ASAP7_75t_SL g5144 ( 
.A(n_4375),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_4376),
.Y(n_5145)
);

INVxp33_ASAP7_75t_SL g5146 ( 
.A(n_4421),
.Y(n_5146)
);

INVxp33_ASAP7_75t_L g5147 ( 
.A(n_4457),
.Y(n_5147)
);

HB1xp67_ASAP7_75t_L g5148 ( 
.A(n_4423),
.Y(n_5148)
);

CKINVDCx5p33_ASAP7_75t_R g5149 ( 
.A(n_4426),
.Y(n_5149)
);

CKINVDCx20_ASAP7_75t_R g5150 ( 
.A(n_4427),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_4377),
.Y(n_5151)
);

INVxp67_ASAP7_75t_SL g5152 ( 
.A(n_4379),
.Y(n_5152)
);

CKINVDCx5p33_ASAP7_75t_R g5153 ( 
.A(n_4432),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_4380),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_4385),
.Y(n_5155)
);

CKINVDCx20_ASAP7_75t_R g5156 ( 
.A(n_4434),
.Y(n_5156)
);

BUFx6f_ASAP7_75t_L g5157 ( 
.A(n_4387),
.Y(n_5157)
);

INVxp67_ASAP7_75t_SL g5158 ( 
.A(n_4386),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_4388),
.Y(n_5159)
);

HB1xp67_ASAP7_75t_L g5160 ( 
.A(n_4435),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_4398),
.Y(n_5161)
);

INVx3_ASAP7_75t_L g5162 ( 
.A(n_4387),
.Y(n_5162)
);

BUFx3_ASAP7_75t_L g5163 ( 
.A(n_4403),
.Y(n_5163)
);

CKINVDCx5p33_ASAP7_75t_R g5164 ( 
.A(n_4438),
.Y(n_5164)
);

CKINVDCx5p33_ASAP7_75t_R g5165 ( 
.A(n_4440),
.Y(n_5165)
);

INVx2_ASAP7_75t_L g5166 ( 
.A(n_4387),
.Y(n_5166)
);

CKINVDCx20_ASAP7_75t_R g5167 ( 
.A(n_4443),
.Y(n_5167)
);

CKINVDCx5p33_ASAP7_75t_R g5168 ( 
.A(n_4444),
.Y(n_5168)
);

BUFx6f_ASAP7_75t_L g5169 ( 
.A(n_4431),
.Y(n_5169)
);

CKINVDCx5p33_ASAP7_75t_R g5170 ( 
.A(n_4445),
.Y(n_5170)
);

CKINVDCx5p33_ASAP7_75t_R g5171 ( 
.A(n_4446),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4404),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_4406),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_4410),
.Y(n_5174)
);

INVx1_ASAP7_75t_L g5175 ( 
.A(n_4417),
.Y(n_5175)
);

CKINVDCx20_ASAP7_75t_R g5176 ( 
.A(n_4447),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_4418),
.Y(n_5177)
);

CKINVDCx20_ASAP7_75t_R g5178 ( 
.A(n_4455),
.Y(n_5178)
);

INVxp67_ASAP7_75t_SL g5179 ( 
.A(n_4419),
.Y(n_5179)
);

CKINVDCx5p33_ASAP7_75t_R g5180 ( 
.A(n_4458),
.Y(n_5180)
);

CKINVDCx14_ASAP7_75t_R g5181 ( 
.A(n_4290),
.Y(n_5181)
);

INVxp33_ASAP7_75t_L g5182 ( 
.A(n_4257),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_4420),
.Y(n_5183)
);

HB1xp67_ASAP7_75t_L g5184 ( 
.A(n_4466),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_4428),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_4429),
.Y(n_5186)
);

CKINVDCx5p33_ASAP7_75t_R g5187 ( 
.A(n_4468),
.Y(n_5187)
);

INVxp33_ASAP7_75t_SL g5188 ( 
.A(n_4476),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_4467),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4474),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_4478),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_4486),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_4504),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_4516),
.Y(n_5194)
);

CKINVDCx5p33_ASAP7_75t_R g5195 ( 
.A(n_4480),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_4530),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_4539),
.Y(n_5197)
);

INVx2_ASAP7_75t_L g5198 ( 
.A(n_4431),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_4584),
.Y(n_5199)
);

INVxp33_ASAP7_75t_SL g5200 ( 
.A(n_4481),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_4591),
.Y(n_5201)
);

CKINVDCx5p33_ASAP7_75t_R g5202 ( 
.A(n_4484),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_4595),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_4641),
.Y(n_5204)
);

INVxp67_ASAP7_75t_SL g5205 ( 
.A(n_4350),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4680),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_4685),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_4350),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_4535),
.Y(n_5209)
);

CKINVDCx5p33_ASAP7_75t_R g5210 ( 
.A(n_4496),
.Y(n_5210)
);

INVxp67_ASAP7_75t_SL g5211 ( 
.A(n_4355),
.Y(n_5211)
);

CKINVDCx20_ASAP7_75t_R g5212 ( 
.A(n_4499),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_4431),
.Y(n_5213)
);

BUFx2_ASAP7_75t_L g5214 ( 
.A(n_4512),
.Y(n_5214)
);

INVxp67_ASAP7_75t_L g5215 ( 
.A(n_4513),
.Y(n_5215)
);

INVxp67_ASAP7_75t_SL g5216 ( 
.A(n_4453),
.Y(n_5216)
);

INVxp67_ASAP7_75t_SL g5217 ( 
.A(n_4453),
.Y(n_5217)
);

CKINVDCx5p33_ASAP7_75t_R g5218 ( 
.A(n_4518),
.Y(n_5218)
);

CKINVDCx5p33_ASAP7_75t_R g5219 ( 
.A(n_4522),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_4574),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_4593),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_4682),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_4687),
.Y(n_5223)
);

CKINVDCx5p33_ASAP7_75t_R g5224 ( 
.A(n_4523),
.Y(n_5224)
);

INVx1_ASAP7_75t_L g5225 ( 
.A(n_4700),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4707),
.Y(n_5226)
);

INVx1_ASAP7_75t_L g5227 ( 
.A(n_4285),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_4286),
.Y(n_5228)
);

CKINVDCx5p33_ASAP7_75t_R g5229 ( 
.A(n_4525),
.Y(n_5229)
);

CKINVDCx5p33_ASAP7_75t_R g5230 ( 
.A(n_4526),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_4289),
.Y(n_5231)
);

INVx1_ASAP7_75t_L g5232 ( 
.A(n_4301),
.Y(n_5232)
);

HB1xp67_ASAP7_75t_L g5233 ( 
.A(n_4527),
.Y(n_5233)
);

CKINVDCx5p33_ASAP7_75t_R g5234 ( 
.A(n_4531),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_4305),
.Y(n_5235)
);

BUFx6f_ASAP7_75t_L g5236 ( 
.A(n_4453),
.Y(n_5236)
);

CKINVDCx20_ASAP7_75t_R g5237 ( 
.A(n_4532),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_4313),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_4329),
.Y(n_5239)
);

CKINVDCx5p33_ASAP7_75t_R g5240 ( 
.A(n_4534),
.Y(n_5240)
);

INVx1_ASAP7_75t_L g5241 ( 
.A(n_4354),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_4472),
.Y(n_5242)
);

CKINVDCx20_ASAP7_75t_R g5243 ( 
.A(n_4540),
.Y(n_5243)
);

BUFx3_ASAP7_75t_L g5244 ( 
.A(n_4472),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_4356),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_4194),
.Y(n_5246)
);

INVxp67_ASAP7_75t_L g5247 ( 
.A(n_4541),
.Y(n_5247)
);

INVx2_ASAP7_75t_L g5248 ( 
.A(n_4472),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_4196),
.Y(n_5249)
);

INVxp67_ASAP7_75t_L g5250 ( 
.A(n_4543),
.Y(n_5250)
);

CKINVDCx5p33_ASAP7_75t_R g5251 ( 
.A(n_4548),
.Y(n_5251)
);

INVx2_ASAP7_75t_L g5252 ( 
.A(n_4542),
.Y(n_5252)
);

HB1xp67_ASAP7_75t_L g5253 ( 
.A(n_4552),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_4198),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_4200),
.Y(n_5255)
);

CKINVDCx20_ASAP7_75t_R g5256 ( 
.A(n_4555),
.Y(n_5256)
);

CKINVDCx5p33_ASAP7_75t_R g5257 ( 
.A(n_4560),
.Y(n_5257)
);

INVxp67_ASAP7_75t_L g5258 ( 
.A(n_4562),
.Y(n_5258)
);

CKINVDCx16_ASAP7_75t_R g5259 ( 
.A(n_4363),
.Y(n_5259)
);

CKINVDCx5p33_ASAP7_75t_R g5260 ( 
.A(n_4564),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_4201),
.Y(n_5261)
);

CKINVDCx5p33_ASAP7_75t_R g5262 ( 
.A(n_4565),
.Y(n_5262)
);

CKINVDCx16_ASAP7_75t_R g5263 ( 
.A(n_4422),
.Y(n_5263)
);

CKINVDCx5p33_ASAP7_75t_R g5264 ( 
.A(n_4566),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_4211),
.Y(n_5265)
);

INVxp33_ASAP7_75t_L g5266 ( 
.A(n_4069),
.Y(n_5266)
);

CKINVDCx20_ASAP7_75t_R g5267 ( 
.A(n_4572),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_4214),
.Y(n_5268)
);

CKINVDCx5p33_ASAP7_75t_R g5269 ( 
.A(n_4573),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_4216),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_4217),
.Y(n_5271)
);

BUFx3_ASAP7_75t_L g5272 ( 
.A(n_4542),
.Y(n_5272)
);

INVxp67_ASAP7_75t_SL g5273 ( 
.A(n_4533),
.Y(n_5273)
);

CKINVDCx5p33_ASAP7_75t_R g5274 ( 
.A(n_4576),
.Y(n_5274)
);

CKINVDCx20_ASAP7_75t_R g5275 ( 
.A(n_4583),
.Y(n_5275)
);

HB1xp67_ASAP7_75t_L g5276 ( 
.A(n_4586),
.Y(n_5276)
);

BUFx10_ASAP7_75t_L g5277 ( 
.A(n_4590),
.Y(n_5277)
);

INVx1_ASAP7_75t_L g5278 ( 
.A(n_4220),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_4223),
.Y(n_5279)
);

CKINVDCx5p33_ASAP7_75t_R g5280 ( 
.A(n_4597),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_4225),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_4229),
.Y(n_5282)
);

CKINVDCx5p33_ASAP7_75t_R g5283 ( 
.A(n_4602),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_4230),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_4231),
.Y(n_5285)
);

CKINVDCx5p33_ASAP7_75t_R g5286 ( 
.A(n_4604),
.Y(n_5286)
);

CKINVDCx20_ASAP7_75t_R g5287 ( 
.A(n_4608),
.Y(n_5287)
);

INVxp67_ASAP7_75t_SL g5288 ( 
.A(n_4632),
.Y(n_5288)
);

CKINVDCx14_ASAP7_75t_R g5289 ( 
.A(n_4314),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_4238),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_4240),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_4247),
.Y(n_5292)
);

CKINVDCx16_ASAP7_75t_R g5293 ( 
.A(n_4399),
.Y(n_5293)
);

CKINVDCx5p33_ASAP7_75t_R g5294 ( 
.A(n_4610),
.Y(n_5294)
);

BUFx2_ASAP7_75t_L g5295 ( 
.A(n_4611),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_4248),
.Y(n_5296)
);

INVxp33_ASAP7_75t_SL g5297 ( 
.A(n_4613),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_4249),
.Y(n_5298)
);

CKINVDCx20_ASAP7_75t_R g5299 ( 
.A(n_4614),
.Y(n_5299)
);

CKINVDCx20_ASAP7_75t_R g5300 ( 
.A(n_4619),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_4251),
.Y(n_5301)
);

CKINVDCx5p33_ASAP7_75t_R g5302 ( 
.A(n_4621),
.Y(n_5302)
);

INVx1_ASAP7_75t_L g5303 ( 
.A(n_4259),
.Y(n_5303)
);

INVxp67_ASAP7_75t_SL g5304 ( 
.A(n_4670),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4262),
.Y(n_5305)
);

INVx2_ASAP7_75t_L g5306 ( 
.A(n_4542),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_4264),
.Y(n_5307)
);

INVx1_ASAP7_75t_L g5308 ( 
.A(n_4265),
.Y(n_5308)
);

CKINVDCx5p33_ASAP7_75t_R g5309 ( 
.A(n_4624),
.Y(n_5309)
);

INVxp67_ASAP7_75t_L g5310 ( 
.A(n_4627),
.Y(n_5310)
);

CKINVDCx20_ASAP7_75t_R g5311 ( 
.A(n_4629),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_4269),
.Y(n_5312)
);

CKINVDCx5p33_ASAP7_75t_R g5313 ( 
.A(n_4638),
.Y(n_5313)
);

CKINVDCx14_ASAP7_75t_R g5314 ( 
.A(n_4473),
.Y(n_5314)
);

INVx1_ASAP7_75t_L g5315 ( 
.A(n_4271),
.Y(n_5315)
);

INVxp67_ASAP7_75t_L g5316 ( 
.A(n_4639),
.Y(n_5316)
);

INVx3_ASAP7_75t_L g5317 ( 
.A(n_4628),
.Y(n_5317)
);

INVxp67_ASAP7_75t_L g5318 ( 
.A(n_4640),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_4272),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_4273),
.Y(n_5320)
);

INVx1_ASAP7_75t_L g5321 ( 
.A(n_4275),
.Y(n_5321)
);

CKINVDCx5p33_ASAP7_75t_R g5322 ( 
.A(n_4647),
.Y(n_5322)
);

CKINVDCx5p33_ASAP7_75t_R g5323 ( 
.A(n_4649),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_4276),
.Y(n_5324)
);

INVxp67_ASAP7_75t_SL g5325 ( 
.A(n_4679),
.Y(n_5325)
);

CKINVDCx5p33_ASAP7_75t_R g5326 ( 
.A(n_4653),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_4279),
.Y(n_5327)
);

CKINVDCx5p33_ASAP7_75t_R g5328 ( 
.A(n_4654),
.Y(n_5328)
);

BUFx10_ASAP7_75t_L g5329 ( 
.A(n_4714),
.Y(n_5329)
);

BUFx3_ASAP7_75t_L g5330 ( 
.A(n_4628),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_4281),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_4284),
.Y(n_5332)
);

CKINVDCx20_ASAP7_75t_R g5333 ( 
.A(n_4656),
.Y(n_5333)
);

INVxp67_ASAP7_75t_L g5334 ( 
.A(n_4657),
.Y(n_5334)
);

INVxp67_ASAP7_75t_L g5335 ( 
.A(n_4659),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_4291),
.Y(n_5336)
);

CKINVDCx5p33_ASAP7_75t_R g5337 ( 
.A(n_4662),
.Y(n_5337)
);

CKINVDCx14_ASAP7_75t_R g5338 ( 
.A(n_4663),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_4292),
.Y(n_5339)
);

CKINVDCx20_ASAP7_75t_R g5340 ( 
.A(n_4665),
.Y(n_5340)
);

INVxp33_ASAP7_75t_L g5341 ( 
.A(n_4648),
.Y(n_5341)
);

CKINVDCx5p33_ASAP7_75t_R g5342 ( 
.A(n_4666),
.Y(n_5342)
);

CKINVDCx20_ASAP7_75t_R g5343 ( 
.A(n_4667),
.Y(n_5343)
);

INVxp33_ASAP7_75t_SL g5344 ( 
.A(n_4668),
.Y(n_5344)
);

CKINVDCx5p33_ASAP7_75t_R g5345 ( 
.A(n_4669),
.Y(n_5345)
);

HB1xp67_ASAP7_75t_L g5346 ( 
.A(n_4678),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4295),
.Y(n_5347)
);

INVxp33_ASAP7_75t_SL g5348 ( 
.A(n_4692),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_4297),
.Y(n_5349)
);

INVxp33_ASAP7_75t_L g5350 ( 
.A(n_4456),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_4300),
.Y(n_5351)
);

INVxp67_ASAP7_75t_L g5352 ( 
.A(n_4696),
.Y(n_5352)
);

CKINVDCx20_ASAP7_75t_R g5353 ( 
.A(n_4697),
.Y(n_5353)
);

CKINVDCx20_ASAP7_75t_R g5354 ( 
.A(n_4705),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_4302),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_4306),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_4308),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_4310),
.Y(n_5358)
);

CKINVDCx20_ASAP7_75t_R g5359 ( 
.A(n_4711),
.Y(n_5359)
);

HB1xp67_ASAP7_75t_L g5360 ( 
.A(n_4713),
.Y(n_5360)
);

CKINVDCx5p33_ASAP7_75t_R g5361 ( 
.A(n_4267),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_4312),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_4316),
.Y(n_5363)
);

INVxp67_ASAP7_75t_L g5364 ( 
.A(n_4366),
.Y(n_5364)
);

HB1xp67_ASAP7_75t_L g5365 ( 
.A(n_4055),
.Y(n_5365)
);

CKINVDCx5p33_ASAP7_75t_R g5366 ( 
.A(n_4139),
.Y(n_5366)
);

CKINVDCx5p33_ASAP7_75t_R g5367 ( 
.A(n_4071),
.Y(n_5367)
);

INVx2_ASAP7_75t_L g5368 ( 
.A(n_4628),
.Y(n_5368)
);

INVxp33_ASAP7_75t_SL g5369 ( 
.A(n_4100),
.Y(n_5369)
);

CKINVDCx16_ASAP7_75t_R g5370 ( 
.A(n_4341),
.Y(n_5370)
);

INVxp67_ASAP7_75t_SL g5371 ( 
.A(n_4515),
.Y(n_5371)
);

CKINVDCx20_ASAP7_75t_R g5372 ( 
.A(n_4169),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_4319),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_4320),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_4324),
.Y(n_5375)
);

INVx1_ASAP7_75t_L g5376 ( 
.A(n_4327),
.Y(n_5376)
);

INVxp67_ASAP7_75t_SL g5377 ( 
.A(n_4244),
.Y(n_5377)
);

INVx2_ASAP7_75t_L g5378 ( 
.A(n_4645),
.Y(n_5378)
);

BUFx3_ASAP7_75t_L g5379 ( 
.A(n_4645),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_4328),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_4330),
.Y(n_5381)
);

CKINVDCx5p33_ASAP7_75t_R g5382 ( 
.A(n_4383),
.Y(n_5382)
);

INVxp67_ASAP7_75t_SL g5383 ( 
.A(n_4378),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_4332),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_4334),
.Y(n_5385)
);

BUFx3_ASAP7_75t_L g5386 ( 
.A(n_4645),
.Y(n_5386)
);

INVxp67_ASAP7_75t_SL g5387 ( 
.A(n_4245),
.Y(n_5387)
);

INVx1_ASAP7_75t_L g5388 ( 
.A(n_4336),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_4338),
.Y(n_5389)
);

CKINVDCx16_ASAP7_75t_R g5390 ( 
.A(n_4391),
.Y(n_5390)
);

BUFx3_ASAP7_75t_L g5391 ( 
.A(n_4703),
.Y(n_5391)
);

CKINVDCx5p33_ASAP7_75t_R g5392 ( 
.A(n_4414),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_4340),
.Y(n_5393)
);

BUFx3_ASAP7_75t_L g5394 ( 
.A(n_4703),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_4348),
.Y(n_5395)
);

CKINVDCx5p33_ASAP7_75t_R g5396 ( 
.A(n_4460),
.Y(n_5396)
);

INVx1_ASAP7_75t_L g5397 ( 
.A(n_4351),
.Y(n_5397)
);

CKINVDCx20_ASAP7_75t_R g5398 ( 
.A(n_4509),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_4703),
.Y(n_5399)
);

INVx1_ASAP7_75t_L g5400 ( 
.A(n_4622),
.Y(n_5400)
);

CKINVDCx5p33_ASAP7_75t_R g5401 ( 
.A(n_4528),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_4501),
.Y(n_5402)
);

CKINVDCx20_ASAP7_75t_R g5403 ( 
.A(n_4612),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_4599),
.Y(n_5404)
);

CKINVDCx20_ASAP7_75t_R g5405 ( 
.A(n_4061),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_4424),
.Y(n_5406)
);

INVx3_ASAP7_75t_L g5407 ( 
.A(n_4425),
.Y(n_5407)
);

INVx3_ASAP7_75t_L g5408 ( 
.A(n_4433),
.Y(n_5408)
);

BUFx6f_ASAP7_75t_L g5409 ( 
.A(n_4436),
.Y(n_5409)
);

INVxp67_ASAP7_75t_SL g5410 ( 
.A(n_4157),
.Y(n_5410)
);

INVx2_ASAP7_75t_L g5411 ( 
.A(n_4437),
.Y(n_5411)
);

BUFx3_ASAP7_75t_L g5412 ( 
.A(n_4439),
.Y(n_5412)
);

CKINVDCx20_ASAP7_75t_R g5413 ( 
.A(n_4317),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_4441),
.Y(n_5414)
);

BUFx2_ASAP7_75t_L g5415 ( 
.A(n_4450),
.Y(n_5415)
);

CKINVDCx5p33_ASAP7_75t_R g5416 ( 
.A(n_4475),
.Y(n_5416)
);

CKINVDCx5p33_ASAP7_75t_R g5417 ( 
.A(n_4459),
.Y(n_5417)
);

CKINVDCx20_ASAP7_75t_R g5418 ( 
.A(n_4463),
.Y(n_5418)
);

HB1xp67_ASAP7_75t_L g5419 ( 
.A(n_4465),
.Y(n_5419)
);

INVx1_ASAP7_75t_L g5420 ( 
.A(n_4442),
.Y(n_5420)
);

CKINVDCx5p33_ASAP7_75t_R g5421 ( 
.A(n_4469),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_4448),
.Y(n_5422)
);

CKINVDCx5p33_ASAP7_75t_R g5423 ( 
.A(n_4470),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_4449),
.Y(n_5424)
);

CKINVDCx16_ASAP7_75t_R g5425 ( 
.A(n_4471),
.Y(n_5425)
);

HB1xp67_ASAP7_75t_L g5426 ( 
.A(n_4718),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_5317),
.Y(n_5427)
);

OAI21x1_ASAP7_75t_L g5428 ( 
.A1(n_5105),
.A2(n_2756),
.B(n_2729),
.Y(n_5428)
);

AND2x4_ASAP7_75t_L g5429 ( 
.A(n_4794),
.B(n_4451),
.Y(n_5429)
);

NAND2xp5_ASAP7_75t_SL g5430 ( 
.A(n_4797),
.B(n_4126),
.Y(n_5430)
);

OA21x2_ASAP7_75t_L g5431 ( 
.A1(n_5113),
.A2(n_3038),
.B(n_3032),
.Y(n_5431)
);

NAND2xp5_ASAP7_75t_L g5432 ( 
.A(n_5093),
.B(n_2921),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_4993),
.Y(n_5433)
);

OAI22x1_ASAP7_75t_L g5434 ( 
.A1(n_4817),
.A2(n_4452),
.B1(n_3016),
.B2(n_3048),
.Y(n_5434)
);

INVx5_ASAP7_75t_L g5435 ( 
.A(n_4788),
.Y(n_5435)
);

AND2x2_ASAP7_75t_L g5436 ( 
.A(n_4970),
.B(n_3283),
.Y(n_5436)
);

INVx2_ASAP7_75t_SL g5437 ( 
.A(n_4776),
.Y(n_5437)
);

BUFx6f_ASAP7_75t_L g5438 ( 
.A(n_4918),
.Y(n_5438)
);

BUFx8_ASAP7_75t_SL g5439 ( 
.A(n_4719),
.Y(n_5439)
);

INVxp67_ASAP7_75t_L g5440 ( 
.A(n_4822),
.Y(n_5440)
);

BUFx12f_ASAP7_75t_L g5441 ( 
.A(n_5277),
.Y(n_5441)
);

NOR2x1_ASAP7_75t_L g5442 ( 
.A(n_4942),
.B(n_3039),
.Y(n_5442)
);

INVx2_ASAP7_75t_L g5443 ( 
.A(n_5317),
.Y(n_5443)
);

CKINVDCx6p67_ASAP7_75t_R g5444 ( 
.A(n_4987),
.Y(n_5444)
);

AND2x2_ASAP7_75t_L g5445 ( 
.A(n_5038),
.B(n_3293),
.Y(n_5445)
);

AOI22xp5_ASAP7_75t_L g5446 ( 
.A1(n_5369),
.A2(n_2878),
.B1(n_2879),
.B2(n_2876),
.Y(n_5446)
);

AOI22xp5_ASAP7_75t_L g5447 ( 
.A1(n_5211),
.A2(n_5370),
.B1(n_5371),
.B2(n_5410),
.Y(n_5447)
);

AND2x2_ASAP7_75t_L g5448 ( 
.A(n_4722),
.B(n_4775),
.Y(n_5448)
);

AOI22xp5_ASAP7_75t_L g5449 ( 
.A1(n_5387),
.A2(n_2884),
.B1(n_2886),
.B2(n_2883),
.Y(n_5449)
);

BUFx2_ASAP7_75t_L g5450 ( 
.A(n_5405),
.Y(n_5450)
);

INVx2_ASAP7_75t_L g5451 ( 
.A(n_5272),
.Y(n_5451)
);

INVx2_ASAP7_75t_L g5452 ( 
.A(n_5330),
.Y(n_5452)
);

NOR2xp33_ASAP7_75t_L g5453 ( 
.A(n_5273),
.B(n_2953),
.Y(n_5453)
);

BUFx8_ASAP7_75t_SL g5454 ( 
.A(n_4728),
.Y(n_5454)
);

OA21x2_ASAP7_75t_L g5455 ( 
.A1(n_5114),
.A2(n_3043),
.B(n_3040),
.Y(n_5455)
);

INVx2_ASAP7_75t_L g5456 ( 
.A(n_5379),
.Y(n_5456)
);

NAND2xp5_ASAP7_75t_L g5457 ( 
.A(n_5377),
.B(n_2972),
.Y(n_5457)
);

AND2x4_ASAP7_75t_L g5458 ( 
.A(n_4789),
.B(n_2805),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_5001),
.Y(n_5459)
);

INVx4_ASAP7_75t_L g5460 ( 
.A(n_4745),
.Y(n_5460)
);

INVx2_ASAP7_75t_L g5461 ( 
.A(n_5386),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_4833),
.Y(n_5462)
);

CKINVDCx16_ASAP7_75t_R g5463 ( 
.A(n_4800),
.Y(n_5463)
);

NOR2xp33_ASAP7_75t_L g5464 ( 
.A(n_5288),
.B(n_5304),
.Y(n_5464)
);

BUFx12f_ASAP7_75t_L g5465 ( 
.A(n_5277),
.Y(n_5465)
);

BUFx3_ASAP7_75t_L g5466 ( 
.A(n_4992),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_4834),
.Y(n_5467)
);

INVx4_ASAP7_75t_L g5468 ( 
.A(n_4753),
.Y(n_5468)
);

OA21x2_ASAP7_75t_L g5469 ( 
.A1(n_5115),
.A2(n_3060),
.B(n_3053),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_4839),
.Y(n_5470)
);

BUFx6f_ASAP7_75t_L g5471 ( 
.A(n_5391),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_4840),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_4841),
.Y(n_5473)
);

BUFx6f_ASAP7_75t_L g5474 ( 
.A(n_5394),
.Y(n_5474)
);

INVx2_ASAP7_75t_SL g5475 ( 
.A(n_4858),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_SL g5476 ( 
.A(n_4975),
.B(n_2887),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_4842),
.Y(n_5477)
);

INVx2_ASAP7_75t_L g5478 ( 
.A(n_5252),
.Y(n_5478)
);

BUFx12f_ASAP7_75t_L g5479 ( 
.A(n_5329),
.Y(n_5479)
);

BUFx6f_ASAP7_75t_L g5480 ( 
.A(n_5157),
.Y(n_5480)
);

HB1xp67_ASAP7_75t_L g5481 ( 
.A(n_4799),
.Y(n_5481)
);

OA21x2_ASAP7_75t_L g5482 ( 
.A1(n_5117),
.A2(n_3063),
.B(n_3061),
.Y(n_5482)
);

BUFx6f_ASAP7_75t_L g5483 ( 
.A(n_5157),
.Y(n_5483)
);

AND2x4_ASAP7_75t_L g5484 ( 
.A(n_4819),
.B(n_2983),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_4843),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_5306),
.Y(n_5486)
);

INVx3_ASAP7_75t_L g5487 ( 
.A(n_5072),
.Y(n_5487)
);

AOI22xp5_ASAP7_75t_L g5488 ( 
.A1(n_5383),
.A2(n_2891),
.B1(n_2893),
.B2(n_2888),
.Y(n_5488)
);

BUFx8_ASAP7_75t_L g5489 ( 
.A(n_4835),
.Y(n_5489)
);

BUFx6f_ASAP7_75t_L g5490 ( 
.A(n_5157),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_4846),
.Y(n_5491)
);

BUFx6f_ASAP7_75t_L g5492 ( 
.A(n_5169),
.Y(n_5492)
);

NAND2xp33_ASAP7_75t_L g5493 ( 
.A(n_4820),
.B(n_2894),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_4847),
.Y(n_5494)
);

CKINVDCx11_ASAP7_75t_R g5495 ( 
.A(n_5015),
.Y(n_5495)
);

NOR2xp33_ASAP7_75t_L g5496 ( 
.A(n_5325),
.B(n_3010),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_5138),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5139),
.Y(n_5498)
);

INVx4_ASAP7_75t_L g5499 ( 
.A(n_4761),
.Y(n_5499)
);

NAND2xp5_ASAP7_75t_L g5500 ( 
.A(n_4725),
.B(n_3160),
.Y(n_5500)
);

AOI22xp5_ASAP7_75t_L g5501 ( 
.A1(n_5059),
.A2(n_4963),
.B1(n_4936),
.B2(n_5338),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_5140),
.Y(n_5502)
);

CKINVDCx8_ASAP7_75t_R g5503 ( 
.A(n_4823),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_4729),
.B(n_3229),
.Y(n_5504)
);

AND2x2_ASAP7_75t_L g5505 ( 
.A(n_4827),
.B(n_3293),
.Y(n_5505)
);

AND2x4_ASAP7_75t_L g5506 ( 
.A(n_4851),
.B(n_3058),
.Y(n_5506)
);

OAI22xp5_ASAP7_75t_L g5507 ( 
.A1(n_5400),
.A2(n_2896),
.B1(n_2906),
.B2(n_2902),
.Y(n_5507)
);

AND2x2_ASAP7_75t_L g5508 ( 
.A(n_4870),
.B(n_3311),
.Y(n_5508)
);

HB1xp67_ASAP7_75t_L g5509 ( 
.A(n_4930),
.Y(n_5509)
);

AOI22xp5_ASAP7_75t_L g5510 ( 
.A1(n_5027),
.A2(n_2909),
.B1(n_2910),
.B2(n_2907),
.Y(n_5510)
);

NAND2xp5_ASAP7_75t_L g5511 ( 
.A(n_4736),
.B(n_3304),
.Y(n_5511)
);

AND2x4_ASAP7_75t_L g5512 ( 
.A(n_4857),
.B(n_3066),
.Y(n_5512)
);

INVx3_ASAP7_75t_L g5513 ( 
.A(n_5163),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5145),
.Y(n_5514)
);

AND2x6_ASAP7_75t_L g5515 ( 
.A(n_5118),
.B(n_5402),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5151),
.Y(n_5516)
);

NAND2xp5_ASAP7_75t_L g5517 ( 
.A(n_4737),
.B(n_4738),
.Y(n_5517)
);

BUFx6f_ASAP7_75t_L g5518 ( 
.A(n_5169),
.Y(n_5518)
);

INVx1_ASAP7_75t_L g5519 ( 
.A(n_5154),
.Y(n_5519)
);

CKINVDCx20_ASAP7_75t_R g5520 ( 
.A(n_5017),
.Y(n_5520)
);

AND2x4_ASAP7_75t_L g5521 ( 
.A(n_4892),
.B(n_3171),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_5368),
.Y(n_5522)
);

BUFx6f_ASAP7_75t_L g5523 ( 
.A(n_5169),
.Y(n_5523)
);

INVx3_ASAP7_75t_L g5524 ( 
.A(n_5244),
.Y(n_5524)
);

INVx1_ASAP7_75t_L g5525 ( 
.A(n_5155),
.Y(n_5525)
);

BUFx6f_ASAP7_75t_L g5526 ( 
.A(n_5236),
.Y(n_5526)
);

AND2x6_ASAP7_75t_L g5527 ( 
.A(n_5404),
.B(n_3215),
.Y(n_5527)
);

AOI22xp5_ASAP7_75t_L g5528 ( 
.A1(n_4941),
.A2(n_5021),
.B1(n_5146),
.B2(n_5012),
.Y(n_5528)
);

NAND2xp5_ASAP7_75t_L g5529 ( 
.A(n_4739),
.B(n_3334),
.Y(n_5529)
);

AND2x4_ASAP7_75t_L g5530 ( 
.A(n_4911),
.B(n_3303),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_5159),
.Y(n_5531)
);

CKINVDCx5p33_ASAP7_75t_R g5532 ( 
.A(n_4945),
.Y(n_5532)
);

BUFx2_ASAP7_75t_L g5533 ( 
.A(n_5413),
.Y(n_5533)
);

INVx2_ASAP7_75t_L g5534 ( 
.A(n_5378),
.Y(n_5534)
);

CKINVDCx11_ASAP7_75t_R g5535 ( 
.A(n_5041),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_5161),
.Y(n_5536)
);

AND2x2_ASAP7_75t_L g5537 ( 
.A(n_5147),
.B(n_3311),
.Y(n_5537)
);

OAI22xp5_ASAP7_75t_SL g5538 ( 
.A1(n_5372),
.A2(n_3290),
.B1(n_3379),
.B2(n_3274),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_5172),
.Y(n_5539)
);

NAND2xp5_ASAP7_75t_L g5540 ( 
.A(n_4741),
.B(n_3380),
.Y(n_5540)
);

INVx2_ASAP7_75t_L g5541 ( 
.A(n_5399),
.Y(n_5541)
);

INVx2_ASAP7_75t_L g5542 ( 
.A(n_5183),
.Y(n_5542)
);

INVx1_ASAP7_75t_L g5543 ( 
.A(n_5173),
.Y(n_5543)
);

AND2x2_ASAP7_75t_L g5544 ( 
.A(n_5415),
.B(n_3321),
.Y(n_5544)
);

AOI22xp33_ASAP7_75t_SL g5545 ( 
.A1(n_5425),
.A2(n_3419),
.B1(n_3444),
.B2(n_3422),
.Y(n_5545)
);

OAI22xp5_ASAP7_75t_L g5546 ( 
.A1(n_5080),
.A2(n_2913),
.B1(n_2915),
.B2(n_2914),
.Y(n_5546)
);

NAND2xp5_ASAP7_75t_SL g5547 ( 
.A(n_5188),
.B(n_2917),
.Y(n_5547)
);

INVx3_ASAP7_75t_L g5548 ( 
.A(n_5409),
.Y(n_5548)
);

NAND2xp5_ASAP7_75t_L g5549 ( 
.A(n_4742),
.B(n_3402),
.Y(n_5549)
);

INVx3_ASAP7_75t_L g5550 ( 
.A(n_5409),
.Y(n_5550)
);

AND2x2_ASAP7_75t_L g5551 ( 
.A(n_5350),
.B(n_3321),
.Y(n_5551)
);

INVx2_ASAP7_75t_L g5552 ( 
.A(n_5185),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5174),
.Y(n_5553)
);

INVx2_ASAP7_75t_L g5554 ( 
.A(n_5186),
.Y(n_5554)
);

INVx1_ASAP7_75t_L g5555 ( 
.A(n_5175),
.Y(n_5555)
);

NOR2xp33_ASAP7_75t_L g5556 ( 
.A(n_4723),
.B(n_3417),
.Y(n_5556)
);

AND2x4_ASAP7_75t_L g5557 ( 
.A(n_4733),
.B(n_3428),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_5177),
.Y(n_5558)
);

AND2x4_ASAP7_75t_L g5559 ( 
.A(n_4768),
.B(n_4824),
.Y(n_5559)
);

INVx3_ASAP7_75t_L g5560 ( 
.A(n_5409),
.Y(n_5560)
);

AND2x4_ASAP7_75t_L g5561 ( 
.A(n_4837),
.B(n_3459),
.Y(n_5561)
);

AND2x4_ASAP7_75t_L g5562 ( 
.A(n_4912),
.B(n_3538),
.Y(n_5562)
);

INVx2_ASAP7_75t_L g5563 ( 
.A(n_5189),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_4744),
.Y(n_5564)
);

BUFx6f_ASAP7_75t_L g5565 ( 
.A(n_5236),
.Y(n_5565)
);

INVx3_ASAP7_75t_L g5566 ( 
.A(n_5412),
.Y(n_5566)
);

INVx2_ASAP7_75t_L g5567 ( 
.A(n_5190),
.Y(n_5567)
);

INVx2_ASAP7_75t_L g5568 ( 
.A(n_5191),
.Y(n_5568)
);

INVx2_ASAP7_75t_SL g5569 ( 
.A(n_5329),
.Y(n_5569)
);

AND2x2_ASAP7_75t_L g5570 ( 
.A(n_5365),
.B(n_3580),
.Y(n_5570)
);

INVx2_ASAP7_75t_L g5571 ( 
.A(n_5192),
.Y(n_5571)
);

OA21x2_ASAP7_75t_L g5572 ( 
.A1(n_5119),
.A2(n_3069),
.B(n_3068),
.Y(n_5572)
);

BUFx6f_ASAP7_75t_L g5573 ( 
.A(n_5236),
.Y(n_5573)
);

BUFx6f_ASAP7_75t_L g5574 ( 
.A(n_4749),
.Y(n_5574)
);

NAND2xp5_ASAP7_75t_L g5575 ( 
.A(n_4746),
.B(n_3558),
.Y(n_5575)
);

AND2x2_ASAP7_75t_L g5576 ( 
.A(n_4763),
.B(n_3580),
.Y(n_5576)
);

AND2x2_ASAP7_75t_SL g5577 ( 
.A(n_4743),
.B(n_2769),
.Y(n_5577)
);

BUFx2_ASAP7_75t_L g5578 ( 
.A(n_5181),
.Y(n_5578)
);

INVx5_ASAP7_75t_L g5579 ( 
.A(n_4855),
.Y(n_5579)
);

BUFx2_ASAP7_75t_L g5580 ( 
.A(n_5289),
.Y(n_5580)
);

HB1xp67_ASAP7_75t_L g5581 ( 
.A(n_4958),
.Y(n_5581)
);

INVx1_ASAP7_75t_L g5582 ( 
.A(n_4748),
.Y(n_5582)
);

INVx2_ASAP7_75t_L g5583 ( 
.A(n_5193),
.Y(n_5583)
);

INVx3_ASAP7_75t_L g5584 ( 
.A(n_5407),
.Y(n_5584)
);

INVx2_ASAP7_75t_L g5585 ( 
.A(n_5194),
.Y(n_5585)
);

AOI22xp5_ASAP7_75t_L g5586 ( 
.A1(n_5200),
.A2(n_2922),
.B1(n_2927),
.B2(n_2925),
.Y(n_5586)
);

NAND2xp5_ASAP7_75t_L g5587 ( 
.A(n_4750),
.B(n_4752),
.Y(n_5587)
);

INVx2_ASAP7_75t_L g5588 ( 
.A(n_5196),
.Y(n_5588)
);

INVx1_ASAP7_75t_L g5589 ( 
.A(n_4754),
.Y(n_5589)
);

CKINVDCx6p67_ASAP7_75t_R g5590 ( 
.A(n_5046),
.Y(n_5590)
);

INVx2_ASAP7_75t_L g5591 ( 
.A(n_5197),
.Y(n_5591)
);

NAND2xp5_ASAP7_75t_L g5592 ( 
.A(n_4755),
.B(n_3599),
.Y(n_5592)
);

BUFx6f_ASAP7_75t_L g5593 ( 
.A(n_4749),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_4758),
.Y(n_5594)
);

HB1xp67_ASAP7_75t_L g5595 ( 
.A(n_4966),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_5199),
.Y(n_5596)
);

AOI22xp5_ASAP7_75t_L g5597 ( 
.A1(n_5297),
.A2(n_2929),
.B1(n_2933),
.B2(n_2931),
.Y(n_5597)
);

INVx2_ASAP7_75t_L g5598 ( 
.A(n_5201),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5203),
.Y(n_5599)
);

NAND2xp5_ASAP7_75t_L g5600 ( 
.A(n_4765),
.B(n_3631),
.Y(n_5600)
);

HB1xp67_ASAP7_75t_L g5601 ( 
.A(n_5314),
.Y(n_5601)
);

INVx2_ASAP7_75t_L g5602 ( 
.A(n_5204),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_4766),
.Y(n_5603)
);

BUFx3_ASAP7_75t_L g5604 ( 
.A(n_5047),
.Y(n_5604)
);

HB1xp67_ASAP7_75t_L g5605 ( 
.A(n_4974),
.Y(n_5605)
);

OA22x2_ASAP7_75t_SL g5606 ( 
.A1(n_5344),
.A2(n_3168),
.B1(n_3759),
.B2(n_2961),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_4767),
.Y(n_5607)
);

INVx2_ASAP7_75t_L g5608 ( 
.A(n_5206),
.Y(n_5608)
);

INVx1_ASAP7_75t_L g5609 ( 
.A(n_4769),
.Y(n_5609)
);

NAND2xp5_ASAP7_75t_L g5610 ( 
.A(n_4771),
.B(n_3722),
.Y(n_5610)
);

INVx3_ASAP7_75t_L g5611 ( 
.A(n_5407),
.Y(n_5611)
);

BUFx6f_ASAP7_75t_L g5612 ( 
.A(n_4749),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_4772),
.Y(n_5613)
);

NAND2xp5_ASAP7_75t_L g5614 ( 
.A(n_4778),
.B(n_3966),
.Y(n_5614)
);

BUFx2_ASAP7_75t_L g5615 ( 
.A(n_5049),
.Y(n_5615)
);

CKINVDCx20_ASAP7_75t_R g5616 ( 
.A(n_5057),
.Y(n_5616)
);

BUFx6f_ASAP7_75t_L g5617 ( 
.A(n_4891),
.Y(n_5617)
);

AND2x2_ASAP7_75t_L g5618 ( 
.A(n_4784),
.B(n_4786),
.Y(n_5618)
);

AND2x2_ASAP7_75t_L g5619 ( 
.A(n_5182),
.B(n_3707),
.Y(n_5619)
);

HB1xp67_ASAP7_75t_L g5620 ( 
.A(n_5293),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_4780),
.Y(n_5621)
);

INVx2_ASAP7_75t_L g5622 ( 
.A(n_5207),
.Y(n_5622)
);

INVx1_ASAP7_75t_L g5623 ( 
.A(n_4781),
.Y(n_5623)
);

AND2x2_ASAP7_75t_L g5624 ( 
.A(n_4882),
.B(n_3707),
.Y(n_5624)
);

INVx2_ASAP7_75t_SL g5625 ( 
.A(n_4988),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_4782),
.Y(n_5626)
);

INVx2_ASAP7_75t_L g5627 ( 
.A(n_5208),
.Y(n_5627)
);

BUFx3_ASAP7_75t_L g5628 ( 
.A(n_5075),
.Y(n_5628)
);

BUFx6f_ASAP7_75t_L g5629 ( 
.A(n_4891),
.Y(n_5629)
);

BUFx6f_ASAP7_75t_L g5630 ( 
.A(n_4891),
.Y(n_5630)
);

INVx2_ASAP7_75t_L g5631 ( 
.A(n_5246),
.Y(n_5631)
);

AND2x2_ASAP7_75t_L g5632 ( 
.A(n_4886),
.B(n_3746),
.Y(n_5632)
);

NAND2xp5_ASAP7_75t_L g5633 ( 
.A(n_4787),
.B(n_4790),
.Y(n_5633)
);

INVx5_ASAP7_75t_L g5634 ( 
.A(n_4759),
.Y(n_5634)
);

INVx4_ASAP7_75t_L g5635 ( 
.A(n_4777),
.Y(n_5635)
);

BUFx6f_ASAP7_75t_L g5636 ( 
.A(n_4907),
.Y(n_5636)
);

CKINVDCx5p33_ASAP7_75t_R g5637 ( 
.A(n_4946),
.Y(n_5637)
);

OAI22xp5_ASAP7_75t_L g5638 ( 
.A1(n_5215),
.A2(n_2934),
.B1(n_2937),
.B2(n_2935),
.Y(n_5638)
);

INVx2_ASAP7_75t_L g5639 ( 
.A(n_5249),
.Y(n_5639)
);

BUFx6f_ASAP7_75t_L g5640 ( 
.A(n_4907),
.Y(n_5640)
);

BUFx3_ASAP7_75t_L g5641 ( 
.A(n_5077),
.Y(n_5641)
);

INVx2_ASAP7_75t_L g5642 ( 
.A(n_5254),
.Y(n_5642)
);

AOI22xp5_ASAP7_75t_L g5643 ( 
.A1(n_5348),
.A2(n_2943),
.B1(n_2950),
.B2(n_2944),
.Y(n_5643)
);

AND2x4_ASAP7_75t_L g5644 ( 
.A(n_4924),
.B(n_3549),
.Y(n_5644)
);

NAND2xp5_ASAP7_75t_L g5645 ( 
.A(n_4803),
.B(n_3968),
.Y(n_5645)
);

BUFx2_ASAP7_75t_L g5646 ( 
.A(n_5095),
.Y(n_5646)
);

INVx3_ASAP7_75t_L g5647 ( 
.A(n_5408),
.Y(n_5647)
);

NAND2xp5_ASAP7_75t_L g5648 ( 
.A(n_4807),
.B(n_3977),
.Y(n_5648)
);

INVx2_ASAP7_75t_L g5649 ( 
.A(n_5255),
.Y(n_5649)
);

BUFx6f_ASAP7_75t_L g5650 ( 
.A(n_4907),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_4808),
.Y(n_5651)
);

INVx1_ASAP7_75t_L g5652 ( 
.A(n_4810),
.Y(n_5652)
);

BUFx2_ASAP7_75t_L g5653 ( 
.A(n_5099),
.Y(n_5653)
);

INVx2_ASAP7_75t_L g5654 ( 
.A(n_5261),
.Y(n_5654)
);

BUFx6f_ASAP7_75t_L g5655 ( 
.A(n_5092),
.Y(n_5655)
);

OA21x2_ASAP7_75t_L g5656 ( 
.A1(n_5120),
.A2(n_3075),
.B(n_3071),
.Y(n_5656)
);

NAND2xp5_ASAP7_75t_L g5657 ( 
.A(n_4812),
.B(n_3081),
.Y(n_5657)
);

BUFx6f_ASAP7_75t_L g5658 ( 
.A(n_5092),
.Y(n_5658)
);

BUFx6f_ASAP7_75t_L g5659 ( 
.A(n_5092),
.Y(n_5659)
);

INVx2_ASAP7_75t_L g5660 ( 
.A(n_5265),
.Y(n_5660)
);

AND2x2_ASAP7_75t_L g5661 ( 
.A(n_4897),
.B(n_3746),
.Y(n_5661)
);

INVx6_ASAP7_75t_L g5662 ( 
.A(n_5141),
.Y(n_5662)
);

INVx3_ASAP7_75t_L g5663 ( 
.A(n_5408),
.Y(n_5663)
);

INVxp67_ASAP7_75t_L g5664 ( 
.A(n_5048),
.Y(n_5664)
);

NAND2xp5_ASAP7_75t_L g5665 ( 
.A(n_4813),
.B(n_4818),
.Y(n_5665)
);

INVx3_ASAP7_75t_L g5666 ( 
.A(n_5209),
.Y(n_5666)
);

BUFx6f_ASAP7_75t_L g5667 ( 
.A(n_5162),
.Y(n_5667)
);

INVx4_ASAP7_75t_L g5668 ( 
.A(n_4783),
.Y(n_5668)
);

BUFx6f_ASAP7_75t_L g5669 ( 
.A(n_5162),
.Y(n_5669)
);

AND2x4_ASAP7_75t_L g5670 ( 
.A(n_4928),
.B(n_3565),
.Y(n_5670)
);

AND2x2_ASAP7_75t_L g5671 ( 
.A(n_5058),
.B(n_5110),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_4825),
.Y(n_5672)
);

OAI22xp5_ASAP7_75t_L g5673 ( 
.A1(n_5247),
.A2(n_2957),
.B1(n_2959),
.B2(n_2958),
.Y(n_5673)
);

OAI21x1_ASAP7_75t_L g5674 ( 
.A1(n_5122),
.A2(n_2873),
.B(n_2841),
.Y(n_5674)
);

INVx2_ASAP7_75t_L g5675 ( 
.A(n_5268),
.Y(n_5675)
);

NOR2x1_ASAP7_75t_L g5676 ( 
.A(n_5035),
.B(n_3083),
.Y(n_5676)
);

AND2x4_ASAP7_75t_L g5677 ( 
.A(n_4933),
.B(n_4938),
.Y(n_5677)
);

INVx2_ASAP7_75t_L g5678 ( 
.A(n_5270),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_4826),
.Y(n_5679)
);

BUFx6f_ASAP7_75t_L g5680 ( 
.A(n_5025),
.Y(n_5680)
);

AND2x4_ASAP7_75t_L g5681 ( 
.A(n_4951),
.B(n_3596),
.Y(n_5681)
);

INVx1_ASAP7_75t_L g5682 ( 
.A(n_4828),
.Y(n_5682)
);

CKINVDCx16_ASAP7_75t_R g5683 ( 
.A(n_4859),
.Y(n_5683)
);

HB1xp67_ASAP7_75t_L g5684 ( 
.A(n_5367),
.Y(n_5684)
);

INVxp67_ASAP7_75t_SL g5685 ( 
.A(n_4732),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_4830),
.Y(n_5686)
);

AND2x4_ASAP7_75t_L g5687 ( 
.A(n_5214),
.B(n_3617),
.Y(n_5687)
);

BUFx12f_ASAP7_75t_L g5688 ( 
.A(n_4720),
.Y(n_5688)
);

AOI22xp5_ASAP7_75t_L g5689 ( 
.A1(n_5416),
.A2(n_2967),
.B1(n_2973),
.B2(n_2971),
.Y(n_5689)
);

INVx2_ASAP7_75t_L g5690 ( 
.A(n_5271),
.Y(n_5690)
);

OA21x2_ASAP7_75t_L g5691 ( 
.A1(n_5123),
.A2(n_3093),
.B(n_3085),
.Y(n_5691)
);

BUFx6f_ASAP7_75t_L g5692 ( 
.A(n_5025),
.Y(n_5692)
);

INVx2_ASAP7_75t_L g5693 ( 
.A(n_5278),
.Y(n_5693)
);

INVx3_ASAP7_75t_L g5694 ( 
.A(n_5220),
.Y(n_5694)
);

OAI22xp5_ASAP7_75t_L g5695 ( 
.A1(n_5250),
.A2(n_2974),
.B1(n_2976),
.B2(n_2975),
.Y(n_5695)
);

INVx2_ASAP7_75t_L g5696 ( 
.A(n_5279),
.Y(n_5696)
);

OAI22xp5_ASAP7_75t_L g5697 ( 
.A1(n_5258),
.A2(n_2982),
.B1(n_2989),
.B2(n_2987),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_4871),
.Y(n_5698)
);

NAND2xp5_ASAP7_75t_SL g5699 ( 
.A(n_4950),
.B(n_2990),
.Y(n_5699)
);

INVx2_ASAP7_75t_L g5700 ( 
.A(n_5281),
.Y(n_5700)
);

INVx2_ASAP7_75t_SL g5701 ( 
.A(n_4994),
.Y(n_5701)
);

AND2x2_ASAP7_75t_L g5702 ( 
.A(n_5295),
.B(n_3844),
.Y(n_5702)
);

INVx3_ASAP7_75t_L g5703 ( 
.A(n_5221),
.Y(n_5703)
);

INVx2_ASAP7_75t_L g5704 ( 
.A(n_5282),
.Y(n_5704)
);

BUFx6f_ASAP7_75t_L g5705 ( 
.A(n_5039),
.Y(n_5705)
);

INVx2_ASAP7_75t_L g5706 ( 
.A(n_5284),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_4872),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_4873),
.Y(n_5708)
);

INVx2_ASAP7_75t_L g5709 ( 
.A(n_5285),
.Y(n_5709)
);

NAND2xp5_ASAP7_75t_L g5710 ( 
.A(n_5124),
.B(n_3097),
.Y(n_5710)
);

NOR2xp33_ASAP7_75t_L g5711 ( 
.A(n_5364),
.B(n_2792),
.Y(n_5711)
);

INVx2_ASAP7_75t_L g5712 ( 
.A(n_5290),
.Y(n_5712)
);

INVx2_ASAP7_75t_L g5713 ( 
.A(n_5291),
.Y(n_5713)
);

INVx2_ASAP7_75t_SL g5714 ( 
.A(n_5390),
.Y(n_5714)
);

AND2x4_ASAP7_75t_L g5715 ( 
.A(n_5310),
.B(n_3636),
.Y(n_5715)
);

INVx3_ASAP7_75t_L g5716 ( 
.A(n_5222),
.Y(n_5716)
);

INVx1_ASAP7_75t_L g5717 ( 
.A(n_4874),
.Y(n_5717)
);

INVx3_ASAP7_75t_L g5718 ( 
.A(n_5223),
.Y(n_5718)
);

NOR2x1_ASAP7_75t_L g5719 ( 
.A(n_5097),
.B(n_3099),
.Y(n_5719)
);

BUFx3_ASAP7_75t_L g5720 ( 
.A(n_5112),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_4876),
.Y(n_5721)
);

INVx1_ASAP7_75t_L g5722 ( 
.A(n_4877),
.Y(n_5722)
);

NAND2xp5_ASAP7_75t_L g5723 ( 
.A(n_5129),
.B(n_3100),
.Y(n_5723)
);

AND2x2_ASAP7_75t_L g5724 ( 
.A(n_4798),
.B(n_3844),
.Y(n_5724)
);

BUFx12f_ASAP7_75t_L g5725 ( 
.A(n_4724),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_4883),
.Y(n_5726)
);

AND2x4_ASAP7_75t_L g5727 ( 
.A(n_5316),
.B(n_3651),
.Y(n_5727)
);

BUFx6f_ASAP7_75t_L g5728 ( 
.A(n_5039),
.Y(n_5728)
);

INVx2_ASAP7_75t_L g5729 ( 
.A(n_5292),
.Y(n_5729)
);

INVx2_ASAP7_75t_L g5730 ( 
.A(n_5296),
.Y(n_5730)
);

BUFx8_ASAP7_75t_L g5731 ( 
.A(n_4835),
.Y(n_5731)
);

AND2x4_ASAP7_75t_L g5732 ( 
.A(n_5318),
.B(n_5334),
.Y(n_5732)
);

HB1xp67_ASAP7_75t_L g5733 ( 
.A(n_5259),
.Y(n_5733)
);

INVx2_ASAP7_75t_L g5734 ( 
.A(n_5298),
.Y(n_5734)
);

INVx2_ASAP7_75t_L g5735 ( 
.A(n_5301),
.Y(n_5735)
);

AND2x2_ASAP7_75t_L g5736 ( 
.A(n_4923),
.B(n_3884),
.Y(n_5736)
);

CKINVDCx5p33_ASAP7_75t_R g5737 ( 
.A(n_4957),
.Y(n_5737)
);

INVx2_ASAP7_75t_L g5738 ( 
.A(n_5303),
.Y(n_5738)
);

INVx2_ASAP7_75t_L g5739 ( 
.A(n_5305),
.Y(n_5739)
);

INVx3_ASAP7_75t_L g5740 ( 
.A(n_5225),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_4884),
.Y(n_5741)
);

NAND2xp33_ASAP7_75t_L g5742 ( 
.A(n_4785),
.B(n_2992),
.Y(n_5742)
);

BUFx3_ASAP7_75t_L g5743 ( 
.A(n_5142),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_4885),
.Y(n_5744)
);

OAI22xp5_ASAP7_75t_SL g5745 ( 
.A1(n_4730),
.A2(n_3456),
.B1(n_3464),
.B2(n_3454),
.Y(n_5745)
);

OAI22xp5_ASAP7_75t_SL g5746 ( 
.A1(n_4731),
.A2(n_3526),
.B1(n_3555),
.B2(n_3500),
.Y(n_5746)
);

INVx2_ASAP7_75t_L g5747 ( 
.A(n_5307),
.Y(n_5747)
);

BUFx6f_ASAP7_75t_L g5748 ( 
.A(n_5166),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_4887),
.Y(n_5749)
);

AND2x2_ASAP7_75t_L g5750 ( 
.A(n_4944),
.B(n_3884),
.Y(n_5750)
);

INVx2_ASAP7_75t_L g5751 ( 
.A(n_5308),
.Y(n_5751)
);

BUFx6f_ASAP7_75t_L g5752 ( 
.A(n_5198),
.Y(n_5752)
);

NAND2xp5_ASAP7_75t_L g5753 ( 
.A(n_5132),
.B(n_3105),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_4889),
.Y(n_5754)
);

OR2x2_ASAP7_75t_L g5755 ( 
.A(n_5263),
.B(n_3677),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_4894),
.Y(n_5756)
);

NOR2xp33_ASAP7_75t_L g5757 ( 
.A(n_5102),
.B(n_5103),
.Y(n_5757)
);

INVx2_ASAP7_75t_SL g5758 ( 
.A(n_5382),
.Y(n_5758)
);

HB1xp67_ASAP7_75t_L g5759 ( 
.A(n_5417),
.Y(n_5759)
);

NAND2xp5_ASAP7_75t_L g5760 ( 
.A(n_5133),
.B(n_3109),
.Y(n_5760)
);

OAI22xp5_ASAP7_75t_SL g5761 ( 
.A1(n_4735),
.A2(n_3608),
.B1(n_3613),
.B2(n_3597),
.Y(n_5761)
);

OAI22x1_ASAP7_75t_SL g5762 ( 
.A1(n_5150),
.A2(n_3690),
.B1(n_3741),
.B2(n_3626),
.Y(n_5762)
);

BUFx6f_ASAP7_75t_L g5763 ( 
.A(n_5213),
.Y(n_5763)
);

CKINVDCx5p33_ASAP7_75t_R g5764 ( 
.A(n_4964),
.Y(n_5764)
);

INVx3_ASAP7_75t_L g5765 ( 
.A(n_5226),
.Y(n_5765)
);

INVx2_ASAP7_75t_L g5766 ( 
.A(n_5312),
.Y(n_5766)
);

OAI22xp5_ASAP7_75t_SL g5767 ( 
.A1(n_4740),
.A2(n_3775),
.B1(n_3824),
.B2(n_3774),
.Y(n_5767)
);

INVx3_ASAP7_75t_L g5768 ( 
.A(n_5411),
.Y(n_5768)
);

BUFx6f_ASAP7_75t_L g5769 ( 
.A(n_5242),
.Y(n_5769)
);

INVx2_ASAP7_75t_L g5770 ( 
.A(n_5315),
.Y(n_5770)
);

INVx5_ASAP7_75t_L g5771 ( 
.A(n_4779),
.Y(n_5771)
);

AND2x4_ASAP7_75t_L g5772 ( 
.A(n_5335),
.B(n_3734),
.Y(n_5772)
);

INVx2_ASAP7_75t_L g5773 ( 
.A(n_5319),
.Y(n_5773)
);

BUFx6f_ASAP7_75t_L g5774 ( 
.A(n_5248),
.Y(n_5774)
);

OAI22xp5_ASAP7_75t_L g5775 ( 
.A1(n_5352),
.A2(n_2994),
.B1(n_2995),
.B2(n_2993),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_4895),
.Y(n_5776)
);

AND2x4_ASAP7_75t_L g5777 ( 
.A(n_5406),
.B(n_3815),
.Y(n_5777)
);

BUFx8_ASAP7_75t_L g5778 ( 
.A(n_4838),
.Y(n_5778)
);

AND2x2_ASAP7_75t_SL g5779 ( 
.A(n_4878),
.B(n_2881),
.Y(n_5779)
);

BUFx6f_ASAP7_75t_L g5780 ( 
.A(n_4734),
.Y(n_5780)
);

BUFx6f_ASAP7_75t_L g5781 ( 
.A(n_4757),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_4898),
.Y(n_5782)
);

HB1xp67_ASAP7_75t_L g5783 ( 
.A(n_5421),
.Y(n_5783)
);

BUFx6f_ASAP7_75t_L g5784 ( 
.A(n_4796),
.Y(n_5784)
);

INVx2_ASAP7_75t_L g5785 ( 
.A(n_5320),
.Y(n_5785)
);

CKINVDCx5p33_ASAP7_75t_R g5786 ( 
.A(n_4965),
.Y(n_5786)
);

NOR2x1_ASAP7_75t_L g5787 ( 
.A(n_4901),
.B(n_3110),
.Y(n_5787)
);

BUFx6f_ASAP7_75t_L g5788 ( 
.A(n_4801),
.Y(n_5788)
);

INVx1_ASAP7_75t_L g5789 ( 
.A(n_4904),
.Y(n_5789)
);

OAI21x1_ASAP7_75t_L g5790 ( 
.A1(n_5134),
.A2(n_2912),
.B(n_2908),
.Y(n_5790)
);

INVx5_ASAP7_75t_L g5791 ( 
.A(n_4902),
.Y(n_5791)
);

AND2x2_ASAP7_75t_L g5792 ( 
.A(n_5423),
.B(n_4973),
.Y(n_5792)
);

INVx3_ASAP7_75t_L g5793 ( 
.A(n_4905),
.Y(n_5793)
);

BUFx6f_ASAP7_75t_L g5794 ( 
.A(n_4802),
.Y(n_5794)
);

AND2x2_ASAP7_75t_L g5795 ( 
.A(n_4978),
.B(n_3945),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_4906),
.Y(n_5796)
);

BUFx6f_ASAP7_75t_L g5797 ( 
.A(n_4804),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_4915),
.Y(n_5798)
);

INVx6_ASAP7_75t_L g5799 ( 
.A(n_4996),
.Y(n_5799)
);

NOR2x1_ASAP7_75t_L g5800 ( 
.A(n_4916),
.B(n_3115),
.Y(n_5800)
);

INVx1_ASAP7_75t_L g5801 ( 
.A(n_4920),
.Y(n_5801)
);

BUFx6f_ASAP7_75t_L g5802 ( 
.A(n_4831),
.Y(n_5802)
);

OAI22x1_ASAP7_75t_R g5803 ( 
.A1(n_5156),
.A2(n_3870),
.B1(n_3903),
.B2(n_3858),
.Y(n_5803)
);

INVx2_ASAP7_75t_L g5804 ( 
.A(n_5321),
.Y(n_5804)
);

NAND2xp5_ASAP7_75t_L g5805 ( 
.A(n_5135),
.B(n_3117),
.Y(n_5805)
);

BUFx3_ASAP7_75t_L g5806 ( 
.A(n_5167),
.Y(n_5806)
);

AND2x2_ASAP7_75t_L g5807 ( 
.A(n_4990),
.B(n_3945),
.Y(n_5807)
);

AND2x2_ASAP7_75t_L g5808 ( 
.A(n_4997),
.B(n_3980),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_4925),
.Y(n_5809)
);

BUFx6f_ASAP7_75t_L g5810 ( 
.A(n_4850),
.Y(n_5810)
);

NAND2xp5_ASAP7_75t_L g5811 ( 
.A(n_4849),
.B(n_3133),
.Y(n_5811)
);

AND2x2_ASAP7_75t_L g5812 ( 
.A(n_4999),
.B(n_3980),
.Y(n_5812)
);

AND2x2_ASAP7_75t_L g5813 ( 
.A(n_5009),
.B(n_4009),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_4927),
.Y(n_5814)
);

OAI22xp5_ASAP7_75t_SL g5815 ( 
.A1(n_4747),
.A2(n_3938),
.B1(n_3955),
.B2(n_3916),
.Y(n_5815)
);

INVx2_ASAP7_75t_L g5816 ( 
.A(n_5324),
.Y(n_5816)
);

INVx1_ASAP7_75t_L g5817 ( 
.A(n_4929),
.Y(n_5817)
);

BUFx6f_ASAP7_75t_L g5818 ( 
.A(n_4880),
.Y(n_5818)
);

NOR2xp33_ASAP7_75t_L g5819 ( 
.A(n_4716),
.B(n_3169),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_4931),
.Y(n_5820)
);

BUFx6f_ASAP7_75t_L g5821 ( 
.A(n_4909),
.Y(n_5821)
);

CKINVDCx20_ASAP7_75t_R g5822 ( 
.A(n_5176),
.Y(n_5822)
);

BUFx6f_ASAP7_75t_L g5823 ( 
.A(n_4949),
.Y(n_5823)
);

NAND2xp33_ASAP7_75t_L g5824 ( 
.A(n_4791),
.B(n_2996),
.Y(n_5824)
);

BUFx2_ASAP7_75t_L g5825 ( 
.A(n_5178),
.Y(n_5825)
);

INVxp67_ASAP7_75t_L g5826 ( 
.A(n_5010),
.Y(n_5826)
);

INVx4_ASAP7_75t_L g5827 ( 
.A(n_4795),
.Y(n_5827)
);

NAND2xp5_ASAP7_75t_L g5828 ( 
.A(n_4852),
.B(n_3136),
.Y(n_5828)
);

INVx3_ASAP7_75t_L g5829 ( 
.A(n_4935),
.Y(n_5829)
);

INVx2_ASAP7_75t_L g5830 ( 
.A(n_5327),
.Y(n_5830)
);

NAND2xp5_ASAP7_75t_L g5831 ( 
.A(n_4853),
.B(n_3138),
.Y(n_5831)
);

INVx2_ASAP7_75t_L g5832 ( 
.A(n_5331),
.Y(n_5832)
);

AND2x2_ASAP7_75t_L g5833 ( 
.A(n_5028),
.B(n_4009),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_4937),
.Y(n_5834)
);

INVx3_ASAP7_75t_L g5835 ( 
.A(n_4940),
.Y(n_5835)
);

INVx2_ASAP7_75t_L g5836 ( 
.A(n_5332),
.Y(n_5836)
);

INVx2_ASAP7_75t_L g5837 ( 
.A(n_5336),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_4943),
.Y(n_5838)
);

BUFx2_ASAP7_75t_L g5839 ( 
.A(n_5212),
.Y(n_5839)
);

INVx3_ASAP7_75t_L g5840 ( 
.A(n_4947),
.Y(n_5840)
);

INVx2_ASAP7_75t_L g5841 ( 
.A(n_5339),
.Y(n_5841)
);

INVx1_ASAP7_75t_L g5842 ( 
.A(n_4954),
.Y(n_5842)
);

INVx2_ASAP7_75t_L g5843 ( 
.A(n_5347),
.Y(n_5843)
);

INVx2_ASAP7_75t_L g5844 ( 
.A(n_5349),
.Y(n_5844)
);

AND2x4_ASAP7_75t_L g5845 ( 
.A(n_5414),
.B(n_3825),
.Y(n_5845)
);

AND2x2_ASAP7_75t_L g5846 ( 
.A(n_5031),
.B(n_3833),
.Y(n_5846)
);

AND2x6_ASAP7_75t_L g5847 ( 
.A(n_5420),
.B(n_3998),
.Y(n_5847)
);

INVx2_ASAP7_75t_L g5848 ( 
.A(n_5351),
.Y(n_5848)
);

CKINVDCx5p33_ASAP7_75t_R g5849 ( 
.A(n_5032),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_4955),
.Y(n_5850)
);

NAND2xp5_ASAP7_75t_L g5851 ( 
.A(n_4861),
.B(n_3139),
.Y(n_5851)
);

OAI21x1_ASAP7_75t_L g5852 ( 
.A1(n_4862),
.A2(n_2936),
.B(n_2920),
.Y(n_5852)
);

INVx3_ASAP7_75t_L g5853 ( 
.A(n_4956),
.Y(n_5853)
);

NAND2xp5_ASAP7_75t_L g5854 ( 
.A(n_4863),
.B(n_3143),
.Y(n_5854)
);

BUFx12f_ASAP7_75t_L g5855 ( 
.A(n_4726),
.Y(n_5855)
);

AND2x2_ASAP7_75t_L g5856 ( 
.A(n_5034),
.B(n_3135),
.Y(n_5856)
);

INVx2_ASAP7_75t_L g5857 ( 
.A(n_5355),
.Y(n_5857)
);

OAI21x1_ASAP7_75t_L g5858 ( 
.A1(n_4865),
.A2(n_2947),
.B(n_2939),
.Y(n_5858)
);

INVx2_ASAP7_75t_L g5859 ( 
.A(n_5356),
.Y(n_5859)
);

AOI22xp5_ASAP7_75t_L g5860 ( 
.A1(n_5043),
.A2(n_3003),
.B1(n_3006),
.B2(n_2997),
.Y(n_5860)
);

OAI21x1_ASAP7_75t_L g5861 ( 
.A1(n_4866),
.A2(n_4869),
.B(n_4868),
.Y(n_5861)
);

INVx2_ASAP7_75t_L g5862 ( 
.A(n_5357),
.Y(n_5862)
);

CKINVDCx20_ASAP7_75t_R g5863 ( 
.A(n_5237),
.Y(n_5863)
);

INVx2_ASAP7_75t_L g5864 ( 
.A(n_5358),
.Y(n_5864)
);

BUFx6f_ASAP7_75t_L g5865 ( 
.A(n_4971),
.Y(n_5865)
);

INVx1_ASAP7_75t_L g5866 ( 
.A(n_4959),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_4960),
.Y(n_5867)
);

AND2x2_ASAP7_75t_L g5868 ( 
.A(n_5056),
.B(n_3159),
.Y(n_5868)
);

INVx2_ASAP7_75t_L g5869 ( 
.A(n_5362),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_4961),
.Y(n_5870)
);

AND2x4_ASAP7_75t_L g5871 ( 
.A(n_5422),
.B(n_3145),
.Y(n_5871)
);

INVx2_ASAP7_75t_L g5872 ( 
.A(n_5363),
.Y(n_5872)
);

NOR2x1_ASAP7_75t_L g5873 ( 
.A(n_4962),
.B(n_3151),
.Y(n_5873)
);

INVx3_ASAP7_75t_L g5874 ( 
.A(n_4968),
.Y(n_5874)
);

CKINVDCx5p33_ASAP7_75t_R g5875 ( 
.A(n_5062),
.Y(n_5875)
);

INVxp67_ASAP7_75t_L g5876 ( 
.A(n_5036),
.Y(n_5876)
);

AOI22x1_ASAP7_75t_SL g5877 ( 
.A1(n_4751),
.A2(n_3981),
.B1(n_3996),
.B2(n_3975),
.Y(n_5877)
);

INVx3_ASAP7_75t_L g5878 ( 
.A(n_4969),
.Y(n_5878)
);

BUFx6f_ASAP7_75t_L g5879 ( 
.A(n_4998),
.Y(n_5879)
);

OAI21x1_ASAP7_75t_L g5880 ( 
.A1(n_4972),
.A2(n_2986),
.B(n_2984),
.Y(n_5880)
);

INVx2_ASAP7_75t_L g5881 ( 
.A(n_5373),
.Y(n_5881)
);

INVx2_ASAP7_75t_SL g5882 ( 
.A(n_5392),
.Y(n_5882)
);

NOR2xp33_ASAP7_75t_L g5883 ( 
.A(n_4717),
.B(n_3279),
.Y(n_5883)
);

INVx2_ASAP7_75t_L g5884 ( 
.A(n_5374),
.Y(n_5884)
);

AOI22x1_ASAP7_75t_SL g5885 ( 
.A1(n_4756),
.A2(n_4002),
.B1(n_4008),
.B2(n_3999),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_4976),
.Y(n_5886)
);

INVx2_ASAP7_75t_L g5887 ( 
.A(n_5375),
.Y(n_5887)
);

HB1xp67_ASAP7_75t_L g5888 ( 
.A(n_5008),
.Y(n_5888)
);

INVx2_ASAP7_75t_L g5889 ( 
.A(n_5376),
.Y(n_5889)
);

BUFx3_ASAP7_75t_L g5890 ( 
.A(n_5243),
.Y(n_5890)
);

BUFx2_ASAP7_75t_L g5891 ( 
.A(n_5256),
.Y(n_5891)
);

AND2x2_ASAP7_75t_SL g5892 ( 
.A(n_4952),
.B(n_3052),
.Y(n_5892)
);

INVx2_ASAP7_75t_L g5893 ( 
.A(n_5380),
.Y(n_5893)
);

INVx2_ASAP7_75t_L g5894 ( 
.A(n_5381),
.Y(n_5894)
);

INVxp33_ASAP7_75t_SL g5895 ( 
.A(n_4727),
.Y(n_5895)
);

INVx1_ASAP7_75t_L g5896 ( 
.A(n_4979),
.Y(n_5896)
);

XNOR2xp5_ASAP7_75t_L g5897 ( 
.A(n_4760),
.B(n_4019),
.Y(n_5897)
);

INVx3_ASAP7_75t_L g5898 ( 
.A(n_4980),
.Y(n_5898)
);

INVx3_ASAP7_75t_L g5899 ( 
.A(n_4981),
.Y(n_5899)
);

BUFx6f_ASAP7_75t_L g5900 ( 
.A(n_5000),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5384),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_4982),
.Y(n_5902)
);

INVx5_ASAP7_75t_L g5903 ( 
.A(n_4985),
.Y(n_5903)
);

OAI22xp5_ASAP7_75t_L g5904 ( 
.A1(n_5396),
.A2(n_3008),
.B1(n_3009),
.B2(n_3007),
.Y(n_5904)
);

INVx1_ASAP7_75t_L g5905 ( 
.A(n_4983),
.Y(n_5905)
);

BUFx6f_ASAP7_75t_L g5906 ( 
.A(n_5002),
.Y(n_5906)
);

INVx3_ASAP7_75t_L g5907 ( 
.A(n_4984),
.Y(n_5907)
);

AND2x2_ASAP7_75t_L g5908 ( 
.A(n_5078),
.B(n_3792),
.Y(n_5908)
);

AND2x2_ASAP7_75t_L g5909 ( 
.A(n_5087),
.B(n_3011),
.Y(n_5909)
);

NAND2xp5_ASAP7_75t_L g5910 ( 
.A(n_4721),
.B(n_3156),
.Y(n_5910)
);

INVx2_ASAP7_75t_L g5911 ( 
.A(n_5385),
.Y(n_5911)
);

BUFx6f_ASAP7_75t_L g5912 ( 
.A(n_5013),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_4986),
.Y(n_5913)
);

OAI21x1_ASAP7_75t_L g5914 ( 
.A1(n_4989),
.A2(n_3111),
.B(n_3082),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_4991),
.Y(n_5915)
);

INVx3_ASAP7_75t_L g5916 ( 
.A(n_4995),
.Y(n_5916)
);

INVxp67_ASAP7_75t_SL g5917 ( 
.A(n_5205),
.Y(n_5917)
);

INVx2_ASAP7_75t_SL g5918 ( 
.A(n_5401),
.Y(n_5918)
);

INVx4_ASAP7_75t_L g5919 ( 
.A(n_4805),
.Y(n_5919)
);

INVx1_ASAP7_75t_L g5920 ( 
.A(n_5003),
.Y(n_5920)
);

INVx2_ASAP7_75t_L g5921 ( 
.A(n_5388),
.Y(n_5921)
);

OAI22x1_ASAP7_75t_SL g5922 ( 
.A1(n_5267),
.A2(n_3018),
.B1(n_3019),
.B2(n_3015),
.Y(n_5922)
);

NAND2xp5_ASAP7_75t_L g5923 ( 
.A(n_5130),
.B(n_5131),
.Y(n_5923)
);

HB1xp67_ASAP7_75t_L g5924 ( 
.A(n_5106),
.Y(n_5924)
);

OA21x2_ASAP7_75t_L g5925 ( 
.A1(n_5004),
.A2(n_3167),
.B(n_3161),
.Y(n_5925)
);

CKINVDCx5p33_ASAP7_75t_R g5926 ( 
.A(n_5088),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_5006),
.Y(n_5927)
);

AND2x2_ASAP7_75t_SL g5928 ( 
.A(n_5040),
.B(n_5079),
.Y(n_5928)
);

INVx3_ASAP7_75t_L g5929 ( 
.A(n_5007),
.Y(n_5929)
);

INVx1_ASAP7_75t_L g5930 ( 
.A(n_5011),
.Y(n_5930)
);

INVx2_ASAP7_75t_SL g5931 ( 
.A(n_5090),
.Y(n_5931)
);

CKINVDCx5p33_ASAP7_75t_R g5932 ( 
.A(n_5094),
.Y(n_5932)
);

AND2x4_ASAP7_75t_L g5933 ( 
.A(n_5424),
.B(n_5419),
.Y(n_5933)
);

INVx3_ASAP7_75t_L g5934 ( 
.A(n_5014),
.Y(n_5934)
);

INVx6_ASAP7_75t_L g5935 ( 
.A(n_5111),
.Y(n_5935)
);

AND2x4_ASAP7_75t_L g5936 ( 
.A(n_5096),
.B(n_3179),
.Y(n_5936)
);

AND2x4_ASAP7_75t_L g5937 ( 
.A(n_5107),
.B(n_3181),
.Y(n_5937)
);

OAI22x1_ASAP7_75t_L g5938 ( 
.A1(n_5101),
.A2(n_3022),
.B1(n_3024),
.B2(n_3020),
.Y(n_5938)
);

INVx1_ASAP7_75t_L g5939 ( 
.A(n_5019),
.Y(n_5939)
);

BUFx2_ASAP7_75t_L g5940 ( 
.A(n_5275),
.Y(n_5940)
);

BUFx6f_ASAP7_75t_L g5941 ( 
.A(n_5018),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5020),
.Y(n_5942)
);

NOR2xp33_ASAP7_75t_L g5943 ( 
.A(n_4816),
.B(n_4829),
.Y(n_5943)
);

AOI22xp5_ASAP7_75t_L g5944 ( 
.A1(n_5104),
.A2(n_5125),
.B1(n_5126),
.B2(n_5116),
.Y(n_5944)
);

NAND2xp5_ASAP7_75t_L g5945 ( 
.A(n_5144),
.B(n_3185),
.Y(n_5945)
);

OAI22xp5_ASAP7_75t_SL g5946 ( 
.A1(n_4762),
.A2(n_3028),
.B1(n_3031),
.B2(n_3025),
.Y(n_5946)
);

INVx2_ASAP7_75t_L g5947 ( 
.A(n_5389),
.Y(n_5947)
);

NAND2xp5_ASAP7_75t_L g5948 ( 
.A(n_5152),
.B(n_3188),
.Y(n_5948)
);

INVx2_ASAP7_75t_L g5949 ( 
.A(n_5393),
.Y(n_5949)
);

INVx3_ASAP7_75t_L g5950 ( 
.A(n_5022),
.Y(n_5950)
);

INVx2_ASAP7_75t_L g5951 ( 
.A(n_5395),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5023),
.Y(n_5952)
);

NAND2xp5_ASAP7_75t_L g5953 ( 
.A(n_5158),
.B(n_3191),
.Y(n_5953)
);

BUFx3_ASAP7_75t_L g5954 ( 
.A(n_5287),
.Y(n_5954)
);

BUFx2_ASAP7_75t_L g5955 ( 
.A(n_5299),
.Y(n_5955)
);

NAND2xp33_ASAP7_75t_L g5956 ( 
.A(n_4806),
.B(n_3033),
.Y(n_5956)
);

OAI21x1_ASAP7_75t_L g5957 ( 
.A1(n_5024),
.A2(n_3124),
.B(n_3120),
.Y(n_5957)
);

INVx2_ASAP7_75t_SL g5958 ( 
.A(n_5127),
.Y(n_5958)
);

AOI22xp5_ASAP7_75t_L g5959 ( 
.A1(n_5128),
.A2(n_3037),
.B1(n_3042),
.B2(n_3035),
.Y(n_5959)
);

INVx5_ASAP7_75t_L g5960 ( 
.A(n_5042),
.Y(n_5960)
);

NAND2xp5_ASAP7_75t_L g5961 ( 
.A(n_5179),
.B(n_3193),
.Y(n_5961)
);

HB1xp67_ASAP7_75t_L g5962 ( 
.A(n_5136),
.Y(n_5962)
);

BUFx3_ASAP7_75t_L g5963 ( 
.A(n_5300),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5026),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5030),
.Y(n_5965)
);

INVx3_ASAP7_75t_L g5966 ( 
.A(n_5033),
.Y(n_5966)
);

AND2x4_ASAP7_75t_L g5967 ( 
.A(n_5109),
.B(n_3196),
.Y(n_5967)
);

OAI21x1_ASAP7_75t_L g5968 ( 
.A1(n_5037),
.A2(n_5045),
.B(n_5044),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5050),
.Y(n_5969)
);

BUFx6f_ASAP7_75t_L g5970 ( 
.A(n_5060),
.Y(n_5970)
);

INVx4_ASAP7_75t_L g5971 ( 
.A(n_4809),
.Y(n_5971)
);

NAND2xp5_ASAP7_75t_L g5972 ( 
.A(n_5051),
.B(n_5052),
.Y(n_5972)
);

INVx2_ASAP7_75t_L g5973 ( 
.A(n_5397),
.Y(n_5973)
);

INVx1_ASAP7_75t_L g5974 ( 
.A(n_5053),
.Y(n_5974)
);

BUFx8_ASAP7_75t_L g5975 ( 
.A(n_4838),
.Y(n_5975)
);

INVx2_ASAP7_75t_L g5976 ( 
.A(n_5061),
.Y(n_5976)
);

BUFx2_ASAP7_75t_L g5977 ( 
.A(n_5311),
.Y(n_5977)
);

BUFx2_ASAP7_75t_L g5978 ( 
.A(n_5333),
.Y(n_5978)
);

INVx5_ASAP7_75t_L g5979 ( 
.A(n_5266),
.Y(n_5979)
);

CKINVDCx11_ASAP7_75t_R g5980 ( 
.A(n_5340),
.Y(n_5980)
);

NAND2xp5_ASAP7_75t_L g5981 ( 
.A(n_5054),
.B(n_3198),
.Y(n_5981)
);

INVx2_ASAP7_75t_L g5982 ( 
.A(n_5227),
.Y(n_5982)
);

INVx3_ASAP7_75t_L g5983 ( 
.A(n_5055),
.Y(n_5983)
);

OAI21x1_ASAP7_75t_L g5984 ( 
.A1(n_5063),
.A2(n_3131),
.B(n_3126),
.Y(n_5984)
);

NAND2xp5_ASAP7_75t_L g5985 ( 
.A(n_5064),
.B(n_3203),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5065),
.Y(n_5986)
);

NAND2xp5_ASAP7_75t_L g5987 ( 
.A(n_5066),
.B(n_3204),
.Y(n_5987)
);

INVx2_ASAP7_75t_L g5988 ( 
.A(n_5228),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5231),
.Y(n_5989)
);

CKINVDCx6p67_ASAP7_75t_R g5990 ( 
.A(n_5343),
.Y(n_5990)
);

NOR2x1_ASAP7_75t_L g5991 ( 
.A(n_5067),
.B(n_3205),
.Y(n_5991)
);

OAI22xp5_ASAP7_75t_L g5992 ( 
.A1(n_5137),
.A2(n_3045),
.B1(n_3046),
.B2(n_3044),
.Y(n_5992)
);

AND2x4_ASAP7_75t_L g5993 ( 
.A(n_5121),
.B(n_3214),
.Y(n_5993)
);

BUFx6f_ASAP7_75t_L g5994 ( 
.A(n_5143),
.Y(n_5994)
);

OAI22x1_ASAP7_75t_SL g5995 ( 
.A1(n_5353),
.A2(n_3051),
.B1(n_3055),
.B2(n_3049),
.Y(n_5995)
);

NOR2xp33_ASAP7_75t_L g5996 ( 
.A(n_4921),
.B(n_3337),
.Y(n_5996)
);

AND2x4_ASAP7_75t_L g5997 ( 
.A(n_5148),
.B(n_5160),
.Y(n_5997)
);

HB1xp67_ASAP7_75t_L g5998 ( 
.A(n_5149),
.Y(n_5998)
);

INVx2_ASAP7_75t_L g5999 ( 
.A(n_5232),
.Y(n_5999)
);

BUFx2_ASAP7_75t_L g6000 ( 
.A(n_5354),
.Y(n_6000)
);

NAND2xp5_ASAP7_75t_L g6001 ( 
.A(n_5068),
.B(n_3216),
.Y(n_6001)
);

INVx2_ASAP7_75t_L g6002 ( 
.A(n_5235),
.Y(n_6002)
);

INVx5_ASAP7_75t_L g6003 ( 
.A(n_5005),
.Y(n_6003)
);

INVx3_ASAP7_75t_L g6004 ( 
.A(n_5069),
.Y(n_6004)
);

INVx2_ASAP7_75t_L g6005 ( 
.A(n_5238),
.Y(n_6005)
);

AND2x4_ASAP7_75t_L g6006 ( 
.A(n_5184),
.B(n_3218),
.Y(n_6006)
);

BUFx6f_ASAP7_75t_L g6007 ( 
.A(n_5153),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5070),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5071),
.Y(n_6009)
);

NAND2xp33_ASAP7_75t_L g6010 ( 
.A(n_4811),
.B(n_3057),
.Y(n_6010)
);

INVx2_ASAP7_75t_L g6011 ( 
.A(n_5239),
.Y(n_6011)
);

OA21x2_ASAP7_75t_L g6012 ( 
.A1(n_5073),
.A2(n_3233),
.B(n_3228),
.Y(n_6012)
);

INVx2_ASAP7_75t_L g6013 ( 
.A(n_5241),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5074),
.Y(n_6014)
);

CKINVDCx5p33_ASAP7_75t_R g6015 ( 
.A(n_5164),
.Y(n_6015)
);

CKINVDCx5p33_ASAP7_75t_R g6016 ( 
.A(n_5165),
.Y(n_6016)
);

OA21x2_ASAP7_75t_L g6017 ( 
.A1(n_5076),
.A2(n_5082),
.B(n_5081),
.Y(n_6017)
);

BUFx12f_ASAP7_75t_L g6018 ( 
.A(n_5168),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5083),
.Y(n_6019)
);

BUFx6f_ASAP7_75t_L g6020 ( 
.A(n_5170),
.Y(n_6020)
);

BUFx6f_ASAP7_75t_L g6021 ( 
.A(n_5171),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_5084),
.Y(n_6022)
);

AOI22xp5_ASAP7_75t_L g6023 ( 
.A1(n_5180),
.A2(n_3062),
.B1(n_3064),
.B2(n_3059),
.Y(n_6023)
);

NAND2xp5_ASAP7_75t_L g6024 ( 
.A(n_5085),
.B(n_3238),
.Y(n_6024)
);

HB1xp67_ASAP7_75t_L g6025 ( 
.A(n_5187),
.Y(n_6025)
);

BUFx6f_ASAP7_75t_L g6026 ( 
.A(n_5195),
.Y(n_6026)
);

NOR2xp33_ASAP7_75t_L g6027 ( 
.A(n_4922),
.B(n_3386),
.Y(n_6027)
);

HB1xp67_ASAP7_75t_L g6028 ( 
.A(n_5202),
.Y(n_6028)
);

HB1xp67_ASAP7_75t_L g6029 ( 
.A(n_5210),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_5086),
.Y(n_6030)
);

BUFx6f_ASAP7_75t_L g6031 ( 
.A(n_5218),
.Y(n_6031)
);

OAI22xp5_ASAP7_75t_L g6032 ( 
.A1(n_5219),
.A2(n_3067),
.B1(n_3070),
.B2(n_3065),
.Y(n_6032)
);

BUFx6f_ASAP7_75t_L g6033 ( 
.A(n_5224),
.Y(n_6033)
);

INVx3_ASAP7_75t_L g6034 ( 
.A(n_5091),
.Y(n_6034)
);

BUFx6f_ASAP7_75t_L g6035 ( 
.A(n_5229),
.Y(n_6035)
);

NAND2xp5_ASAP7_75t_L g6036 ( 
.A(n_5216),
.B(n_3241),
.Y(n_6036)
);

NOR2xp33_ASAP7_75t_L g6037 ( 
.A(n_4770),
.B(n_3436),
.Y(n_6037)
);

BUFx6f_ASAP7_75t_L g6038 ( 
.A(n_5230),
.Y(n_6038)
);

CKINVDCx11_ASAP7_75t_R g6039 ( 
.A(n_5359),
.Y(n_6039)
);

HB1xp67_ASAP7_75t_L g6040 ( 
.A(n_5234),
.Y(n_6040)
);

OA21x2_ASAP7_75t_L g6041 ( 
.A1(n_5089),
.A2(n_5100),
.B(n_5098),
.Y(n_6041)
);

NAND2xp5_ASAP7_75t_L g6042 ( 
.A(n_5217),
.B(n_3245),
.Y(n_6042)
);

INVx4_ASAP7_75t_L g6043 ( 
.A(n_4814),
.Y(n_6043)
);

BUFx6f_ASAP7_75t_L g6044 ( 
.A(n_5240),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5108),
.Y(n_6045)
);

NAND2xp5_ASAP7_75t_L g6046 ( 
.A(n_5245),
.B(n_3246),
.Y(n_6046)
);

BUFx6f_ASAP7_75t_L g6047 ( 
.A(n_5251),
.Y(n_6047)
);

AND2x2_ASAP7_75t_L g6048 ( 
.A(n_5257),
.B(n_3072),
.Y(n_6048)
);

BUFx6f_ASAP7_75t_L g6049 ( 
.A(n_5260),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_5233),
.Y(n_6050)
);

OAI22xp5_ASAP7_75t_L g6051 ( 
.A1(n_5262),
.A2(n_3076),
.B1(n_3078),
.B2(n_3074),
.Y(n_6051)
);

INVx2_ASAP7_75t_L g6052 ( 
.A(n_5253),
.Y(n_6052)
);

AND2x6_ASAP7_75t_L g6053 ( 
.A(n_4815),
.B(n_3247),
.Y(n_6053)
);

INVx3_ASAP7_75t_L g6054 ( 
.A(n_5264),
.Y(n_6054)
);

NAND2xp5_ASAP7_75t_L g6055 ( 
.A(n_5269),
.B(n_3249),
.Y(n_6055)
);

INVx2_ASAP7_75t_L g6056 ( 
.A(n_5276),
.Y(n_6056)
);

BUFx6f_ASAP7_75t_L g6057 ( 
.A(n_5274),
.Y(n_6057)
);

INVx2_ASAP7_75t_L g6058 ( 
.A(n_5346),
.Y(n_6058)
);

BUFx6f_ASAP7_75t_L g6059 ( 
.A(n_5280),
.Y(n_6059)
);

INVx2_ASAP7_75t_L g6060 ( 
.A(n_5360),
.Y(n_6060)
);

AND2x2_ASAP7_75t_L g6061 ( 
.A(n_5283),
.B(n_3079),
.Y(n_6061)
);

INVx2_ASAP7_75t_L g6062 ( 
.A(n_5029),
.Y(n_6062)
);

BUFx2_ASAP7_75t_L g6063 ( 
.A(n_5286),
.Y(n_6063)
);

INVx6_ASAP7_75t_L g6064 ( 
.A(n_4764),
.Y(n_6064)
);

AND2x4_ASAP7_75t_L g6065 ( 
.A(n_5398),
.B(n_3256),
.Y(n_6065)
);

INVx1_ASAP7_75t_L g6066 ( 
.A(n_5294),
.Y(n_6066)
);

INVx4_ASAP7_75t_L g6067 ( 
.A(n_4821),
.Y(n_6067)
);

AND2x6_ASAP7_75t_L g6068 ( 
.A(n_5029),
.B(n_3262),
.Y(n_6068)
);

INVx2_ASAP7_75t_L g6069 ( 
.A(n_5302),
.Y(n_6069)
);

BUFx3_ASAP7_75t_L g6070 ( 
.A(n_5309),
.Y(n_6070)
);

CKINVDCx11_ASAP7_75t_R g6071 ( 
.A(n_4773),
.Y(n_6071)
);

INVx3_ASAP7_75t_L g6072 ( 
.A(n_5313),
.Y(n_6072)
);

BUFx6f_ASAP7_75t_L g6073 ( 
.A(n_5322),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_5323),
.Y(n_6074)
);

BUFx6f_ASAP7_75t_L g6075 ( 
.A(n_5326),
.Y(n_6075)
);

INVx1_ASAP7_75t_L g6076 ( 
.A(n_5328),
.Y(n_6076)
);

INVx2_ASAP7_75t_L g6077 ( 
.A(n_5337),
.Y(n_6077)
);

AND2x2_ASAP7_75t_L g6078 ( 
.A(n_5342),
.B(n_3086),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5345),
.Y(n_6079)
);

AOI22xp5_ASAP7_75t_L g6080 ( 
.A1(n_4836),
.A2(n_3088),
.B1(n_3089),
.B2(n_3087),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_4845),
.Y(n_6081)
);

INVx1_ASAP7_75t_L g6082 ( 
.A(n_4848),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_4856),
.Y(n_6083)
);

CKINVDCx5p33_ASAP7_75t_R g6084 ( 
.A(n_4860),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_4864),
.Y(n_6085)
);

BUFx6f_ASAP7_75t_L g6086 ( 
.A(n_4867),
.Y(n_6086)
);

AND2x2_ASAP7_75t_SL g6087 ( 
.A(n_4879),
.B(n_3172),
.Y(n_6087)
);

INVx2_ASAP7_75t_L g6088 ( 
.A(n_4890),
.Y(n_6088)
);

INVx2_ASAP7_75t_L g6089 ( 
.A(n_4896),
.Y(n_6089)
);

NOR2xp33_ASAP7_75t_L g6090 ( 
.A(n_4900),
.B(n_3562),
.Y(n_6090)
);

NOR2x1_ASAP7_75t_L g6091 ( 
.A(n_5403),
.B(n_3272),
.Y(n_6091)
);

INVx6_ASAP7_75t_L g6092 ( 
.A(n_4774),
.Y(n_6092)
);

CKINVDCx5p33_ASAP7_75t_R g6093 ( 
.A(n_4903),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_4908),
.B(n_4910),
.Y(n_6094)
);

BUFx8_ASAP7_75t_L g6095 ( 
.A(n_4792),
.Y(n_6095)
);

AND2x2_ASAP7_75t_SL g6096 ( 
.A(n_4934),
.B(n_3173),
.Y(n_6096)
);

INVx2_ASAP7_75t_L g6097 ( 
.A(n_5418),
.Y(n_6097)
);

NAND2xp5_ASAP7_75t_L g6098 ( 
.A(n_5016),
.B(n_3282),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_5366),
.Y(n_6099)
);

NAND2xp5_ASAP7_75t_L g6100 ( 
.A(n_4948),
.B(n_3284),
.Y(n_6100)
);

INVx2_ASAP7_75t_L g6101 ( 
.A(n_4953),
.Y(n_6101)
);

INVx3_ASAP7_75t_L g6102 ( 
.A(n_5361),
.Y(n_6102)
);

AND2x2_ASAP7_75t_L g6103 ( 
.A(n_4967),
.B(n_3090),
.Y(n_6103)
);

OAI22xp5_ASAP7_75t_L g6104 ( 
.A1(n_4977),
.A2(n_3092),
.B1(n_3094),
.B2(n_3091),
.Y(n_6104)
);

INVx1_ASAP7_75t_L g6105 ( 
.A(n_4793),
.Y(n_6105)
);

INVx3_ASAP7_75t_L g6106 ( 
.A(n_4832),
.Y(n_6106)
);

INVx1_ASAP7_75t_L g6107 ( 
.A(n_4844),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_4854),
.Y(n_6108)
);

OAI21x1_ASAP7_75t_L g6109 ( 
.A1(n_4875),
.A2(n_3211),
.B(n_3180),
.Y(n_6109)
);

INVx1_ASAP7_75t_L g6110 ( 
.A(n_4881),
.Y(n_6110)
);

INVx2_ASAP7_75t_L g6111 ( 
.A(n_4888),
.Y(n_6111)
);

INVx3_ASAP7_75t_L g6112 ( 
.A(n_4893),
.Y(n_6112)
);

AND2x2_ASAP7_75t_L g6113 ( 
.A(n_5341),
.B(n_3095),
.Y(n_6113)
);

AOI22xp5_ASAP7_75t_L g6114 ( 
.A1(n_4899),
.A2(n_3102),
.B1(n_3103),
.B2(n_3098),
.Y(n_6114)
);

BUFx12f_ASAP7_75t_L g6115 ( 
.A(n_4913),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_4914),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_4917),
.Y(n_6117)
);

NAND2xp33_ASAP7_75t_L g6118 ( 
.A(n_4919),
.B(n_3104),
.Y(n_6118)
);

INVx2_ASAP7_75t_L g6119 ( 
.A(n_4926),
.Y(n_6119)
);

INVx3_ASAP7_75t_L g6120 ( 
.A(n_4932),
.Y(n_6120)
);

BUFx6f_ASAP7_75t_L g6121 ( 
.A(n_4939),
.Y(n_6121)
);

BUFx3_ASAP7_75t_L g6122 ( 
.A(n_4918),
.Y(n_6122)
);

BUFx6f_ASAP7_75t_L g6123 ( 
.A(n_4918),
.Y(n_6123)
);

BUFx8_ASAP7_75t_L g6124 ( 
.A(n_4835),
.Y(n_6124)
);

AND2x4_ASAP7_75t_L g6125 ( 
.A(n_4718),
.B(n_3285),
.Y(n_6125)
);

INVx3_ASAP7_75t_L g6126 ( 
.A(n_4918),
.Y(n_6126)
);

BUFx3_ASAP7_75t_L g6127 ( 
.A(n_4918),
.Y(n_6127)
);

INVx2_ASAP7_75t_L g6128 ( 
.A(n_5317),
.Y(n_6128)
);

INVx5_ASAP7_75t_L g6129 ( 
.A(n_4743),
.Y(n_6129)
);

INVx2_ASAP7_75t_L g6130 ( 
.A(n_5317),
.Y(n_6130)
);

AND2x4_ASAP7_75t_L g6131 ( 
.A(n_4718),
.B(n_3286),
.Y(n_6131)
);

INVx3_ASAP7_75t_L g6132 ( 
.A(n_4918),
.Y(n_6132)
);

INVx2_ASAP7_75t_L g6133 ( 
.A(n_5317),
.Y(n_6133)
);

INVx2_ASAP7_75t_L g6134 ( 
.A(n_5317),
.Y(n_6134)
);

INVx1_ASAP7_75t_L g6135 ( 
.A(n_4993),
.Y(n_6135)
);

BUFx12f_ASAP7_75t_L g6136 ( 
.A(n_5277),
.Y(n_6136)
);

OA21x2_ASAP7_75t_L g6137 ( 
.A1(n_5105),
.A2(n_3288),
.B(n_3287),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_4993),
.Y(n_6138)
);

OA21x2_ASAP7_75t_L g6139 ( 
.A1(n_5105),
.A2(n_3306),
.B(n_3299),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_4993),
.Y(n_6140)
);

CKINVDCx8_ASAP7_75t_R g6141 ( 
.A(n_4788),
.Y(n_6141)
);

CKINVDCx5p33_ASAP7_75t_R g6142 ( 
.A(n_4718),
.Y(n_6142)
);

BUFx6f_ASAP7_75t_L g6143 ( 
.A(n_4918),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_4993),
.Y(n_6144)
);

INVx1_ASAP7_75t_L g6145 ( 
.A(n_4993),
.Y(n_6145)
);

INVx5_ASAP7_75t_L g6146 ( 
.A(n_4788),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_4993),
.Y(n_6147)
);

INVx2_ASAP7_75t_L g6148 ( 
.A(n_5317),
.Y(n_6148)
);

INVx2_ASAP7_75t_L g6149 ( 
.A(n_5317),
.Y(n_6149)
);

NAND2xp5_ASAP7_75t_L g6150 ( 
.A(n_5093),
.B(n_3312),
.Y(n_6150)
);

NOR2xp33_ASAP7_75t_SL g6151 ( 
.A(n_4975),
.B(n_3106),
.Y(n_6151)
);

BUFx6f_ASAP7_75t_L g6152 ( 
.A(n_4918),
.Y(n_6152)
);

INVx2_ASAP7_75t_L g6153 ( 
.A(n_5317),
.Y(n_6153)
);

NAND2xp5_ASAP7_75t_L g6154 ( 
.A(n_5093),
.B(n_3319),
.Y(n_6154)
);

BUFx6f_ASAP7_75t_L g6155 ( 
.A(n_4918),
.Y(n_6155)
);

AND2x4_ASAP7_75t_L g6156 ( 
.A(n_4718),
.B(n_3325),
.Y(n_6156)
);

BUFx6f_ASAP7_75t_L g6157 ( 
.A(n_4918),
.Y(n_6157)
);

INVx2_ASAP7_75t_L g6158 ( 
.A(n_5317),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_4993),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_4993),
.Y(n_6160)
);

OA21x2_ASAP7_75t_L g6161 ( 
.A1(n_5105),
.A2(n_3350),
.B(n_3338),
.Y(n_6161)
);

INVx2_ASAP7_75t_L g6162 ( 
.A(n_5317),
.Y(n_6162)
);

INVx2_ASAP7_75t_SL g6163 ( 
.A(n_4718),
.Y(n_6163)
);

INVx2_ASAP7_75t_L g6164 ( 
.A(n_5317),
.Y(n_6164)
);

AND2x2_ASAP7_75t_SL g6165 ( 
.A(n_4743),
.B(n_3227),
.Y(n_6165)
);

INVx3_ASAP7_75t_L g6166 ( 
.A(n_4918),
.Y(n_6166)
);

AND2x4_ASAP7_75t_L g6167 ( 
.A(n_4718),
.B(n_3351),
.Y(n_6167)
);

BUFx6f_ASAP7_75t_L g6168 ( 
.A(n_4918),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_4993),
.Y(n_6169)
);

BUFx6f_ASAP7_75t_L g6170 ( 
.A(n_4918),
.Y(n_6170)
);

NOR2xp33_ASAP7_75t_L g6171 ( 
.A(n_5093),
.B(n_3817),
.Y(n_6171)
);

BUFx8_ASAP7_75t_L g6172 ( 
.A(n_4835),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_4993),
.Y(n_6173)
);

NAND2xp5_ASAP7_75t_L g6174 ( 
.A(n_5093),
.B(n_3356),
.Y(n_6174)
);

INVx1_ASAP7_75t_L g6175 ( 
.A(n_4993),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_4993),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_4993),
.Y(n_6177)
);

INVx1_ASAP7_75t_L g6178 ( 
.A(n_4993),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_4993),
.Y(n_6179)
);

CKINVDCx11_ASAP7_75t_R g6180 ( 
.A(n_4992),
.Y(n_6180)
);

AND2x2_ASAP7_75t_SL g6181 ( 
.A(n_4743),
.B(n_3263),
.Y(n_6181)
);

BUFx6f_ASAP7_75t_L g6182 ( 
.A(n_4918),
.Y(n_6182)
);

AND2x4_ASAP7_75t_L g6183 ( 
.A(n_4718),
.B(n_3357),
.Y(n_6183)
);

NAND2xp5_ASAP7_75t_L g6184 ( 
.A(n_5093),
.B(n_3360),
.Y(n_6184)
);

AND2x4_ASAP7_75t_L g6185 ( 
.A(n_4718),
.B(n_3368),
.Y(n_6185)
);

AND2x2_ASAP7_75t_L g6186 ( 
.A(n_4970),
.B(n_3112),
.Y(n_6186)
);

CKINVDCx20_ASAP7_75t_R g6187 ( 
.A(n_4719),
.Y(n_6187)
);

AOI22xp5_ASAP7_75t_SL g6188 ( 
.A1(n_5405),
.A2(n_3116),
.B1(n_3119),
.B2(n_3113),
.Y(n_6188)
);

INVx5_ASAP7_75t_L g6189 ( 
.A(n_4788),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_4993),
.Y(n_6190)
);

AND2x2_ASAP7_75t_L g6191 ( 
.A(n_4970),
.B(n_3121),
.Y(n_6191)
);

CKINVDCx5p33_ASAP7_75t_R g6192 ( 
.A(n_4718),
.Y(n_6192)
);

XNOR2x2_ASAP7_75t_R g6193 ( 
.A(n_5944),
.B(n_3503),
.Y(n_6193)
);

AND2x4_ASAP7_75t_L g6194 ( 
.A(n_6163),
.B(n_3372),
.Y(n_6194)
);

INVx1_ASAP7_75t_L g6195 ( 
.A(n_5968),
.Y(n_6195)
);

INVx2_ASAP7_75t_L g6196 ( 
.A(n_5627),
.Y(n_6196)
);

INVx3_ASAP7_75t_L g6197 ( 
.A(n_5979),
.Y(n_6197)
);

INVx1_ASAP7_75t_L g6198 ( 
.A(n_6017),
.Y(n_6198)
);

NAND2xp5_ASAP7_75t_L g6199 ( 
.A(n_6186),
.B(n_3122),
.Y(n_6199)
);

INVx1_ASAP7_75t_L g6200 ( 
.A(n_5564),
.Y(n_6200)
);

AND2x2_ASAP7_75t_L g6201 ( 
.A(n_5448),
.B(n_3123),
.Y(n_6201)
);

INVx2_ASAP7_75t_L g6202 ( 
.A(n_5542),
.Y(n_6202)
);

INVx3_ASAP7_75t_L g6203 ( 
.A(n_5799),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_5582),
.Y(n_6204)
);

INVx2_ASAP7_75t_L g6205 ( 
.A(n_5552),
.Y(n_6205)
);

INVx2_ASAP7_75t_L g6206 ( 
.A(n_5554),
.Y(n_6206)
);

NAND2xp5_ASAP7_75t_L g6207 ( 
.A(n_6191),
.B(n_3127),
.Y(n_6207)
);

NAND2xp5_ASAP7_75t_SL g6208 ( 
.A(n_6151),
.B(n_3129),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_5589),
.Y(n_6209)
);

BUFx6f_ASAP7_75t_L g6210 ( 
.A(n_5438),
.Y(n_6210)
);

INVx3_ASAP7_75t_L g6211 ( 
.A(n_5935),
.Y(n_6211)
);

BUFx6f_ASAP7_75t_L g6212 ( 
.A(n_6123),
.Y(n_6212)
);

BUFx6f_ASAP7_75t_L g6213 ( 
.A(n_6143),
.Y(n_6213)
);

INVx2_ASAP7_75t_L g6214 ( 
.A(n_5563),
.Y(n_6214)
);

NAND2xp5_ASAP7_75t_L g6215 ( 
.A(n_5757),
.B(n_3130),
.Y(n_6215)
);

NAND2xp5_ASAP7_75t_SL g6216 ( 
.A(n_5732),
.B(n_3132),
.Y(n_6216)
);

INVx1_ASAP7_75t_L g6217 ( 
.A(n_5594),
.Y(n_6217)
);

AND2x2_ASAP7_75t_L g6218 ( 
.A(n_5429),
.B(n_3134),
.Y(n_6218)
);

OAI22xp5_ASAP7_75t_SL g6219 ( 
.A1(n_5745),
.A2(n_3142),
.B1(n_3144),
.B2(n_3140),
.Y(n_6219)
);

INVx2_ASAP7_75t_L g6220 ( 
.A(n_5567),
.Y(n_6220)
);

BUFx6f_ASAP7_75t_L g6221 ( 
.A(n_6152),
.Y(n_6221)
);

BUFx6f_ASAP7_75t_L g6222 ( 
.A(n_6155),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_5603),
.Y(n_6223)
);

AND2x4_ASAP7_75t_L g6224 ( 
.A(n_5426),
.B(n_3382),
.Y(n_6224)
);

INVx2_ASAP7_75t_L g6225 ( 
.A(n_5568),
.Y(n_6225)
);

AND2x6_ASAP7_75t_L g6226 ( 
.A(n_5676),
.B(n_3383),
.Y(n_6226)
);

BUFx6f_ASAP7_75t_L g6227 ( 
.A(n_6157),
.Y(n_6227)
);

INVxp67_ASAP7_75t_L g6228 ( 
.A(n_5481),
.Y(n_6228)
);

INVx3_ASAP7_75t_L g6229 ( 
.A(n_6122),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_5607),
.Y(n_6230)
);

NAND2xp5_ASAP7_75t_L g6231 ( 
.A(n_5464),
.B(n_3150),
.Y(n_6231)
);

OR2x2_ASAP7_75t_L g6232 ( 
.A(n_5733),
.B(n_3152),
.Y(n_6232)
);

NAND2xp5_ASAP7_75t_SL g6233 ( 
.A(n_5447),
.B(n_5715),
.Y(n_6233)
);

BUFx6f_ASAP7_75t_L g6234 ( 
.A(n_6168),
.Y(n_6234)
);

INVx3_ASAP7_75t_L g6235 ( 
.A(n_6127),
.Y(n_6235)
);

NAND2xp33_ASAP7_75t_L g6236 ( 
.A(n_5532),
.B(n_3155),
.Y(n_6236)
);

INVx2_ASAP7_75t_L g6237 ( 
.A(n_5571),
.Y(n_6237)
);

INVx2_ASAP7_75t_L g6238 ( 
.A(n_5583),
.Y(n_6238)
);

BUFx6f_ASAP7_75t_L g6239 ( 
.A(n_6170),
.Y(n_6239)
);

HB1xp67_ASAP7_75t_L g6240 ( 
.A(n_5620),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_5609),
.Y(n_6241)
);

INVx2_ASAP7_75t_L g6242 ( 
.A(n_5585),
.Y(n_6242)
);

INVx2_ASAP7_75t_L g6243 ( 
.A(n_5588),
.Y(n_6243)
);

AND2x4_ASAP7_75t_L g6244 ( 
.A(n_5435),
.B(n_3385),
.Y(n_6244)
);

INVx2_ASAP7_75t_L g6245 ( 
.A(n_5591),
.Y(n_6245)
);

BUFx8_ASAP7_75t_L g6246 ( 
.A(n_5578),
.Y(n_6246)
);

INVx2_ASAP7_75t_L g6247 ( 
.A(n_5596),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_5598),
.Y(n_6248)
);

XOR2xp5_ASAP7_75t_L g6249 ( 
.A(n_5520),
.B(n_3157),
.Y(n_6249)
);

INVx2_ASAP7_75t_L g6250 ( 
.A(n_5599),
.Y(n_6250)
);

BUFx6f_ASAP7_75t_L g6251 ( 
.A(n_6182),
.Y(n_6251)
);

CKINVDCx5p33_ASAP7_75t_R g6252 ( 
.A(n_5637),
.Y(n_6252)
);

AND2x2_ASAP7_75t_L g6253 ( 
.A(n_5846),
.B(n_3158),
.Y(n_6253)
);

INVx2_ASAP7_75t_L g6254 ( 
.A(n_5602),
.Y(n_6254)
);

NAND2xp33_ASAP7_75t_SL g6255 ( 
.A(n_5460),
.B(n_3162),
.Y(n_6255)
);

AND2x4_ASAP7_75t_L g6256 ( 
.A(n_6146),
.B(n_3388),
.Y(n_6256)
);

BUFx6f_ASAP7_75t_L g6257 ( 
.A(n_6189),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_5613),
.Y(n_6258)
);

NAND2xp5_ASAP7_75t_L g6259 ( 
.A(n_5917),
.B(n_3170),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_SL g6260 ( 
.A(n_5727),
.B(n_3174),
.Y(n_6260)
);

NAND2xp5_ASAP7_75t_L g6261 ( 
.A(n_5556),
.B(n_5923),
.Y(n_6261)
);

INVxp67_ASAP7_75t_L g6262 ( 
.A(n_5618),
.Y(n_6262)
);

INVx2_ASAP7_75t_L g6263 ( 
.A(n_5608),
.Y(n_6263)
);

INVx2_ASAP7_75t_L g6264 ( 
.A(n_5622),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5621),
.Y(n_6265)
);

OAI22xp5_ASAP7_75t_SL g6266 ( 
.A1(n_5746),
.A2(n_5767),
.B1(n_5815),
.B2(n_5761),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_5623),
.Y(n_6267)
);

INVx1_ASAP7_75t_L g6268 ( 
.A(n_5626),
.Y(n_6268)
);

OAI21x1_ASAP7_75t_L g6269 ( 
.A1(n_5428),
.A2(n_3270),
.B(n_3267),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_5651),
.Y(n_6270)
);

HB1xp67_ASAP7_75t_L g6271 ( 
.A(n_5450),
.Y(n_6271)
);

INVx2_ASAP7_75t_L g6272 ( 
.A(n_6041),
.Y(n_6272)
);

BUFx6f_ASAP7_75t_L g6273 ( 
.A(n_5471),
.Y(n_6273)
);

XOR2xp5_ASAP7_75t_L g6274 ( 
.A(n_5616),
.B(n_3175),
.Y(n_6274)
);

INVx2_ASAP7_75t_L g6275 ( 
.A(n_5982),
.Y(n_6275)
);

INVx3_ASAP7_75t_L g6276 ( 
.A(n_5662),
.Y(n_6276)
);

INVx1_ASAP7_75t_L g6277 ( 
.A(n_5652),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_5988),
.Y(n_6278)
);

INVx2_ASAP7_75t_L g6279 ( 
.A(n_5989),
.Y(n_6279)
);

INVx2_ASAP7_75t_L g6280 ( 
.A(n_5999),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_5672),
.Y(n_6281)
);

INVx3_ASAP7_75t_L g6282 ( 
.A(n_6142),
.Y(n_6282)
);

NAND2xp5_ASAP7_75t_L g6283 ( 
.A(n_6171),
.B(n_3176),
.Y(n_6283)
);

INVx2_ASAP7_75t_L g6284 ( 
.A(n_6002),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_5679),
.Y(n_6285)
);

CKINVDCx5p33_ASAP7_75t_R g6286 ( 
.A(n_5737),
.Y(n_6286)
);

AND2x6_ASAP7_75t_L g6287 ( 
.A(n_5719),
.B(n_3390),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_5682),
.Y(n_6288)
);

INVx3_ASAP7_75t_L g6289 ( 
.A(n_6192),
.Y(n_6289)
);

INVx1_ASAP7_75t_L g6290 ( 
.A(n_5686),
.Y(n_6290)
);

BUFx6f_ASAP7_75t_L g6291 ( 
.A(n_5474),
.Y(n_6291)
);

INVx2_ASAP7_75t_L g6292 ( 
.A(n_6005),
.Y(n_6292)
);

HB1xp67_ASAP7_75t_L g6293 ( 
.A(n_5533),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_5698),
.Y(n_6294)
);

BUFx6f_ASAP7_75t_L g6295 ( 
.A(n_5634),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_5707),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_5708),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_5717),
.Y(n_6298)
);

BUFx6f_ASAP7_75t_L g6299 ( 
.A(n_5634),
.Y(n_6299)
);

NAND2xp5_ASAP7_75t_L g6300 ( 
.A(n_5685),
.B(n_5793),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_5721),
.Y(n_6301)
);

NOR3xp33_ASAP7_75t_L g6302 ( 
.A(n_5996),
.B(n_3983),
.C(n_3964),
.Y(n_6302)
);

HB1xp67_ASAP7_75t_L g6303 ( 
.A(n_5509),
.Y(n_6303)
);

BUFx6f_ASAP7_75t_L g6304 ( 
.A(n_5771),
.Y(n_6304)
);

INVx2_ASAP7_75t_L g6305 ( 
.A(n_6011),
.Y(n_6305)
);

CKINVDCx16_ASAP7_75t_R g6306 ( 
.A(n_5463),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_5722),
.Y(n_6307)
);

CKINVDCx5p33_ASAP7_75t_R g6308 ( 
.A(n_5764),
.Y(n_6308)
);

HB1xp67_ASAP7_75t_L g6309 ( 
.A(n_5581),
.Y(n_6309)
);

INVx1_ASAP7_75t_L g6310 ( 
.A(n_5726),
.Y(n_6310)
);

INVx3_ASAP7_75t_L g6311 ( 
.A(n_6126),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_5741),
.Y(n_6312)
);

AND2x4_ASAP7_75t_L g6313 ( 
.A(n_5437),
.B(n_3394),
.Y(n_6313)
);

NAND2xp5_ASAP7_75t_L g6314 ( 
.A(n_5829),
.B(n_3182),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_5744),
.Y(n_6315)
);

BUFx6f_ASAP7_75t_L g6316 ( 
.A(n_5771),
.Y(n_6316)
);

INVx1_ASAP7_75t_L g6317 ( 
.A(n_5749),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_5754),
.Y(n_6318)
);

AND2x4_ASAP7_75t_L g6319 ( 
.A(n_5475),
.B(n_3398),
.Y(n_6319)
);

INVx2_ASAP7_75t_L g6320 ( 
.A(n_6013),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_5756),
.Y(n_6321)
);

AND2x2_ASAP7_75t_L g6322 ( 
.A(n_5484),
.B(n_5506),
.Y(n_6322)
);

INVx3_ASAP7_75t_L g6323 ( 
.A(n_6132),
.Y(n_6323)
);

AND2x2_ASAP7_75t_L g6324 ( 
.A(n_5530),
.B(n_3183),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_5776),
.Y(n_6325)
);

AND2x4_ASAP7_75t_L g6326 ( 
.A(n_6129),
.B(n_3404),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_5782),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_5789),
.Y(n_6328)
);

BUFx2_ASAP7_75t_L g6329 ( 
.A(n_6187),
.Y(n_6329)
);

BUFx6f_ASAP7_75t_L g6330 ( 
.A(n_6129),
.Y(n_6330)
);

INVx3_ASAP7_75t_L g6331 ( 
.A(n_6166),
.Y(n_6331)
);

INVx3_ASAP7_75t_L g6332 ( 
.A(n_5503),
.Y(n_6332)
);

AND2x2_ASAP7_75t_L g6333 ( 
.A(n_5671),
.B(n_3184),
.Y(n_6333)
);

INVxp67_ASAP7_75t_L g6334 ( 
.A(n_5888),
.Y(n_6334)
);

AND2x2_ASAP7_75t_L g6335 ( 
.A(n_5440),
.B(n_3186),
.Y(n_6335)
);

INVx2_ASAP7_75t_L g6336 ( 
.A(n_5427),
.Y(n_6336)
);

NAND2xp5_ASAP7_75t_L g6337 ( 
.A(n_5835),
.B(n_3187),
.Y(n_6337)
);

INVx1_ASAP7_75t_L g6338 ( 
.A(n_5796),
.Y(n_6338)
);

INVx2_ASAP7_75t_L g6339 ( 
.A(n_5443),
.Y(n_6339)
);

NAND2xp5_ASAP7_75t_L g6340 ( 
.A(n_5840),
.B(n_3189),
.Y(n_6340)
);

NOR2xp33_ASAP7_75t_L g6341 ( 
.A(n_6027),
.B(n_3190),
.Y(n_6341)
);

NAND2xp5_ASAP7_75t_L g6342 ( 
.A(n_5853),
.B(n_3192),
.Y(n_6342)
);

INVx1_ASAP7_75t_L g6343 ( 
.A(n_5798),
.Y(n_6343)
);

INVx2_ASAP7_75t_L g6344 ( 
.A(n_6128),
.Y(n_6344)
);

HB1xp67_ASAP7_75t_L g6345 ( 
.A(n_5595),
.Y(n_6345)
);

AND2x2_ASAP7_75t_L g6346 ( 
.A(n_5792),
.B(n_3194),
.Y(n_6346)
);

INVx2_ASAP7_75t_L g6347 ( 
.A(n_6130),
.Y(n_6347)
);

NAND2xp5_ASAP7_75t_L g6348 ( 
.A(n_5874),
.B(n_3197),
.Y(n_6348)
);

HB1xp67_ASAP7_75t_L g6349 ( 
.A(n_5601),
.Y(n_6349)
);

INVx2_ASAP7_75t_L g6350 ( 
.A(n_6133),
.Y(n_6350)
);

NAND2xp5_ASAP7_75t_L g6351 ( 
.A(n_5878),
.B(n_3200),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_5801),
.Y(n_6352)
);

INVx2_ASAP7_75t_L g6353 ( 
.A(n_6134),
.Y(n_6353)
);

BUFx2_ASAP7_75t_L g6354 ( 
.A(n_5924),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_5809),
.Y(n_6355)
);

INVx1_ASAP7_75t_L g6356 ( 
.A(n_5814),
.Y(n_6356)
);

NOR2xp33_ASAP7_75t_SL g6357 ( 
.A(n_6141),
.B(n_6018),
.Y(n_6357)
);

AND2x4_ASAP7_75t_L g6358 ( 
.A(n_5580),
.B(n_3406),
.Y(n_6358)
);

BUFx2_ASAP7_75t_L g6359 ( 
.A(n_5822),
.Y(n_6359)
);

NAND2xp5_ASAP7_75t_L g6360 ( 
.A(n_5898),
.B(n_3201),
.Y(n_6360)
);

INVx2_ASAP7_75t_L g6361 ( 
.A(n_6148),
.Y(n_6361)
);

AND2x6_ASAP7_75t_L g6362 ( 
.A(n_5436),
.B(n_3407),
.Y(n_6362)
);

AND2x2_ASAP7_75t_L g6363 ( 
.A(n_6125),
.B(n_3202),
.Y(n_6363)
);

AND2x2_ASAP7_75t_L g6364 ( 
.A(n_6131),
.B(n_3206),
.Y(n_6364)
);

INVx6_ASAP7_75t_L g6365 ( 
.A(n_6095),
.Y(n_6365)
);

INVx3_ASAP7_75t_L g6366 ( 
.A(n_6064),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_5817),
.Y(n_6367)
);

INVx2_ASAP7_75t_L g6368 ( 
.A(n_6149),
.Y(n_6368)
);

INVx1_ASAP7_75t_L g6369 ( 
.A(n_5820),
.Y(n_6369)
);

NAND2xp5_ASAP7_75t_SL g6370 ( 
.A(n_5772),
.B(n_3208),
.Y(n_6370)
);

INVx2_ASAP7_75t_L g6371 ( 
.A(n_6153),
.Y(n_6371)
);

NAND2xp5_ASAP7_75t_L g6372 ( 
.A(n_5899),
.B(n_3209),
.Y(n_6372)
);

INVx2_ASAP7_75t_L g6373 ( 
.A(n_6158),
.Y(n_6373)
);

INVx1_ASAP7_75t_L g6374 ( 
.A(n_5834),
.Y(n_6374)
);

BUFx2_ASAP7_75t_L g6375 ( 
.A(n_5863),
.Y(n_6375)
);

CKINVDCx20_ASAP7_75t_R g6376 ( 
.A(n_5439),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_5838),
.Y(n_6377)
);

NAND2xp5_ASAP7_75t_SL g6378 ( 
.A(n_5468),
.B(n_3210),
.Y(n_6378)
);

INVx1_ASAP7_75t_L g6379 ( 
.A(n_5842),
.Y(n_6379)
);

CKINVDCx20_ASAP7_75t_R g6380 ( 
.A(n_5454),
.Y(n_6380)
);

OA21x2_ASAP7_75t_L g6381 ( 
.A1(n_5674),
.A2(n_3423),
.B(n_3413),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_5850),
.Y(n_6382)
);

NAND2xp5_ASAP7_75t_SL g6383 ( 
.A(n_5499),
.B(n_3212),
.Y(n_6383)
);

NOR2xp33_ASAP7_75t_L g6384 ( 
.A(n_5430),
.B(n_3213),
.Y(n_6384)
);

NAND2xp5_ASAP7_75t_SL g6385 ( 
.A(n_5635),
.B(n_3219),
.Y(n_6385)
);

NAND2xp5_ASAP7_75t_L g6386 ( 
.A(n_5907),
.B(n_3220),
.Y(n_6386)
);

AND2x4_ASAP7_75t_L g6387 ( 
.A(n_5579),
.B(n_3426),
.Y(n_6387)
);

INVx1_ASAP7_75t_L g6388 ( 
.A(n_5866),
.Y(n_6388)
);

NAND2xp5_ASAP7_75t_L g6389 ( 
.A(n_5916),
.B(n_3222),
.Y(n_6389)
);

BUFx6f_ASAP7_75t_L g6390 ( 
.A(n_6071),
.Y(n_6390)
);

INVx2_ASAP7_75t_L g6391 ( 
.A(n_6162),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_5867),
.Y(n_6392)
);

INVx1_ASAP7_75t_L g6393 ( 
.A(n_5870),
.Y(n_6393)
);

INVx2_ASAP7_75t_L g6394 ( 
.A(n_6164),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_5886),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_5896),
.Y(n_6396)
);

AND2x4_ASAP7_75t_L g6397 ( 
.A(n_5903),
.B(n_3429),
.Y(n_6397)
);

BUFx6f_ASAP7_75t_L g6398 ( 
.A(n_5441),
.Y(n_6398)
);

AND2x4_ASAP7_75t_L g6399 ( 
.A(n_6070),
.B(n_3430),
.Y(n_6399)
);

INVx3_ASAP7_75t_L g6400 ( 
.A(n_6092),
.Y(n_6400)
);

INVx3_ASAP7_75t_L g6401 ( 
.A(n_5566),
.Y(n_6401)
);

BUFx6f_ASAP7_75t_L g6402 ( 
.A(n_5465),
.Y(n_6402)
);

HB1xp67_ASAP7_75t_L g6403 ( 
.A(n_5605),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_5902),
.Y(n_6404)
);

INVx1_ASAP7_75t_L g6405 ( 
.A(n_5905),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_5913),
.Y(n_6406)
);

INVx1_ASAP7_75t_L g6407 ( 
.A(n_5915),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_5920),
.Y(n_6408)
);

INVxp67_ASAP7_75t_L g6409 ( 
.A(n_5759),
.Y(n_6409)
);

OAI22xp5_ASAP7_75t_SL g6410 ( 
.A1(n_5538),
.A2(n_3224),
.B1(n_3225),
.B2(n_3223),
.Y(n_6410)
);

INVx2_ASAP7_75t_L g6411 ( 
.A(n_5861),
.Y(n_6411)
);

AND2x4_ASAP7_75t_L g6412 ( 
.A(n_5791),
.B(n_3432),
.Y(n_6412)
);

INVx3_ASAP7_75t_L g6413 ( 
.A(n_6121),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_5927),
.Y(n_6414)
);

NAND2xp5_ASAP7_75t_L g6415 ( 
.A(n_5929),
.B(n_3226),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_5930),
.Y(n_6416)
);

INVx2_ASAP7_75t_L g6417 ( 
.A(n_5631),
.Y(n_6417)
);

INVx1_ASAP7_75t_L g6418 ( 
.A(n_5939),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_5942),
.Y(n_6419)
);

INVx1_ASAP7_75t_L g6420 ( 
.A(n_5952),
.Y(n_6420)
);

INVx2_ASAP7_75t_L g6421 ( 
.A(n_5639),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_5964),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_5965),
.Y(n_6423)
);

NOR2xp33_ASAP7_75t_L g6424 ( 
.A(n_6037),
.B(n_3230),
.Y(n_6424)
);

AND2x4_ASAP7_75t_L g6425 ( 
.A(n_5791),
.B(n_5714),
.Y(n_6425)
);

INVx2_ASAP7_75t_L g6426 ( 
.A(n_5642),
.Y(n_6426)
);

INVx1_ASAP7_75t_L g6427 ( 
.A(n_5969),
.Y(n_6427)
);

AND2x2_ASAP7_75t_L g6428 ( 
.A(n_6156),
.B(n_3231),
.Y(n_6428)
);

INVx1_ASAP7_75t_L g6429 ( 
.A(n_5974),
.Y(n_6429)
);

NAND2xp5_ASAP7_75t_L g6430 ( 
.A(n_5934),
.B(n_3232),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_5986),
.Y(n_6431)
);

OAI22xp5_ASAP7_75t_SL g6432 ( 
.A1(n_5545),
.A2(n_3239),
.B1(n_3240),
.B2(n_3234),
.Y(n_6432)
);

INVx2_ASAP7_75t_L g6433 ( 
.A(n_5649),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_6008),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_6009),
.Y(n_6435)
);

INVx2_ASAP7_75t_L g6436 ( 
.A(n_5654),
.Y(n_6436)
);

INVx2_ASAP7_75t_L g6437 ( 
.A(n_5660),
.Y(n_6437)
);

INVx2_ASAP7_75t_L g6438 ( 
.A(n_5675),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6014),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_6019),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_6022),
.Y(n_6441)
);

NAND2xp5_ASAP7_75t_SL g6442 ( 
.A(n_5668),
.B(n_3242),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_6030),
.Y(n_6443)
);

HB1xp67_ASAP7_75t_L g6444 ( 
.A(n_5687),
.Y(n_6444)
);

INVx2_ASAP7_75t_L g6445 ( 
.A(n_5678),
.Y(n_6445)
);

INVx2_ASAP7_75t_L g6446 ( 
.A(n_5690),
.Y(n_6446)
);

INVx1_ASAP7_75t_L g6447 ( 
.A(n_5497),
.Y(n_6447)
);

INVx2_ASAP7_75t_L g6448 ( 
.A(n_5693),
.Y(n_6448)
);

HB1xp67_ASAP7_75t_L g6449 ( 
.A(n_5537),
.Y(n_6449)
);

HB1xp67_ASAP7_75t_L g6450 ( 
.A(n_5466),
.Y(n_6450)
);

BUFx3_ASAP7_75t_L g6451 ( 
.A(n_5688),
.Y(n_6451)
);

INVx1_ASAP7_75t_L g6452 ( 
.A(n_5498),
.Y(n_6452)
);

INVx1_ASAP7_75t_L g6453 ( 
.A(n_5502),
.Y(n_6453)
);

INVx2_ASAP7_75t_L g6454 ( 
.A(n_5696),
.Y(n_6454)
);

NAND2xp33_ASAP7_75t_L g6455 ( 
.A(n_5786),
.B(n_3250),
.Y(n_6455)
);

AND2x4_ASAP7_75t_L g6456 ( 
.A(n_5604),
.B(n_3438),
.Y(n_6456)
);

NAND2xp5_ASAP7_75t_L g6457 ( 
.A(n_5950),
.B(n_3252),
.Y(n_6457)
);

NAND2xp5_ASAP7_75t_L g6458 ( 
.A(n_5966),
.B(n_3255),
.Y(n_6458)
);

NAND2xp5_ASAP7_75t_L g6459 ( 
.A(n_5983),
.B(n_3258),
.Y(n_6459)
);

AND2x4_ASAP7_75t_L g6460 ( 
.A(n_5628),
.B(n_3450),
.Y(n_6460)
);

INVx2_ASAP7_75t_L g6461 ( 
.A(n_5700),
.Y(n_6461)
);

NAND2xp5_ASAP7_75t_L g6462 ( 
.A(n_6004),
.B(n_3259),
.Y(n_6462)
);

INVx2_ASAP7_75t_L g6463 ( 
.A(n_5704),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_5514),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_5516),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_5519),
.Y(n_6466)
);

NOR2xp33_ASAP7_75t_L g6467 ( 
.A(n_5943),
.B(n_3260),
.Y(n_6467)
);

CKINVDCx8_ASAP7_75t_R g6468 ( 
.A(n_5683),
.Y(n_6468)
);

CKINVDCx8_ASAP7_75t_R g6469 ( 
.A(n_5849),
.Y(n_6469)
);

INVxp67_ASAP7_75t_L g6470 ( 
.A(n_5783),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_5525),
.Y(n_6471)
);

INVx1_ASAP7_75t_SL g6472 ( 
.A(n_5755),
.Y(n_6472)
);

HB1xp67_ASAP7_75t_L g6473 ( 
.A(n_5641),
.Y(n_6473)
);

NAND2xp33_ASAP7_75t_L g6474 ( 
.A(n_5875),
.B(n_5926),
.Y(n_6474)
);

BUFx2_ASAP7_75t_L g6475 ( 
.A(n_6115),
.Y(n_6475)
);

INVx1_ASAP7_75t_L g6476 ( 
.A(n_5531),
.Y(n_6476)
);

NAND2x1p5_ASAP7_75t_L g6477 ( 
.A(n_5827),
.B(n_3460),
.Y(n_6477)
);

INVx1_ASAP7_75t_L g6478 ( 
.A(n_5536),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_5539),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_5543),
.Y(n_6480)
);

INVx1_ASAP7_75t_L g6481 ( 
.A(n_5553),
.Y(n_6481)
);

INVx2_ASAP7_75t_L g6482 ( 
.A(n_5706),
.Y(n_6482)
);

BUFx6f_ASAP7_75t_L g6483 ( 
.A(n_5479),
.Y(n_6483)
);

INVx2_ASAP7_75t_L g6484 ( 
.A(n_5709),
.Y(n_6484)
);

NAND2xp5_ASAP7_75t_L g6485 ( 
.A(n_6034),
.B(n_3264),
.Y(n_6485)
);

INVx1_ASAP7_75t_L g6486 ( 
.A(n_5555),
.Y(n_6486)
);

INVx2_ASAP7_75t_L g6487 ( 
.A(n_5712),
.Y(n_6487)
);

BUFx8_ASAP7_75t_L g6488 ( 
.A(n_5615),
.Y(n_6488)
);

NAND2xp33_ASAP7_75t_SL g6489 ( 
.A(n_5919),
.B(n_3265),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_5558),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_5462),
.Y(n_6491)
);

CKINVDCx20_ASAP7_75t_R g6492 ( 
.A(n_5495),
.Y(n_6492)
);

INVx1_ASAP7_75t_L g6493 ( 
.A(n_5467),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_5470),
.Y(n_6494)
);

NOR2xp33_ASAP7_75t_L g6495 ( 
.A(n_5758),
.B(n_5882),
.Y(n_6495)
);

NAND2xp5_ASAP7_75t_L g6496 ( 
.A(n_6150),
.B(n_3266),
.Y(n_6496)
);

AND2x2_ASAP7_75t_L g6497 ( 
.A(n_6167),
.B(n_3268),
.Y(n_6497)
);

AND2x4_ASAP7_75t_L g6498 ( 
.A(n_5720),
.B(n_3462),
.Y(n_6498)
);

AND2x2_ASAP7_75t_L g6499 ( 
.A(n_6183),
.B(n_3271),
.Y(n_6499)
);

INVx2_ASAP7_75t_L g6500 ( 
.A(n_5713),
.Y(n_6500)
);

NAND2xp5_ASAP7_75t_L g6501 ( 
.A(n_6154),
.B(n_3275),
.Y(n_6501)
);

INVx3_ASAP7_75t_L g6502 ( 
.A(n_5487),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_5472),
.Y(n_6503)
);

INVx3_ASAP7_75t_L g6504 ( 
.A(n_5513),
.Y(n_6504)
);

INVx1_ASAP7_75t_L g6505 ( 
.A(n_5473),
.Y(n_6505)
);

INVx2_ASAP7_75t_L g6506 ( 
.A(n_5729),
.Y(n_6506)
);

INVx2_ASAP7_75t_L g6507 ( 
.A(n_5730),
.Y(n_6507)
);

NAND2xp5_ASAP7_75t_L g6508 ( 
.A(n_6174),
.B(n_3277),
.Y(n_6508)
);

AND2x6_ASAP7_75t_L g6509 ( 
.A(n_5445),
.B(n_3465),
.Y(n_6509)
);

NAND2xp5_ASAP7_75t_L g6510 ( 
.A(n_6184),
.B(n_3278),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_5477),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_5485),
.Y(n_6512)
);

NAND2xp5_ASAP7_75t_L g6513 ( 
.A(n_5584),
.B(n_3280),
.Y(n_6513)
);

AND2x2_ASAP7_75t_L g6514 ( 
.A(n_6185),
.B(n_3292),
.Y(n_6514)
);

NAND2xp5_ASAP7_75t_L g6515 ( 
.A(n_5611),
.B(n_3294),
.Y(n_6515)
);

INVx1_ASAP7_75t_L g6516 ( 
.A(n_5491),
.Y(n_6516)
);

INVx1_ASAP7_75t_L g6517 ( 
.A(n_5494),
.Y(n_6517)
);

INVx2_ASAP7_75t_L g6518 ( 
.A(n_5734),
.Y(n_6518)
);

INVx3_ASAP7_75t_L g6519 ( 
.A(n_5997),
.Y(n_6519)
);

AND2x4_ASAP7_75t_L g6520 ( 
.A(n_5743),
.B(n_3467),
.Y(n_6520)
);

INVx1_ASAP7_75t_L g6521 ( 
.A(n_6046),
.Y(n_6521)
);

INVx1_ASAP7_75t_L g6522 ( 
.A(n_5735),
.Y(n_6522)
);

AND2x2_ASAP7_75t_L g6523 ( 
.A(n_5551),
.B(n_3295),
.Y(n_6523)
);

INVx2_ASAP7_75t_L g6524 ( 
.A(n_5738),
.Y(n_6524)
);

INVx2_ASAP7_75t_L g6525 ( 
.A(n_5739),
.Y(n_6525)
);

BUFx2_ASAP7_75t_L g6526 ( 
.A(n_5806),
.Y(n_6526)
);

OAI21x1_ASAP7_75t_L g6527 ( 
.A1(n_5790),
.A2(n_3305),
.B(n_3273),
.Y(n_6527)
);

NOR2xp33_ASAP7_75t_L g6528 ( 
.A(n_5918),
.B(n_3297),
.Y(n_6528)
);

AND2x4_ASAP7_75t_L g6529 ( 
.A(n_5890),
.B(n_3468),
.Y(n_6529)
);

AND2x4_ASAP7_75t_L g6530 ( 
.A(n_5954),
.B(n_3471),
.Y(n_6530)
);

NAND2xp5_ASAP7_75t_L g6531 ( 
.A(n_5647),
.B(n_3298),
.Y(n_6531)
);

NAND2xp33_ASAP7_75t_L g6532 ( 
.A(n_5932),
.B(n_3301),
.Y(n_6532)
);

INVx2_ASAP7_75t_L g6533 ( 
.A(n_5747),
.Y(n_6533)
);

INVxp67_ASAP7_75t_L g6534 ( 
.A(n_5684),
.Y(n_6534)
);

NAND2xp33_ASAP7_75t_SL g6535 ( 
.A(n_5971),
.B(n_3302),
.Y(n_6535)
);

INVx2_ASAP7_75t_L g6536 ( 
.A(n_5751),
.Y(n_6536)
);

INVx4_ASAP7_75t_L g6537 ( 
.A(n_5725),
.Y(n_6537)
);

HB1xp67_ASAP7_75t_L g6538 ( 
.A(n_5963),
.Y(n_6538)
);

NAND2xp5_ASAP7_75t_L g6539 ( 
.A(n_5663),
.B(n_3308),
.Y(n_6539)
);

OA21x2_ASAP7_75t_L g6540 ( 
.A1(n_5880),
.A2(n_3479),
.B(n_3475),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_5766),
.Y(n_6541)
);

INVx1_ASAP7_75t_L g6542 ( 
.A(n_5770),
.Y(n_6542)
);

INVx2_ASAP7_75t_L g6543 ( 
.A(n_5773),
.Y(n_6543)
);

BUFx6f_ASAP7_75t_L g6544 ( 
.A(n_6136),
.Y(n_6544)
);

BUFx6f_ASAP7_75t_L g6545 ( 
.A(n_5994),
.Y(n_6545)
);

NAND2xp5_ASAP7_75t_L g6546 ( 
.A(n_5453),
.B(n_5496),
.Y(n_6546)
);

INVx1_ASAP7_75t_L g6547 ( 
.A(n_5785),
.Y(n_6547)
);

BUFx6f_ASAP7_75t_L g6548 ( 
.A(n_6007),
.Y(n_6548)
);

INVx2_ASAP7_75t_L g6549 ( 
.A(n_5804),
.Y(n_6549)
);

INVx1_ASAP7_75t_L g6550 ( 
.A(n_5816),
.Y(n_6550)
);

AND2x2_ASAP7_75t_L g6551 ( 
.A(n_5505),
.B(n_3309),
.Y(n_6551)
);

BUFx6f_ASAP7_75t_L g6552 ( 
.A(n_6020),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_5830),
.Y(n_6553)
);

NAND2xp5_ASAP7_75t_SL g6554 ( 
.A(n_6043),
.B(n_3316),
.Y(n_6554)
);

BUFx8_ASAP7_75t_L g6555 ( 
.A(n_5646),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_5832),
.Y(n_6556)
);

OAI21x1_ASAP7_75t_L g6557 ( 
.A1(n_5852),
.A2(n_3362),
.B(n_3329),
.Y(n_6557)
);

NAND2xp5_ASAP7_75t_SL g6558 ( 
.A(n_6067),
.B(n_3317),
.Y(n_6558)
);

OAI22xp5_ASAP7_75t_L g6559 ( 
.A1(n_5446),
.A2(n_3320),
.B1(n_3322),
.B2(n_3318),
.Y(n_6559)
);

HB1xp67_ASAP7_75t_L g6560 ( 
.A(n_5653),
.Y(n_6560)
);

AND2x2_ASAP7_75t_L g6561 ( 
.A(n_5508),
.B(n_3323),
.Y(n_6561)
);

INVx2_ASAP7_75t_L g6562 ( 
.A(n_5836),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_5837),
.Y(n_6563)
);

NAND2xp5_ASAP7_75t_SL g6564 ( 
.A(n_5931),
.B(n_3324),
.Y(n_6564)
);

INVx1_ASAP7_75t_L g6565 ( 
.A(n_5841),
.Y(n_6565)
);

HB1xp67_ASAP7_75t_L g6566 ( 
.A(n_5825),
.Y(n_6566)
);

HB1xp67_ASAP7_75t_L g6567 ( 
.A(n_5839),
.Y(n_6567)
);

AND2x4_ASAP7_75t_L g6568 ( 
.A(n_5625),
.B(n_3480),
.Y(n_6568)
);

NOR2x1_ASAP7_75t_L g6569 ( 
.A(n_6094),
.B(n_3481),
.Y(n_6569)
);

INVx2_ASAP7_75t_L g6570 ( 
.A(n_5843),
.Y(n_6570)
);

BUFx2_ASAP7_75t_L g6571 ( 
.A(n_5891),
.Y(n_6571)
);

INVx1_ASAP7_75t_L g6572 ( 
.A(n_5844),
.Y(n_6572)
);

BUFx2_ASAP7_75t_L g6573 ( 
.A(n_5940),
.Y(n_6573)
);

BUFx3_ASAP7_75t_L g6574 ( 
.A(n_5855),
.Y(n_6574)
);

INVx2_ASAP7_75t_L g6575 ( 
.A(n_5848),
.Y(n_6575)
);

HB1xp67_ASAP7_75t_L g6576 ( 
.A(n_5955),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_5857),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_5859),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_5862),
.Y(n_6579)
);

AND2x2_ASAP7_75t_L g6580 ( 
.A(n_5619),
.B(n_3327),
.Y(n_6580)
);

INVx1_ASAP7_75t_L g6581 ( 
.A(n_5864),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_5869),
.Y(n_6582)
);

BUFx6f_ASAP7_75t_L g6583 ( 
.A(n_6021),
.Y(n_6583)
);

INVx1_ASAP7_75t_L g6584 ( 
.A(n_5872),
.Y(n_6584)
);

INVx1_ASAP7_75t_L g6585 ( 
.A(n_5881),
.Y(n_6585)
);

INVx1_ASAP7_75t_L g6586 ( 
.A(n_5884),
.Y(n_6586)
);

OR2x2_ASAP7_75t_L g6587 ( 
.A(n_6100),
.B(n_3328),
.Y(n_6587)
);

NAND2xp5_ASAP7_75t_SL g6588 ( 
.A(n_5958),
.B(n_3330),
.Y(n_6588)
);

INVx2_ASAP7_75t_L g6589 ( 
.A(n_5887),
.Y(n_6589)
);

INVx2_ASAP7_75t_L g6590 ( 
.A(n_5889),
.Y(n_6590)
);

INVx1_ASAP7_75t_L g6591 ( 
.A(n_5893),
.Y(n_6591)
);

INVx3_ASAP7_75t_L g6592 ( 
.A(n_5667),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_5894),
.Y(n_6593)
);

AND2x2_ASAP7_75t_L g6594 ( 
.A(n_5576),
.B(n_3331),
.Y(n_6594)
);

HB1xp67_ASAP7_75t_L g6595 ( 
.A(n_5977),
.Y(n_6595)
);

INVx2_ASAP7_75t_L g6596 ( 
.A(n_5901),
.Y(n_6596)
);

INVx1_ASAP7_75t_L g6597 ( 
.A(n_5911),
.Y(n_6597)
);

BUFx6f_ASAP7_75t_L g6598 ( 
.A(n_6026),
.Y(n_6598)
);

AND2x2_ASAP7_75t_L g6599 ( 
.A(n_5624),
.B(n_3332),
.Y(n_6599)
);

INVx1_ASAP7_75t_L g6600 ( 
.A(n_5921),
.Y(n_6600)
);

INVx2_ASAP7_75t_L g6601 ( 
.A(n_5947),
.Y(n_6601)
);

INVx1_ASAP7_75t_L g6602 ( 
.A(n_5949),
.Y(n_6602)
);

INVx1_ASAP7_75t_L g6603 ( 
.A(n_5951),
.Y(n_6603)
);

INVx1_ASAP7_75t_L g6604 ( 
.A(n_5973),
.Y(n_6604)
);

INVx1_ASAP7_75t_L g6605 ( 
.A(n_5972),
.Y(n_6605)
);

BUFx6f_ASAP7_75t_L g6606 ( 
.A(n_6031),
.Y(n_6606)
);

INVx1_ASAP7_75t_L g6607 ( 
.A(n_5768),
.Y(n_6607)
);

INVx2_ASAP7_75t_L g6608 ( 
.A(n_5541),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_6036),
.Y(n_6609)
);

INVx1_ASAP7_75t_L g6610 ( 
.A(n_6042),
.Y(n_6610)
);

INVx1_ASAP7_75t_L g6611 ( 
.A(n_5710),
.Y(n_6611)
);

INVx1_ASAP7_75t_L g6612 ( 
.A(n_5723),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_5753),
.Y(n_6613)
);

NAND2xp5_ASAP7_75t_L g6614 ( 
.A(n_5432),
.B(n_3333),
.Y(n_6614)
);

BUFx6f_ASAP7_75t_L g6615 ( 
.A(n_6033),
.Y(n_6615)
);

NAND2xp5_ASAP7_75t_L g6616 ( 
.A(n_5517),
.B(n_3335),
.Y(n_6616)
);

BUFx2_ASAP7_75t_L g6617 ( 
.A(n_5978),
.Y(n_6617)
);

INVx3_ASAP7_75t_L g6618 ( 
.A(n_5669),
.Y(n_6618)
);

NAND2xp5_ASAP7_75t_L g6619 ( 
.A(n_5587),
.B(n_3336),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_5760),
.Y(n_6620)
);

NAND2xp5_ASAP7_75t_L g6621 ( 
.A(n_5633),
.B(n_3341),
.Y(n_6621)
);

INVx2_ASAP7_75t_L g6622 ( 
.A(n_5478),
.Y(n_6622)
);

BUFx6f_ASAP7_75t_L g6623 ( 
.A(n_6035),
.Y(n_6623)
);

INVx5_ASAP7_75t_L g6624 ( 
.A(n_6038),
.Y(n_6624)
);

NAND2xp33_ASAP7_75t_SL g6625 ( 
.A(n_5569),
.B(n_6015),
.Y(n_6625)
);

AND2x2_ASAP7_75t_L g6626 ( 
.A(n_5632),
.B(n_3342),
.Y(n_6626)
);

INVx2_ASAP7_75t_L g6627 ( 
.A(n_5486),
.Y(n_6627)
);

BUFx6f_ASAP7_75t_L g6628 ( 
.A(n_6044),
.Y(n_6628)
);

INVx1_ASAP7_75t_SL g6629 ( 
.A(n_5535),
.Y(n_6629)
);

NAND2xp5_ASAP7_75t_L g6630 ( 
.A(n_5665),
.B(n_3343),
.Y(n_6630)
);

BUFx6f_ASAP7_75t_L g6631 ( 
.A(n_6047),
.Y(n_6631)
);

AND2x4_ASAP7_75t_L g6632 ( 
.A(n_5701),
.B(n_3486),
.Y(n_6632)
);

OAI21x1_ASAP7_75t_L g6633 ( 
.A1(n_5858),
.A2(n_3396),
.B(n_3374),
.Y(n_6633)
);

NAND2xp5_ASAP7_75t_L g6634 ( 
.A(n_5945),
.B(n_3344),
.Y(n_6634)
);

INVx2_ASAP7_75t_L g6635 ( 
.A(n_5522),
.Y(n_6635)
);

HB1xp67_ASAP7_75t_L g6636 ( 
.A(n_6000),
.Y(n_6636)
);

AND2x2_ASAP7_75t_L g6637 ( 
.A(n_5661),
.B(n_3345),
.Y(n_6637)
);

INVx2_ASAP7_75t_L g6638 ( 
.A(n_5534),
.Y(n_6638)
);

INVx2_ASAP7_75t_L g6639 ( 
.A(n_5976),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_5805),
.Y(n_6640)
);

INVx1_ASAP7_75t_L g6641 ( 
.A(n_5811),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_5828),
.Y(n_6642)
);

AND2x4_ASAP7_75t_L g6643 ( 
.A(n_6063),
.B(n_3489),
.Y(n_6643)
);

INVx2_ASAP7_75t_L g6644 ( 
.A(n_6045),
.Y(n_6644)
);

BUFx6f_ASAP7_75t_L g6645 ( 
.A(n_6049),
.Y(n_6645)
);

INVx2_ASAP7_75t_L g6646 ( 
.A(n_5433),
.Y(n_6646)
);

INVx1_ASAP7_75t_SL g6647 ( 
.A(n_5980),
.Y(n_6647)
);

INVx2_ASAP7_75t_L g6648 ( 
.A(n_5459),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_5831),
.Y(n_6649)
);

AND2x2_ASAP7_75t_L g6650 ( 
.A(n_5544),
.B(n_3346),
.Y(n_6650)
);

NOR2xp33_ASAP7_75t_L g6651 ( 
.A(n_5664),
.B(n_3347),
.Y(n_6651)
);

HB1xp67_ASAP7_75t_L g6652 ( 
.A(n_5512),
.Y(n_6652)
);

INVxp67_ASAP7_75t_L g6653 ( 
.A(n_5897),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_5851),
.Y(n_6654)
);

INVx1_ASAP7_75t_L g6655 ( 
.A(n_5854),
.Y(n_6655)
);

HB1xp67_ASAP7_75t_L g6656 ( 
.A(n_5521),
.Y(n_6656)
);

INVx1_ASAP7_75t_L g6657 ( 
.A(n_5657),
.Y(n_6657)
);

AND2x2_ASAP7_75t_L g6658 ( 
.A(n_5909),
.B(n_3348),
.Y(n_6658)
);

BUFx8_ASAP7_75t_L g6659 ( 
.A(n_6057),
.Y(n_6659)
);

INVx1_ASAP7_75t_SL g6660 ( 
.A(n_6039),
.Y(n_6660)
);

INVx1_ASAP7_75t_L g6661 ( 
.A(n_5981),
.Y(n_6661)
);

INVx2_ASAP7_75t_L g6662 ( 
.A(n_6135),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_5985),
.Y(n_6663)
);

BUFx6f_ASAP7_75t_L g6664 ( 
.A(n_6059),
.Y(n_6664)
);

AND2x2_ASAP7_75t_L g6665 ( 
.A(n_6048),
.B(n_3349),
.Y(n_6665)
);

INVxp67_ASAP7_75t_L g6666 ( 
.A(n_5962),
.Y(n_6666)
);

INVx2_ASAP7_75t_L g6667 ( 
.A(n_6138),
.Y(n_6667)
);

NAND2xp5_ASAP7_75t_L g6668 ( 
.A(n_5948),
.B(n_3354),
.Y(n_6668)
);

AND2x2_ASAP7_75t_L g6669 ( 
.A(n_6061),
.B(n_3358),
.Y(n_6669)
);

AND2x2_ASAP7_75t_L g6670 ( 
.A(n_6078),
.B(n_5702),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_5987),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_6001),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_6140),
.Y(n_6673)
);

INVx1_ASAP7_75t_L g6674 ( 
.A(n_6024),
.Y(n_6674)
);

INVx2_ASAP7_75t_L g6675 ( 
.A(n_6144),
.Y(n_6675)
);

INVx2_ASAP7_75t_L g6676 ( 
.A(n_6145),
.Y(n_6676)
);

INVx1_ASAP7_75t_L g6677 ( 
.A(n_5910),
.Y(n_6677)
);

BUFx6f_ASAP7_75t_L g6678 ( 
.A(n_6073),
.Y(n_6678)
);

INVx1_ASAP7_75t_L g6679 ( 
.A(n_5787),
.Y(n_6679)
);

INVx1_ASAP7_75t_L g6680 ( 
.A(n_5800),
.Y(n_6680)
);

BUFx2_ASAP7_75t_L g6681 ( 
.A(n_6016),
.Y(n_6681)
);

INVx2_ASAP7_75t_L g6682 ( 
.A(n_6147),
.Y(n_6682)
);

INVx2_ASAP7_75t_L g6683 ( 
.A(n_6159),
.Y(n_6683)
);

HB1xp67_ASAP7_75t_L g6684 ( 
.A(n_6106),
.Y(n_6684)
);

INVx3_ASAP7_75t_L g6685 ( 
.A(n_5680),
.Y(n_6685)
);

INVx2_ASAP7_75t_L g6686 ( 
.A(n_6160),
.Y(n_6686)
);

INVx3_ASAP7_75t_L g6687 ( 
.A(n_5692),
.Y(n_6687)
);

AND2x2_ASAP7_75t_L g6688 ( 
.A(n_5795),
.B(n_3361),
.Y(n_6688)
);

INVx3_ASAP7_75t_L g6689 ( 
.A(n_5705),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_5873),
.Y(n_6690)
);

NAND2xp5_ASAP7_75t_L g6691 ( 
.A(n_5953),
.B(n_5961),
.Y(n_6691)
);

NAND2xp5_ASAP7_75t_SL g6692 ( 
.A(n_6090),
.B(n_6087),
.Y(n_6692)
);

AND2x4_ASAP7_75t_L g6693 ( 
.A(n_6075),
.B(n_3495),
.Y(n_6693)
);

NAND2xp5_ASAP7_75t_SL g6694 ( 
.A(n_6096),
.B(n_3363),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_5991),
.Y(n_6695)
);

NAND2xp5_ASAP7_75t_L g6696 ( 
.A(n_6055),
.B(n_3364),
.Y(n_6696)
);

BUFx6f_ASAP7_75t_L g6697 ( 
.A(n_6086),
.Y(n_6697)
);

INVx1_ASAP7_75t_L g6698 ( 
.A(n_5925),
.Y(n_6698)
);

HB1xp67_ASAP7_75t_L g6699 ( 
.A(n_6112),
.Y(n_6699)
);

INVx2_ASAP7_75t_L g6700 ( 
.A(n_6169),
.Y(n_6700)
);

INVx1_ASAP7_75t_L g6701 ( 
.A(n_6012),
.Y(n_6701)
);

BUFx6f_ASAP7_75t_L g6702 ( 
.A(n_6180),
.Y(n_6702)
);

INVx1_ASAP7_75t_L g6703 ( 
.A(n_6173),
.Y(n_6703)
);

NOR2xp33_ASAP7_75t_L g6704 ( 
.A(n_5826),
.B(n_3365),
.Y(n_6704)
);

INVx2_ASAP7_75t_L g6705 ( 
.A(n_6175),
.Y(n_6705)
);

INVx3_ASAP7_75t_L g6706 ( 
.A(n_5728),
.Y(n_6706)
);

INVx1_ASAP7_75t_L g6707 ( 
.A(n_6176),
.Y(n_6707)
);

INVx1_ASAP7_75t_L g6708 ( 
.A(n_6177),
.Y(n_6708)
);

HB1xp67_ASAP7_75t_L g6709 ( 
.A(n_6120),
.Y(n_6709)
);

INVx1_ASAP7_75t_L g6710 ( 
.A(n_6178),
.Y(n_6710)
);

AND2x4_ASAP7_75t_L g6711 ( 
.A(n_6054),
.B(n_3498),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_6179),
.Y(n_6712)
);

INVx1_ASAP7_75t_L g6713 ( 
.A(n_6190),
.Y(n_6713)
);

INVx2_ASAP7_75t_L g6714 ( 
.A(n_5451),
.Y(n_6714)
);

INVx2_ASAP7_75t_L g6715 ( 
.A(n_5452),
.Y(n_6715)
);

INVx2_ASAP7_75t_L g6716 ( 
.A(n_5456),
.Y(n_6716)
);

INVx3_ASAP7_75t_L g6717 ( 
.A(n_5480),
.Y(n_6717)
);

INVx1_ASAP7_75t_L g6718 ( 
.A(n_5500),
.Y(n_6718)
);

INVx3_ASAP7_75t_L g6719 ( 
.A(n_5483),
.Y(n_6719)
);

INVx2_ASAP7_75t_L g6720 ( 
.A(n_5461),
.Y(n_6720)
);

AND2x2_ASAP7_75t_L g6721 ( 
.A(n_5807),
.B(n_5808),
.Y(n_6721)
);

BUFx6f_ASAP7_75t_L g6722 ( 
.A(n_5490),
.Y(n_6722)
);

INVx1_ASAP7_75t_L g6723 ( 
.A(n_5504),
.Y(n_6723)
);

NAND2xp5_ASAP7_75t_L g6724 ( 
.A(n_5557),
.B(n_3366),
.Y(n_6724)
);

AOI22xp5_ASAP7_75t_L g6725 ( 
.A1(n_5515),
.A2(n_3367),
.B1(n_3371),
.B2(n_3369),
.Y(n_6725)
);

OA21x2_ASAP7_75t_L g6726 ( 
.A1(n_5914),
.A2(n_3514),
.B(n_3501),
.Y(n_6726)
);

AND2x2_ASAP7_75t_L g6727 ( 
.A(n_5812),
.B(n_5813),
.Y(n_6727)
);

BUFx6f_ASAP7_75t_L g6728 ( 
.A(n_5492),
.Y(n_6728)
);

BUFx6f_ASAP7_75t_L g6729 ( 
.A(n_5518),
.Y(n_6729)
);

BUFx8_ASAP7_75t_L g6730 ( 
.A(n_6101),
.Y(n_6730)
);

INVx1_ASAP7_75t_L g6731 ( 
.A(n_5511),
.Y(n_6731)
);

NAND2xp5_ASAP7_75t_L g6732 ( 
.A(n_5561),
.B(n_3373),
.Y(n_6732)
);

BUFx2_ASAP7_75t_L g6733 ( 
.A(n_6084),
.Y(n_6733)
);

INVx2_ASAP7_75t_L g6734 ( 
.A(n_5748),
.Y(n_6734)
);

BUFx6f_ASAP7_75t_L g6735 ( 
.A(n_5523),
.Y(n_6735)
);

INVx1_ASAP7_75t_L g6736 ( 
.A(n_5529),
.Y(n_6736)
);

CKINVDCx5p33_ASAP7_75t_R g6737 ( 
.A(n_6093),
.Y(n_6737)
);

INVx2_ASAP7_75t_L g6738 ( 
.A(n_5752),
.Y(n_6738)
);

INVx1_ASAP7_75t_L g6739 ( 
.A(n_5540),
.Y(n_6739)
);

INVx1_ASAP7_75t_L g6740 ( 
.A(n_5549),
.Y(n_6740)
);

OA21x2_ASAP7_75t_L g6741 ( 
.A1(n_5957),
.A2(n_3517),
.B(n_3516),
.Y(n_6741)
);

NAND2xp5_ASAP7_75t_L g6742 ( 
.A(n_5562),
.B(n_3376),
.Y(n_6742)
);

NAND2xp5_ASAP7_75t_L g6743 ( 
.A(n_5644),
.B(n_3387),
.Y(n_6743)
);

INVx1_ASAP7_75t_L g6744 ( 
.A(n_5575),
.Y(n_6744)
);

NAND2xp5_ASAP7_75t_SL g6745 ( 
.A(n_5856),
.B(n_3389),
.Y(n_6745)
);

INVx1_ASAP7_75t_L g6746 ( 
.A(n_5592),
.Y(n_6746)
);

INVx2_ASAP7_75t_L g6747 ( 
.A(n_5763),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_5769),
.Y(n_6748)
);

INVx1_ASAP7_75t_L g6749 ( 
.A(n_5600),
.Y(n_6749)
);

INVx4_ASAP7_75t_L g6750 ( 
.A(n_6003),
.Y(n_6750)
);

INVx3_ASAP7_75t_L g6751 ( 
.A(n_5526),
.Y(n_6751)
);

INVx3_ASAP7_75t_L g6752 ( 
.A(n_5565),
.Y(n_6752)
);

NAND2xp5_ASAP7_75t_SL g6753 ( 
.A(n_5868),
.B(n_3391),
.Y(n_6753)
);

BUFx6f_ASAP7_75t_L g6754 ( 
.A(n_5573),
.Y(n_6754)
);

INVx1_ASAP7_75t_L g6755 ( 
.A(n_5610),
.Y(n_6755)
);

INVx2_ASAP7_75t_L g6756 ( 
.A(n_5774),
.Y(n_6756)
);

INVx1_ASAP7_75t_L g6757 ( 
.A(n_5614),
.Y(n_6757)
);

AND2x2_ASAP7_75t_L g6758 ( 
.A(n_5833),
.B(n_3393),
.Y(n_6758)
);

INVx1_ASAP7_75t_L g6759 ( 
.A(n_5645),
.Y(n_6759)
);

HB1xp67_ASAP7_75t_L g6760 ( 
.A(n_6111),
.Y(n_6760)
);

INVxp67_ASAP7_75t_L g6761 ( 
.A(n_5998),
.Y(n_6761)
);

INVx2_ASAP7_75t_L g6762 ( 
.A(n_5780),
.Y(n_6762)
);

AND2x2_ASAP7_75t_L g6763 ( 
.A(n_5777),
.B(n_3395),
.Y(n_6763)
);

INVx2_ASAP7_75t_L g6764 ( 
.A(n_5781),
.Y(n_6764)
);

NAND2xp5_ASAP7_75t_L g6765 ( 
.A(n_5670),
.B(n_3397),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_5648),
.Y(n_6766)
);

NAND2xp5_ASAP7_75t_L g6767 ( 
.A(n_5681),
.B(n_3399),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_5784),
.Y(n_6768)
);

INVx1_ASAP7_75t_L g6769 ( 
.A(n_5548),
.Y(n_6769)
);

INVx1_ASAP7_75t_SL g6770 ( 
.A(n_5590),
.Y(n_6770)
);

HB1xp67_ASAP7_75t_L g6771 ( 
.A(n_6119),
.Y(n_6771)
);

AND2x4_ASAP7_75t_L g6772 ( 
.A(n_6072),
.B(n_3518),
.Y(n_6772)
);

AND2x2_ASAP7_75t_L g6773 ( 
.A(n_5845),
.B(n_5570),
.Y(n_6773)
);

AND2x2_ASAP7_75t_L g6774 ( 
.A(n_5928),
.B(n_3400),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_5550),
.Y(n_6775)
);

INVx2_ASAP7_75t_L g6776 ( 
.A(n_5788),
.Y(n_6776)
);

INVx2_ASAP7_75t_L g6777 ( 
.A(n_5794),
.Y(n_6777)
);

INVx1_ASAP7_75t_L g6778 ( 
.A(n_5560),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_5457),
.Y(n_6779)
);

INVx1_ASAP7_75t_L g6780 ( 
.A(n_5666),
.Y(n_6780)
);

BUFx2_ASAP7_75t_L g6781 ( 
.A(n_5990),
.Y(n_6781)
);

INVx1_ASAP7_75t_L g6782 ( 
.A(n_5694),
.Y(n_6782)
);

INVx2_ASAP7_75t_L g6783 ( 
.A(n_5797),
.Y(n_6783)
);

AND2x4_ASAP7_75t_L g6784 ( 
.A(n_6025),
.B(n_3521),
.Y(n_6784)
);

AND2x4_ASAP7_75t_L g6785 ( 
.A(n_6028),
.B(n_3530),
.Y(n_6785)
);

NAND2xp5_ASAP7_75t_L g6786 ( 
.A(n_5711),
.B(n_3401),
.Y(n_6786)
);

INVx1_ASAP7_75t_L g6787 ( 
.A(n_5703),
.Y(n_6787)
);

INVx2_ASAP7_75t_L g6788 ( 
.A(n_5802),
.Y(n_6788)
);

NAND2xp5_ASAP7_75t_L g6789 ( 
.A(n_5559),
.B(n_3405),
.Y(n_6789)
);

XOR2xp5_ASAP7_75t_L g6790 ( 
.A(n_5895),
.B(n_3408),
.Y(n_6790)
);

INVx2_ASAP7_75t_L g6791 ( 
.A(n_5810),
.Y(n_6791)
);

AND2x4_ASAP7_75t_L g6792 ( 
.A(n_6029),
.B(n_3544),
.Y(n_6792)
);

INVx3_ASAP7_75t_L g6793 ( 
.A(n_5574),
.Y(n_6793)
);

INVx1_ASAP7_75t_L g6794 ( 
.A(n_5716),
.Y(n_6794)
);

INVx1_ASAP7_75t_L g6795 ( 
.A(n_5718),
.Y(n_6795)
);

NOR2xp33_ASAP7_75t_L g6796 ( 
.A(n_5876),
.B(n_3409),
.Y(n_6796)
);

INVx2_ASAP7_75t_L g6797 ( 
.A(n_5818),
.Y(n_6797)
);

BUFx8_ASAP7_75t_L g6798 ( 
.A(n_5515),
.Y(n_6798)
);

INVx1_ASAP7_75t_L g6799 ( 
.A(n_5740),
.Y(n_6799)
);

INVx1_ASAP7_75t_L g6800 ( 
.A(n_5765),
.Y(n_6800)
);

BUFx2_ASAP7_75t_L g6801 ( 
.A(n_6103),
.Y(n_6801)
);

NAND2xp5_ASAP7_75t_L g6802 ( 
.A(n_5677),
.B(n_5819),
.Y(n_6802)
);

INVx1_ASAP7_75t_L g6803 ( 
.A(n_5431),
.Y(n_6803)
);

INVx1_ASAP7_75t_L g6804 ( 
.A(n_5455),
.Y(n_6804)
);

INVx1_ASAP7_75t_L g6805 ( 
.A(n_5469),
.Y(n_6805)
);

HB1xp67_ASAP7_75t_L g6806 ( 
.A(n_6065),
.Y(n_6806)
);

HB1xp67_ASAP7_75t_L g6807 ( 
.A(n_5933),
.Y(n_6807)
);

INVx1_ASAP7_75t_SL g6808 ( 
.A(n_6097),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_5482),
.Y(n_6809)
);

BUFx2_ASAP7_75t_L g6810 ( 
.A(n_6040),
.Y(n_6810)
);

INVxp67_ASAP7_75t_L g6811 ( 
.A(n_5527),
.Y(n_6811)
);

INVx1_ASAP7_75t_L g6812 ( 
.A(n_5572),
.Y(n_6812)
);

INVx2_ASAP7_75t_L g6813 ( 
.A(n_5821),
.Y(n_6813)
);

BUFx6f_ASAP7_75t_L g6814 ( 
.A(n_5593),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_5823),
.Y(n_6815)
);

INVx1_ASAP7_75t_L g6816 ( 
.A(n_5656),
.Y(n_6816)
);

INVx1_ASAP7_75t_L g6817 ( 
.A(n_5691),
.Y(n_6817)
);

INVx1_ASAP7_75t_L g6818 ( 
.A(n_6137),
.Y(n_6818)
);

INVx2_ASAP7_75t_L g6819 ( 
.A(n_5865),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6139),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_6161),
.Y(n_6821)
);

INVx2_ASAP7_75t_L g6822 ( 
.A(n_5879),
.Y(n_6822)
);

HB1xp67_ASAP7_75t_L g6823 ( 
.A(n_6105),
.Y(n_6823)
);

NAND2xp5_ASAP7_75t_L g6824 ( 
.A(n_5883),
.B(n_3412),
.Y(n_6824)
);

NAND2xp5_ASAP7_75t_L g6825 ( 
.A(n_5908),
.B(n_3414),
.Y(n_6825)
);

INVx3_ASAP7_75t_L g6826 ( 
.A(n_5612),
.Y(n_6826)
);

INVx1_ASAP7_75t_L g6827 ( 
.A(n_5984),
.Y(n_6827)
);

HB1xp67_ASAP7_75t_L g6828 ( 
.A(n_6107),
.Y(n_6828)
);

BUFx6f_ASAP7_75t_L g6829 ( 
.A(n_5617),
.Y(n_6829)
);

NAND2xp5_ASAP7_75t_L g6830 ( 
.A(n_5871),
.B(n_3415),
.Y(n_6830)
);

INVx2_ASAP7_75t_L g6831 ( 
.A(n_5900),
.Y(n_6831)
);

NAND2xp5_ASAP7_75t_L g6832 ( 
.A(n_5458),
.B(n_3416),
.Y(n_6832)
);

INVx1_ASAP7_75t_L g6833 ( 
.A(n_5629),
.Y(n_6833)
);

INVx2_ASAP7_75t_L g6834 ( 
.A(n_5906),
.Y(n_6834)
);

NAND2xp33_ASAP7_75t_L g6835 ( 
.A(n_6069),
.B(n_3418),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_5912),
.Y(n_6836)
);

CKINVDCx5p33_ASAP7_75t_R g6837 ( 
.A(n_5444),
.Y(n_6837)
);

INVx2_ASAP7_75t_L g6838 ( 
.A(n_5941),
.Y(n_6838)
);

BUFx3_ASAP7_75t_L g6839 ( 
.A(n_5489),
.Y(n_6839)
);

INVx1_ASAP7_75t_L g6840 ( 
.A(n_5630),
.Y(n_6840)
);

INVx1_ASAP7_75t_L g6841 ( 
.A(n_5636),
.Y(n_6841)
);

INVx3_ASAP7_75t_L g6842 ( 
.A(n_5640),
.Y(n_6842)
);

BUFx6f_ASAP7_75t_L g6843 ( 
.A(n_5650),
.Y(n_6843)
);

INVxp67_ASAP7_75t_L g6844 ( 
.A(n_5527),
.Y(n_6844)
);

INVx2_ASAP7_75t_L g6845 ( 
.A(n_5970),
.Y(n_6845)
);

INVx1_ASAP7_75t_L g6846 ( 
.A(n_5655),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_5658),
.Y(n_6847)
);

INVx3_ASAP7_75t_L g6848 ( 
.A(n_5659),
.Y(n_6848)
);

INVx2_ASAP7_75t_L g6849 ( 
.A(n_5960),
.Y(n_6849)
);

INVxp67_ASAP7_75t_L g6850 ( 
.A(n_5847),
.Y(n_6850)
);

HB1xp67_ASAP7_75t_L g6851 ( 
.A(n_6108),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_5442),
.Y(n_6852)
);

INVx2_ASAP7_75t_L g6853 ( 
.A(n_5524),
.Y(n_6853)
);

INVx3_ASAP7_75t_L g6854 ( 
.A(n_6077),
.Y(n_6854)
);

INVx1_ASAP7_75t_L g6855 ( 
.A(n_6109),
.Y(n_6855)
);

BUFx6f_ASAP7_75t_L g6856 ( 
.A(n_5577),
.Y(n_6856)
);

NAND2xp5_ASAP7_75t_L g6857 ( 
.A(n_6098),
.B(n_3421),
.Y(n_6857)
);

CKINVDCx20_ASAP7_75t_R g6858 ( 
.A(n_5731),
.Y(n_6858)
);

INVx3_ASAP7_75t_L g6859 ( 
.A(n_6088),
.Y(n_6859)
);

INVx1_ASAP7_75t_L g6860 ( 
.A(n_5936),
.Y(n_6860)
);

INVx1_ASAP7_75t_L g6861 ( 
.A(n_5937),
.Y(n_6861)
);

INVx1_ASAP7_75t_L g6862 ( 
.A(n_5967),
.Y(n_6862)
);

AND2x2_ASAP7_75t_L g6863 ( 
.A(n_6113),
.B(n_5779),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_5993),
.Y(n_6864)
);

NAND2xp5_ASAP7_75t_L g6865 ( 
.A(n_6006),
.B(n_3424),
.Y(n_6865)
);

NAND2xp5_ASAP7_75t_L g6866 ( 
.A(n_5689),
.B(n_3425),
.Y(n_6866)
);

NOR2xp33_ASAP7_75t_L g6867 ( 
.A(n_6050),
.B(n_3431),
.Y(n_6867)
);

HB1xp67_ASAP7_75t_L g6868 ( 
.A(n_6110),
.Y(n_6868)
);

INVx1_ASAP7_75t_L g6869 ( 
.A(n_6052),
.Y(n_6869)
);

INVx2_ASAP7_75t_L g6870 ( 
.A(n_5606),
.Y(n_6870)
);

INVx2_ASAP7_75t_L g6871 ( 
.A(n_6056),
.Y(n_6871)
);

INVx1_ASAP7_75t_L g6872 ( 
.A(n_6058),
.Y(n_6872)
);

INVx3_ASAP7_75t_L g6873 ( 
.A(n_6089),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6060),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_5449),
.Y(n_6875)
);

INVx1_ASAP7_75t_L g6876 ( 
.A(n_5488),
.Y(n_6876)
);

OA21x2_ASAP7_75t_L g6877 ( 
.A1(n_5476),
.A2(n_5699),
.B(n_5547),
.Y(n_6877)
);

INVx1_ASAP7_75t_L g6878 ( 
.A(n_5847),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_5493),
.Y(n_6879)
);

INVx1_ASAP7_75t_L g6880 ( 
.A(n_5742),
.Y(n_6880)
);

INVx2_ASAP7_75t_L g6881 ( 
.A(n_5938),
.Y(n_6881)
);

BUFx6f_ASAP7_75t_L g6882 ( 
.A(n_6165),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_5824),
.Y(n_6883)
);

HB1xp67_ASAP7_75t_L g6884 ( 
.A(n_6116),
.Y(n_6884)
);

INVx1_ASAP7_75t_L g6885 ( 
.A(n_5956),
.Y(n_6885)
);

AND2x4_ASAP7_75t_L g6886 ( 
.A(n_5724),
.B(n_3550),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6010),
.Y(n_6887)
);

NAND2xp5_ASAP7_75t_SL g6888 ( 
.A(n_5510),
.B(n_3433),
.Y(n_6888)
);

OAI21x1_ASAP7_75t_L g6889 ( 
.A1(n_6062),
.A2(n_3507),
.B(n_3427),
.Y(n_6889)
);

BUFx3_ASAP7_75t_L g6890 ( 
.A(n_5778),
.Y(n_6890)
);

INVx3_ASAP7_75t_L g6891 ( 
.A(n_6053),
.Y(n_6891)
);

HB1xp67_ASAP7_75t_L g6892 ( 
.A(n_6117),
.Y(n_6892)
);

NAND2xp5_ASAP7_75t_SL g6893 ( 
.A(n_6066),
.B(n_3435),
.Y(n_6893)
);

NAND2xp5_ASAP7_75t_L g6894 ( 
.A(n_5586),
.B(n_3437),
.Y(n_6894)
);

INVx1_ASAP7_75t_L g6895 ( 
.A(n_5507),
.Y(n_6895)
);

NAND2xp5_ASAP7_75t_L g6896 ( 
.A(n_5597),
.B(n_3439),
.Y(n_6896)
);

AND2x4_ASAP7_75t_L g6897 ( 
.A(n_5736),
.B(n_3551),
.Y(n_6897)
);

INVx2_ASAP7_75t_L g6898 ( 
.A(n_6074),
.Y(n_6898)
);

INVx6_ASAP7_75t_L g6899 ( 
.A(n_5975),
.Y(n_6899)
);

BUFx6f_ASAP7_75t_L g6900 ( 
.A(n_6181),
.Y(n_6900)
);

NAND2xp33_ASAP7_75t_L g6901 ( 
.A(n_6068),
.B(n_3443),
.Y(n_6901)
);

INVx2_ASAP7_75t_L g6902 ( 
.A(n_6076),
.Y(n_6902)
);

HB1xp67_ASAP7_75t_L g6903 ( 
.A(n_6104),
.Y(n_6903)
);

INVx2_ASAP7_75t_L g6904 ( 
.A(n_6079),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6081),
.Y(n_6905)
);

AND2x2_ASAP7_75t_L g6906 ( 
.A(n_5892),
.B(n_3445),
.Y(n_6906)
);

INVx2_ASAP7_75t_L g6907 ( 
.A(n_6082),
.Y(n_6907)
);

OA21x2_ASAP7_75t_L g6908 ( 
.A1(n_5860),
.A2(n_3573),
.B(n_3554),
.Y(n_6908)
);

INVx2_ASAP7_75t_L g6909 ( 
.A(n_6083),
.Y(n_6909)
);

AND2x4_ASAP7_75t_L g6910 ( 
.A(n_5750),
.B(n_3575),
.Y(n_6910)
);

NOR2xp33_ASAP7_75t_L g6911 ( 
.A(n_6085),
.B(n_3446),
.Y(n_6911)
);

INVx1_ASAP7_75t_L g6912 ( 
.A(n_5546),
.Y(n_6912)
);

NOR2xp33_ASAP7_75t_SL g6913 ( 
.A(n_6124),
.B(n_3447),
.Y(n_6913)
);

BUFx6f_ASAP7_75t_L g6914 ( 
.A(n_6068),
.Y(n_6914)
);

AND2x2_ASAP7_75t_L g6915 ( 
.A(n_5528),
.B(n_3451),
.Y(n_6915)
);

BUFx6f_ASAP7_75t_L g6916 ( 
.A(n_6053),
.Y(n_6916)
);

INVx1_ASAP7_75t_L g6917 ( 
.A(n_5638),
.Y(n_6917)
);

NAND2xp5_ASAP7_75t_L g6918 ( 
.A(n_5643),
.B(n_3452),
.Y(n_6918)
);

INVx1_ASAP7_75t_L g6919 ( 
.A(n_5673),
.Y(n_6919)
);

INVx3_ASAP7_75t_L g6920 ( 
.A(n_6099),
.Y(n_6920)
);

INVx1_ASAP7_75t_L g6921 ( 
.A(n_5695),
.Y(n_6921)
);

INVxp67_ASAP7_75t_L g6922 ( 
.A(n_6118),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_5697),
.Y(n_6923)
);

AND2x4_ASAP7_75t_L g6924 ( 
.A(n_6102),
.B(n_3576),
.Y(n_6924)
);

INVx2_ASAP7_75t_L g6925 ( 
.A(n_5434),
.Y(n_6925)
);

INVx1_ASAP7_75t_L g6926 ( 
.A(n_5775),
.Y(n_6926)
);

INVx1_ASAP7_75t_L g6927 ( 
.A(n_5959),
.Y(n_6927)
);

INVx1_ASAP7_75t_L g6928 ( 
.A(n_6023),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_6080),
.Y(n_6929)
);

INVxp67_ASAP7_75t_L g6930 ( 
.A(n_6091),
.Y(n_6930)
);

BUFx6f_ASAP7_75t_L g6931 ( 
.A(n_6172),
.Y(n_6931)
);

OA21x2_ASAP7_75t_L g6932 ( 
.A1(n_6114),
.A2(n_3578),
.B(n_3577),
.Y(n_6932)
);

NAND2xp5_ASAP7_75t_L g6933 ( 
.A(n_5904),
.B(n_5992),
.Y(n_6933)
);

INVxp67_ASAP7_75t_L g6934 ( 
.A(n_6032),
.Y(n_6934)
);

BUFx6f_ASAP7_75t_L g6935 ( 
.A(n_6188),
.Y(n_6935)
);

BUFx2_ASAP7_75t_L g6936 ( 
.A(n_5501),
.Y(n_6936)
);

NAND2xp5_ASAP7_75t_L g6937 ( 
.A(n_6051),
.B(n_3453),
.Y(n_6937)
);

BUFx6f_ASAP7_75t_L g6938 ( 
.A(n_5922),
.Y(n_6938)
);

INVx2_ASAP7_75t_L g6939 ( 
.A(n_5946),
.Y(n_6939)
);

AND2x2_ASAP7_75t_L g6940 ( 
.A(n_5803),
.B(n_3455),
.Y(n_6940)
);

INVx1_ASAP7_75t_L g6941 ( 
.A(n_5995),
.Y(n_6941)
);

NAND2xp5_ASAP7_75t_L g6942 ( 
.A(n_5877),
.B(n_3457),
.Y(n_6942)
);

AND3x1_ASAP7_75t_L g6943 ( 
.A(n_5762),
.B(n_3582),
.C(n_3579),
.Y(n_6943)
);

INVx1_ASAP7_75t_L g6944 ( 
.A(n_5885),
.Y(n_6944)
);

INVx2_ASAP7_75t_L g6945 ( 
.A(n_5627),
.Y(n_6945)
);

NAND2xp5_ASAP7_75t_SL g6946 ( 
.A(n_6151),
.B(n_3458),
.Y(n_6946)
);

INVx2_ASAP7_75t_L g6947 ( 
.A(n_5627),
.Y(n_6947)
);

BUFx6f_ASAP7_75t_L g6948 ( 
.A(n_5438),
.Y(n_6948)
);

INVxp67_ASAP7_75t_L g6949 ( 
.A(n_5426),
.Y(n_6949)
);

INVx3_ASAP7_75t_L g6950 ( 
.A(n_5979),
.Y(n_6950)
);

NAND2xp5_ASAP7_75t_L g6951 ( 
.A(n_6186),
.B(n_3461),
.Y(n_6951)
);

INVx2_ASAP7_75t_L g6952 ( 
.A(n_6196),
.Y(n_6952)
);

NAND2xp5_ASAP7_75t_SL g6953 ( 
.A(n_6261),
.B(n_3463),
.Y(n_6953)
);

AOI22xp33_ASAP7_75t_L g6954 ( 
.A1(n_6939),
.A2(n_3466),
.B1(n_3470),
.B2(n_3469),
.Y(n_6954)
);

INVx2_ASAP7_75t_L g6955 ( 
.A(n_6945),
.Y(n_6955)
);

BUFx3_ASAP7_75t_L g6956 ( 
.A(n_6659),
.Y(n_6956)
);

INVx2_ASAP7_75t_L g6957 ( 
.A(n_6947),
.Y(n_6957)
);

BUFx3_ASAP7_75t_L g6958 ( 
.A(n_6203),
.Y(n_6958)
);

NAND2xp5_ASAP7_75t_SL g6959 ( 
.A(n_6927),
.B(n_3472),
.Y(n_6959)
);

INVx2_ASAP7_75t_L g6960 ( 
.A(n_6202),
.Y(n_6960)
);

INVxp67_ASAP7_75t_SL g6961 ( 
.A(n_6807),
.Y(n_6961)
);

INVx2_ASAP7_75t_L g6962 ( 
.A(n_6205),
.Y(n_6962)
);

NAND2xp5_ASAP7_75t_SL g6963 ( 
.A(n_6928),
.B(n_3473),
.Y(n_6963)
);

INVx1_ASAP7_75t_L g6964 ( 
.A(n_6200),
.Y(n_6964)
);

BUFx6f_ASAP7_75t_L g6965 ( 
.A(n_6257),
.Y(n_6965)
);

NOR2xp33_ASAP7_75t_L g6966 ( 
.A(n_6341),
.B(n_3474),
.Y(n_6966)
);

INVx4_ASAP7_75t_L g6967 ( 
.A(n_6624),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6333),
.B(n_3476),
.Y(n_6968)
);

BUFx3_ASAP7_75t_L g6969 ( 
.A(n_6211),
.Y(n_6969)
);

AOI22xp33_ASAP7_75t_L g6970 ( 
.A1(n_6233),
.A2(n_6432),
.B1(n_6929),
.B2(n_6876),
.Y(n_6970)
);

INVx2_ASAP7_75t_L g6971 ( 
.A(n_6206),
.Y(n_6971)
);

NAND2xp5_ASAP7_75t_SL g6972 ( 
.A(n_6934),
.B(n_3477),
.Y(n_6972)
);

AND2x2_ASAP7_75t_L g6973 ( 
.A(n_6253),
.B(n_3478),
.Y(n_6973)
);

NAND2xp5_ASAP7_75t_SL g6974 ( 
.A(n_6879),
.B(n_3482),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6204),
.Y(n_6975)
);

NAND2xp5_ASAP7_75t_SL g6976 ( 
.A(n_6880),
.B(n_3483),
.Y(n_6976)
);

INVx1_ASAP7_75t_L g6977 ( 
.A(n_6209),
.Y(n_6977)
);

INVx2_ASAP7_75t_L g6978 ( 
.A(n_6214),
.Y(n_6978)
);

INVx2_ASAP7_75t_L g6979 ( 
.A(n_6220),
.Y(n_6979)
);

INVx2_ASAP7_75t_L g6980 ( 
.A(n_6225),
.Y(n_6980)
);

AND2x2_ASAP7_75t_L g6981 ( 
.A(n_6201),
.B(n_3487),
.Y(n_6981)
);

INVx2_ASAP7_75t_L g6982 ( 
.A(n_6237),
.Y(n_6982)
);

INVx4_ASAP7_75t_L g6983 ( 
.A(n_6624),
.Y(n_6983)
);

INVx1_ASAP7_75t_L g6984 ( 
.A(n_6217),
.Y(n_6984)
);

INVx6_ASAP7_75t_L g6985 ( 
.A(n_6246),
.Y(n_6985)
);

INVx4_ASAP7_75t_L g6986 ( 
.A(n_6545),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6223),
.Y(n_6987)
);

INVx2_ASAP7_75t_L g6988 ( 
.A(n_6238),
.Y(n_6988)
);

OR2x6_ASAP7_75t_L g6989 ( 
.A(n_6899),
.B(n_6365),
.Y(n_6989)
);

BUFx6f_ASAP7_75t_L g6990 ( 
.A(n_6257),
.Y(n_6990)
);

NAND2xp5_ASAP7_75t_SL g6991 ( 
.A(n_6883),
.B(n_3488),
.Y(n_6991)
);

INVx3_ASAP7_75t_L g6992 ( 
.A(n_6469),
.Y(n_6992)
);

INVx1_ASAP7_75t_L g6993 ( 
.A(n_6230),
.Y(n_6993)
);

NAND2xp5_ASAP7_75t_L g6994 ( 
.A(n_6691),
.B(n_3491),
.Y(n_6994)
);

INVx2_ASAP7_75t_L g6995 ( 
.A(n_6242),
.Y(n_6995)
);

INVx5_ASAP7_75t_L g6996 ( 
.A(n_6702),
.Y(n_6996)
);

INVx2_ASAP7_75t_L g6997 ( 
.A(n_6243),
.Y(n_6997)
);

AOI22xp5_ASAP7_75t_L g6998 ( 
.A1(n_6424),
.A2(n_3492),
.B1(n_3494),
.B2(n_3493),
.Y(n_6998)
);

OAI22xp33_ASAP7_75t_L g6999 ( 
.A1(n_6933),
.A2(n_3496),
.B1(n_3504),
.B2(n_3502),
.Y(n_6999)
);

NAND2xp5_ASAP7_75t_SL g7000 ( 
.A(n_6885),
.B(n_3505),
.Y(n_7000)
);

BUFx6f_ASAP7_75t_L g7001 ( 
.A(n_6545),
.Y(n_7001)
);

INVx2_ASAP7_75t_L g7002 ( 
.A(n_6245),
.Y(n_7002)
);

NAND2xp5_ASAP7_75t_SL g7003 ( 
.A(n_6887),
.B(n_3506),
.Y(n_7003)
);

NOR2xp33_ASAP7_75t_L g7004 ( 
.A(n_6467),
.B(n_3508),
.Y(n_7004)
);

BUFx6f_ASAP7_75t_L g7005 ( 
.A(n_6548),
.Y(n_7005)
);

INVx2_ASAP7_75t_SL g7006 ( 
.A(n_6329),
.Y(n_7006)
);

OR2x2_ASAP7_75t_L g7007 ( 
.A(n_6306),
.B(n_3509),
.Y(n_7007)
);

INVx1_ASAP7_75t_L g7008 ( 
.A(n_6241),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_6258),
.Y(n_7009)
);

INVx3_ASAP7_75t_L g7010 ( 
.A(n_6548),
.Y(n_7010)
);

INVx1_ASAP7_75t_SL g7011 ( 
.A(n_6354),
.Y(n_7011)
);

NAND3x1_ASAP7_75t_L g7012 ( 
.A(n_6940),
.B(n_2641),
.C(n_2563),
.Y(n_7012)
);

INVx2_ASAP7_75t_L g7013 ( 
.A(n_6247),
.Y(n_7013)
);

INVx1_ASAP7_75t_L g7014 ( 
.A(n_6265),
.Y(n_7014)
);

BUFx3_ASAP7_75t_L g7015 ( 
.A(n_6276),
.Y(n_7015)
);

BUFx4f_ASAP7_75t_L g7016 ( 
.A(n_6702),
.Y(n_7016)
);

INVx2_ASAP7_75t_SL g7017 ( 
.A(n_6282),
.Y(n_7017)
);

INVx1_ASAP7_75t_SL g7018 ( 
.A(n_6472),
.Y(n_7018)
);

AND2x6_ASAP7_75t_L g7019 ( 
.A(n_6914),
.B(n_3601),
.Y(n_7019)
);

INVx2_ASAP7_75t_L g7020 ( 
.A(n_6248),
.Y(n_7020)
);

NOR2xp33_ASAP7_75t_SL g7021 ( 
.A(n_6252),
.B(n_3510),
.Y(n_7021)
);

NAND2xp5_ASAP7_75t_SL g7022 ( 
.A(n_6546),
.B(n_3511),
.Y(n_7022)
);

INVx5_ASAP7_75t_L g7023 ( 
.A(n_6390),
.Y(n_7023)
);

BUFx6f_ASAP7_75t_L g7024 ( 
.A(n_6552),
.Y(n_7024)
);

INVxp33_ASAP7_75t_SL g7025 ( 
.A(n_6286),
.Y(n_7025)
);

INVx2_ASAP7_75t_L g7026 ( 
.A(n_6250),
.Y(n_7026)
);

NAND2xp5_ASAP7_75t_SL g7027 ( 
.A(n_6495),
.B(n_3512),
.Y(n_7027)
);

AND2x2_ASAP7_75t_L g7028 ( 
.A(n_6774),
.B(n_3513),
.Y(n_7028)
);

INVx2_ASAP7_75t_L g7029 ( 
.A(n_6254),
.Y(n_7029)
);

INVx4_ASAP7_75t_L g7030 ( 
.A(n_6552),
.Y(n_7030)
);

INVx3_ASAP7_75t_L g7031 ( 
.A(n_6583),
.Y(n_7031)
);

INVx2_ASAP7_75t_L g7032 ( 
.A(n_6263),
.Y(n_7032)
);

NOR2xp33_ASAP7_75t_L g7033 ( 
.A(n_6949),
.B(n_3519),
.Y(n_7033)
);

NAND2xp5_ASAP7_75t_L g7034 ( 
.A(n_6605),
.B(n_3523),
.Y(n_7034)
);

AOI22xp33_ASAP7_75t_L g7035 ( 
.A1(n_6875),
.A2(n_6903),
.B1(n_6509),
.B2(n_6362),
.Y(n_7035)
);

INVx2_ASAP7_75t_L g7036 ( 
.A(n_6264),
.Y(n_7036)
);

INVx3_ASAP7_75t_L g7037 ( 
.A(n_6583),
.Y(n_7037)
);

INVx2_ASAP7_75t_L g7038 ( 
.A(n_6275),
.Y(n_7038)
);

NOR2xp33_ASAP7_75t_L g7039 ( 
.A(n_6692),
.B(n_3524),
.Y(n_7039)
);

NOR2xp33_ASAP7_75t_L g7040 ( 
.A(n_6409),
.B(n_3525),
.Y(n_7040)
);

INVx2_ASAP7_75t_L g7041 ( 
.A(n_6278),
.Y(n_7041)
);

INVx2_ASAP7_75t_L g7042 ( 
.A(n_6279),
.Y(n_7042)
);

NOR2xp33_ASAP7_75t_L g7043 ( 
.A(n_6470),
.B(n_3528),
.Y(n_7043)
);

INVx3_ASAP7_75t_L g7044 ( 
.A(n_6598),
.Y(n_7044)
);

BUFx3_ASAP7_75t_L g7045 ( 
.A(n_6598),
.Y(n_7045)
);

OR2x6_ASAP7_75t_L g7046 ( 
.A(n_6606),
.B(n_3515),
.Y(n_7046)
);

INVx2_ASAP7_75t_L g7047 ( 
.A(n_6280),
.Y(n_7047)
);

INVx1_ASAP7_75t_L g7048 ( 
.A(n_6267),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_6268),
.Y(n_7049)
);

AND2x2_ASAP7_75t_SL g7050 ( 
.A(n_6935),
.B(n_3532),
.Y(n_7050)
);

AND3x2_ASAP7_75t_L g7051 ( 
.A(n_6357),
.B(n_3607),
.C(n_3588),
.Y(n_7051)
);

INVx1_ASAP7_75t_L g7052 ( 
.A(n_6270),
.Y(n_7052)
);

NOR2xp33_ASAP7_75t_L g7053 ( 
.A(n_6936),
.B(n_3529),
.Y(n_7053)
);

INVx1_ASAP7_75t_L g7054 ( 
.A(n_6277),
.Y(n_7054)
);

INVx1_ASAP7_75t_L g7055 ( 
.A(n_6281),
.Y(n_7055)
);

NAND2xp5_ASAP7_75t_SL g7056 ( 
.A(n_6920),
.B(n_3531),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_6285),
.Y(n_7057)
);

INVx1_ASAP7_75t_L g7058 ( 
.A(n_6288),
.Y(n_7058)
);

BUFx2_ASAP7_75t_L g7059 ( 
.A(n_6240),
.Y(n_7059)
);

NAND2xp33_ASAP7_75t_L g7060 ( 
.A(n_6308),
.B(n_3533),
.Y(n_7060)
);

NAND3xp33_ASAP7_75t_L g7061 ( 
.A(n_6651),
.B(n_3535),
.C(n_3534),
.Y(n_7061)
);

INVx2_ASAP7_75t_L g7062 ( 
.A(n_6284),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_SL g7063 ( 
.A(n_6670),
.B(n_3536),
.Y(n_7063)
);

NAND2xp5_ASAP7_75t_SL g7064 ( 
.A(n_6916),
.B(n_3540),
.Y(n_7064)
);

CKINVDCx5p33_ASAP7_75t_R g7065 ( 
.A(n_6737),
.Y(n_7065)
);

INVx2_ASAP7_75t_L g7066 ( 
.A(n_6292),
.Y(n_7066)
);

NAND2xp5_ASAP7_75t_SL g7067 ( 
.A(n_6916),
.B(n_3542),
.Y(n_7067)
);

INVx4_ASAP7_75t_L g7068 ( 
.A(n_6606),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6290),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_6294),
.Y(n_7070)
);

NAND2xp5_ASAP7_75t_SL g7071 ( 
.A(n_6922),
.B(n_3543),
.Y(n_7071)
);

AO21x2_ASAP7_75t_L g7072 ( 
.A1(n_6198),
.A2(n_3603),
.B(n_3602),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6296),
.Y(n_7073)
);

INVx2_ASAP7_75t_SL g7074 ( 
.A(n_6289),
.Y(n_7074)
);

OR2x6_ASAP7_75t_L g7075 ( 
.A(n_6615),
.B(n_3620),
.Y(n_7075)
);

INVx2_ASAP7_75t_L g7076 ( 
.A(n_6305),
.Y(n_7076)
);

NAND2xp5_ASAP7_75t_L g7077 ( 
.A(n_6677),
.B(n_3546),
.Y(n_7077)
);

NAND2xp5_ASAP7_75t_SL g7078 ( 
.A(n_6519),
.B(n_3547),
.Y(n_7078)
);

INVx2_ASAP7_75t_L g7079 ( 
.A(n_6320),
.Y(n_7079)
);

OR2x2_ASAP7_75t_L g7080 ( 
.A(n_6303),
.B(n_3548),
.Y(n_7080)
);

INVx2_ASAP7_75t_L g7081 ( 
.A(n_6417),
.Y(n_7081)
);

INVx2_ASAP7_75t_L g7082 ( 
.A(n_6421),
.Y(n_7082)
);

INVx2_ASAP7_75t_L g7083 ( 
.A(n_6426),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_6297),
.Y(n_7084)
);

NAND2xp5_ASAP7_75t_L g7085 ( 
.A(n_6609),
.B(n_3552),
.Y(n_7085)
);

INVx3_ASAP7_75t_L g7086 ( 
.A(n_6615),
.Y(n_7086)
);

OR2x6_ASAP7_75t_L g7087 ( 
.A(n_6623),
.B(n_3646),
.Y(n_7087)
);

INVx1_ASAP7_75t_L g7088 ( 
.A(n_6298),
.Y(n_7088)
);

INVx1_ASAP7_75t_SL g7089 ( 
.A(n_6571),
.Y(n_7089)
);

BUFx6f_ASAP7_75t_L g7090 ( 
.A(n_6623),
.Y(n_7090)
);

INVx2_ASAP7_75t_L g7091 ( 
.A(n_6433),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_6301),
.Y(n_7092)
);

INVx2_ASAP7_75t_L g7093 ( 
.A(n_6436),
.Y(n_7093)
);

INVx1_ASAP7_75t_L g7094 ( 
.A(n_6307),
.Y(n_7094)
);

INVx1_ASAP7_75t_L g7095 ( 
.A(n_6310),
.Y(n_7095)
);

INVx2_ASAP7_75t_SL g7096 ( 
.A(n_6425),
.Y(n_7096)
);

NAND2xp5_ASAP7_75t_SL g7097 ( 
.A(n_6898),
.B(n_3553),
.Y(n_7097)
);

INVx1_ASAP7_75t_L g7098 ( 
.A(n_6312),
.Y(n_7098)
);

INVx3_ASAP7_75t_L g7099 ( 
.A(n_6628),
.Y(n_7099)
);

INVx1_ASAP7_75t_L g7100 ( 
.A(n_6315),
.Y(n_7100)
);

OR2x6_ASAP7_75t_L g7101 ( 
.A(n_6628),
.B(n_3670),
.Y(n_7101)
);

OR2x6_ASAP7_75t_L g7102 ( 
.A(n_6631),
.B(n_3703),
.Y(n_7102)
);

INVx2_ASAP7_75t_L g7103 ( 
.A(n_6437),
.Y(n_7103)
);

OR2x6_ASAP7_75t_L g7104 ( 
.A(n_6631),
.B(n_3751),
.Y(n_7104)
);

INVx2_ASAP7_75t_L g7105 ( 
.A(n_6438),
.Y(n_7105)
);

INVx2_ASAP7_75t_SL g7106 ( 
.A(n_6359),
.Y(n_7106)
);

AO21x2_ASAP7_75t_L g7107 ( 
.A1(n_6803),
.A2(n_3627),
.B(n_3624),
.Y(n_7107)
);

AND2x2_ASAP7_75t_L g7108 ( 
.A(n_6773),
.B(n_3556),
.Y(n_7108)
);

NAND2xp5_ASAP7_75t_L g7109 ( 
.A(n_6610),
.B(n_3559),
.Y(n_7109)
);

INVx2_ASAP7_75t_L g7110 ( 
.A(n_6445),
.Y(n_7110)
);

XNOR2xp5_ASAP7_75t_L g7111 ( 
.A(n_6249),
.B(n_3560),
.Y(n_7111)
);

NOR2xp33_ASAP7_75t_L g7112 ( 
.A(n_6534),
.B(n_3561),
.Y(n_7112)
);

INVx1_ASAP7_75t_L g7113 ( 
.A(n_6317),
.Y(n_7113)
);

INVx8_ASAP7_75t_L g7114 ( 
.A(n_6295),
.Y(n_7114)
);

AOI22xp33_ASAP7_75t_L g7115 ( 
.A1(n_6362),
.A2(n_3563),
.B1(n_3566),
.B2(n_3564),
.Y(n_7115)
);

INVx2_ASAP7_75t_L g7116 ( 
.A(n_6446),
.Y(n_7116)
);

OR2x2_ASAP7_75t_L g7117 ( 
.A(n_6309),
.B(n_3569),
.Y(n_7117)
);

INVx4_ASAP7_75t_SL g7118 ( 
.A(n_6931),
.Y(n_7118)
);

INVx1_ASAP7_75t_L g7119 ( 
.A(n_6318),
.Y(n_7119)
);

AOI22xp33_ASAP7_75t_SL g7120 ( 
.A1(n_6266),
.A2(n_3571),
.B1(n_3572),
.B2(n_3570),
.Y(n_7120)
);

AND2x4_ASAP7_75t_L g7121 ( 
.A(n_6366),
.B(n_3630),
.Y(n_7121)
);

INVx2_ASAP7_75t_SL g7122 ( 
.A(n_6375),
.Y(n_7122)
);

INVx2_ASAP7_75t_L g7123 ( 
.A(n_6448),
.Y(n_7123)
);

INVx1_ASAP7_75t_L g7124 ( 
.A(n_6321),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_6325),
.Y(n_7125)
);

INVx1_ASAP7_75t_L g7126 ( 
.A(n_6327),
.Y(n_7126)
);

AO22x2_ASAP7_75t_L g7127 ( 
.A1(n_6274),
.A2(n_3635),
.B1(n_3637),
.B2(n_3632),
.Y(n_7127)
);

INVx1_ASAP7_75t_L g7128 ( 
.A(n_6328),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_6338),
.Y(n_7129)
);

INVx4_ASAP7_75t_L g7130 ( 
.A(n_6645),
.Y(n_7130)
);

BUFx6f_ASAP7_75t_SL g7131 ( 
.A(n_6839),
.Y(n_7131)
);

INVx2_ASAP7_75t_L g7132 ( 
.A(n_6454),
.Y(n_7132)
);

XNOR2xp5_ASAP7_75t_L g7133 ( 
.A(n_6790),
.B(n_3574),
.Y(n_7133)
);

BUFx6f_ASAP7_75t_L g7134 ( 
.A(n_6645),
.Y(n_7134)
);

INVx1_ASAP7_75t_SL g7135 ( 
.A(n_6573),
.Y(n_7135)
);

NAND2xp5_ASAP7_75t_SL g7136 ( 
.A(n_6902),
.B(n_3581),
.Y(n_7136)
);

AND2x2_ASAP7_75t_SL g7137 ( 
.A(n_6935),
.B(n_6474),
.Y(n_7137)
);

NOR2xp33_ASAP7_75t_L g7138 ( 
.A(n_6228),
.B(n_6666),
.Y(n_7138)
);

NOR2xp33_ASAP7_75t_L g7139 ( 
.A(n_6761),
.B(n_3583),
.Y(n_7139)
);

INVx4_ASAP7_75t_L g7140 ( 
.A(n_6664),
.Y(n_7140)
);

INVx2_ASAP7_75t_L g7141 ( 
.A(n_6461),
.Y(n_7141)
);

INVx2_ASAP7_75t_L g7142 ( 
.A(n_6463),
.Y(n_7142)
);

INVx4_ASAP7_75t_L g7143 ( 
.A(n_6664),
.Y(n_7143)
);

AOI22xp33_ASAP7_75t_L g7144 ( 
.A1(n_6362),
.A2(n_3584),
.B1(n_3587),
.B2(n_3585),
.Y(n_7144)
);

INVx2_ASAP7_75t_L g7145 ( 
.A(n_6482),
.Y(n_7145)
);

INVx2_ASAP7_75t_L g7146 ( 
.A(n_6484),
.Y(n_7146)
);

INVx3_ASAP7_75t_L g7147 ( 
.A(n_6678),
.Y(n_7147)
);

INVx2_ASAP7_75t_L g7148 ( 
.A(n_6487),
.Y(n_7148)
);

NAND2xp5_ASAP7_75t_SL g7149 ( 
.A(n_6904),
.B(n_3592),
.Y(n_7149)
);

AOI22xp33_ASAP7_75t_L g7150 ( 
.A1(n_6509),
.A2(n_3593),
.B1(n_3604),
.B2(n_3594),
.Y(n_7150)
);

INVx2_ASAP7_75t_L g7151 ( 
.A(n_6500),
.Y(n_7151)
);

INVx2_ASAP7_75t_L g7152 ( 
.A(n_6506),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_6343),
.Y(n_7153)
);

NOR2xp33_ASAP7_75t_L g7154 ( 
.A(n_6334),
.B(n_3605),
.Y(n_7154)
);

OR2x6_ASAP7_75t_L g7155 ( 
.A(n_6678),
.B(n_3789),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_6352),
.Y(n_7156)
);

INVx3_ASAP7_75t_L g7157 ( 
.A(n_6697),
.Y(n_7157)
);

CKINVDCx5p33_ASAP7_75t_R g7158 ( 
.A(n_6376),
.Y(n_7158)
);

INVx2_ASAP7_75t_L g7159 ( 
.A(n_6507),
.Y(n_7159)
);

NAND2xp5_ASAP7_75t_SL g7160 ( 
.A(n_6907),
.B(n_3606),
.Y(n_7160)
);

INVx2_ASAP7_75t_L g7161 ( 
.A(n_6518),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_6355),
.Y(n_7162)
);

INVx1_ASAP7_75t_L g7163 ( 
.A(n_6356),
.Y(n_7163)
);

AO21x2_ASAP7_75t_L g7164 ( 
.A1(n_6804),
.A2(n_3640),
.B(n_3639),
.Y(n_7164)
);

AOI22xp5_ASAP7_75t_L g7165 ( 
.A1(n_6509),
.A2(n_3609),
.B1(n_3611),
.B2(n_3610),
.Y(n_7165)
);

INVx1_ASAP7_75t_L g7166 ( 
.A(n_6367),
.Y(n_7166)
);

INVx3_ASAP7_75t_L g7167 ( 
.A(n_6697),
.Y(n_7167)
);

INVx2_ASAP7_75t_SL g7168 ( 
.A(n_6617),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_6369),
.Y(n_7169)
);

NAND2xp5_ASAP7_75t_L g7170 ( 
.A(n_6657),
.B(n_3612),
.Y(n_7170)
);

INVx2_ASAP7_75t_L g7171 ( 
.A(n_6524),
.Y(n_7171)
);

INVx2_ASAP7_75t_L g7172 ( 
.A(n_6525),
.Y(n_7172)
);

NAND2xp5_ASAP7_75t_SL g7173 ( 
.A(n_6909),
.B(n_6300),
.Y(n_7173)
);

NAND3xp33_ASAP7_75t_L g7174 ( 
.A(n_6302),
.B(n_6796),
.C(n_6704),
.Y(n_7174)
);

INVx2_ASAP7_75t_L g7175 ( 
.A(n_6533),
.Y(n_7175)
);

INVx2_ASAP7_75t_L g7176 ( 
.A(n_6536),
.Y(n_7176)
);

INVx2_ASAP7_75t_L g7177 ( 
.A(n_6543),
.Y(n_7177)
);

NAND2xp5_ASAP7_75t_SL g7178 ( 
.A(n_6721),
.B(n_3614),
.Y(n_7178)
);

INVx1_ASAP7_75t_L g7179 ( 
.A(n_6374),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_6377),
.Y(n_7180)
);

INVx2_ASAP7_75t_L g7181 ( 
.A(n_6549),
.Y(n_7181)
);

NAND2xp5_ASAP7_75t_L g7182 ( 
.A(n_6661),
.B(n_3615),
.Y(n_7182)
);

INVx1_ASAP7_75t_L g7183 ( 
.A(n_6379),
.Y(n_7183)
);

NAND2xp5_ASAP7_75t_SL g7184 ( 
.A(n_6727),
.B(n_3616),
.Y(n_7184)
);

NAND2xp5_ASAP7_75t_L g7185 ( 
.A(n_6663),
.B(n_3619),
.Y(n_7185)
);

NAND2xp5_ASAP7_75t_SL g7186 ( 
.A(n_6802),
.B(n_3622),
.Y(n_7186)
);

INVx2_ASAP7_75t_L g7187 ( 
.A(n_6562),
.Y(n_7187)
);

NAND2xp5_ASAP7_75t_SL g7188 ( 
.A(n_6905),
.B(n_3623),
.Y(n_7188)
);

INVx1_ASAP7_75t_L g7189 ( 
.A(n_6382),
.Y(n_7189)
);

INVx2_ASAP7_75t_SL g7190 ( 
.A(n_6526),
.Y(n_7190)
);

INVx2_ASAP7_75t_L g7191 ( 
.A(n_6570),
.Y(n_7191)
);

INVx1_ASAP7_75t_L g7192 ( 
.A(n_6388),
.Y(n_7192)
);

BUFx3_ASAP7_75t_L g7193 ( 
.A(n_6295),
.Y(n_7193)
);

NAND2xp5_ASAP7_75t_L g7194 ( 
.A(n_6671),
.B(n_3625),
.Y(n_7194)
);

INVx1_ASAP7_75t_L g7195 ( 
.A(n_6392),
.Y(n_7195)
);

INVx2_ASAP7_75t_L g7196 ( 
.A(n_6575),
.Y(n_7196)
);

INVx2_ASAP7_75t_L g7197 ( 
.A(n_6589),
.Y(n_7197)
);

AND2x2_ASAP7_75t_L g7198 ( 
.A(n_6322),
.B(n_3628),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_6393),
.Y(n_7199)
);

INVx2_ASAP7_75t_L g7200 ( 
.A(n_6590),
.Y(n_7200)
);

AOI22xp33_ASAP7_75t_L g7201 ( 
.A1(n_6863),
.A2(n_3629),
.B1(n_3643),
.B2(n_3633),
.Y(n_7201)
);

NAND2xp5_ASAP7_75t_SL g7202 ( 
.A(n_6891),
.B(n_3644),
.Y(n_7202)
);

INVx1_ASAP7_75t_L g7203 ( 
.A(n_6395),
.Y(n_7203)
);

INVx2_ASAP7_75t_L g7204 ( 
.A(n_6596),
.Y(n_7204)
);

INVx3_ASAP7_75t_L g7205 ( 
.A(n_6468),
.Y(n_7205)
);

INVx1_ASAP7_75t_L g7206 ( 
.A(n_6396),
.Y(n_7206)
);

NAND2xp33_ASAP7_75t_SL g7207 ( 
.A(n_6681),
.B(n_3652),
.Y(n_7207)
);

CKINVDCx5p33_ASAP7_75t_R g7208 ( 
.A(n_6380),
.Y(n_7208)
);

CKINVDCx5p33_ASAP7_75t_R g7209 ( 
.A(n_6492),
.Y(n_7209)
);

INVx1_ASAP7_75t_L g7210 ( 
.A(n_6404),
.Y(n_7210)
);

NOR2xp33_ASAP7_75t_L g7211 ( 
.A(n_6262),
.B(n_3653),
.Y(n_7211)
);

INVx1_ASAP7_75t_L g7212 ( 
.A(n_6405),
.Y(n_7212)
);

INVx5_ASAP7_75t_L g7213 ( 
.A(n_6390),
.Y(n_7213)
);

NAND2xp5_ASAP7_75t_SL g7214 ( 
.A(n_6779),
.B(n_3656),
.Y(n_7214)
);

NAND2xp33_ASAP7_75t_L g7215 ( 
.A(n_6611),
.B(n_3657),
.Y(n_7215)
);

NAND2xp5_ASAP7_75t_SL g7216 ( 
.A(n_6912),
.B(n_3658),
.Y(n_7216)
);

AOI22xp33_ASAP7_75t_L g7217 ( 
.A1(n_6895),
.A2(n_3661),
.B1(n_3663),
.B2(n_3660),
.Y(n_7217)
);

HB1xp67_ASAP7_75t_L g7218 ( 
.A(n_6345),
.Y(n_7218)
);

BUFx3_ASAP7_75t_L g7219 ( 
.A(n_6299),
.Y(n_7219)
);

INVx1_ASAP7_75t_L g7220 ( 
.A(n_6406),
.Y(n_7220)
);

NAND2xp5_ASAP7_75t_L g7221 ( 
.A(n_6672),
.B(n_6674),
.Y(n_7221)
);

NAND2xp33_ASAP7_75t_L g7222 ( 
.A(n_6612),
.B(n_3664),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_6407),
.Y(n_7223)
);

NOR2xp33_ASAP7_75t_L g7224 ( 
.A(n_6449),
.B(n_3665),
.Y(n_7224)
);

NAND2xp5_ASAP7_75t_L g7225 ( 
.A(n_6613),
.B(n_6620),
.Y(n_7225)
);

AND2x4_ASAP7_75t_L g7226 ( 
.A(n_6400),
.B(n_6299),
.Y(n_7226)
);

INVx3_ASAP7_75t_L g7227 ( 
.A(n_6451),
.Y(n_7227)
);

NAND2xp5_ASAP7_75t_SL g7228 ( 
.A(n_6917),
.B(n_3668),
.Y(n_7228)
);

INVx4_ASAP7_75t_SL g7229 ( 
.A(n_6931),
.Y(n_7229)
);

INVx2_ASAP7_75t_SL g7230 ( 
.A(n_6271),
.Y(n_7230)
);

INVx1_ASAP7_75t_L g7231 ( 
.A(n_6408),
.Y(n_7231)
);

NAND2xp5_ASAP7_75t_SL g7232 ( 
.A(n_6919),
.B(n_3669),
.Y(n_7232)
);

NAND2xp33_ASAP7_75t_R g7233 ( 
.A(n_6837),
.B(n_3671),
.Y(n_7233)
);

BUFx6f_ASAP7_75t_L g7234 ( 
.A(n_6304),
.Y(n_7234)
);

BUFx6f_ASAP7_75t_L g7235 ( 
.A(n_6304),
.Y(n_7235)
);

INVx2_ASAP7_75t_SL g7236 ( 
.A(n_6293),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_6414),
.Y(n_7237)
);

INVx2_ASAP7_75t_L g7238 ( 
.A(n_6601),
.Y(n_7238)
);

INVx2_ASAP7_75t_L g7239 ( 
.A(n_6608),
.Y(n_7239)
);

INVx1_ASAP7_75t_L g7240 ( 
.A(n_6416),
.Y(n_7240)
);

NOR2xp33_ASAP7_75t_L g7241 ( 
.A(n_6930),
.B(n_3672),
.Y(n_7241)
);

NOR2xp33_ASAP7_75t_L g7242 ( 
.A(n_6733),
.B(n_3673),
.Y(n_7242)
);

INVx1_ASAP7_75t_L g7243 ( 
.A(n_6418),
.Y(n_7243)
);

BUFx6f_ASAP7_75t_L g7244 ( 
.A(n_6316),
.Y(n_7244)
);

INVx2_ASAP7_75t_L g7245 ( 
.A(n_6622),
.Y(n_7245)
);

OAI22xp33_ASAP7_75t_L g7246 ( 
.A1(n_6824),
.A2(n_3678),
.B1(n_3679),
.B2(n_3675),
.Y(n_7246)
);

INVx1_ASAP7_75t_L g7247 ( 
.A(n_6419),
.Y(n_7247)
);

HB1xp67_ASAP7_75t_L g7248 ( 
.A(n_6560),
.Y(n_7248)
);

INVx2_ASAP7_75t_L g7249 ( 
.A(n_6627),
.Y(n_7249)
);

INVx4_ASAP7_75t_L g7250 ( 
.A(n_6316),
.Y(n_7250)
);

NAND2xp5_ASAP7_75t_L g7251 ( 
.A(n_6640),
.B(n_3680),
.Y(n_7251)
);

OAI22xp33_ASAP7_75t_L g7252 ( 
.A1(n_6283),
.A2(n_3684),
.B1(n_3685),
.B2(n_3681),
.Y(n_7252)
);

INVx1_ASAP7_75t_L g7253 ( 
.A(n_6420),
.Y(n_7253)
);

INVx2_ASAP7_75t_L g7254 ( 
.A(n_6635),
.Y(n_7254)
);

NAND2xp5_ASAP7_75t_SL g7255 ( 
.A(n_6921),
.B(n_3686),
.Y(n_7255)
);

INVx1_ASAP7_75t_L g7256 ( 
.A(n_6422),
.Y(n_7256)
);

INVx2_ASAP7_75t_L g7257 ( 
.A(n_6638),
.Y(n_7257)
);

INVx2_ASAP7_75t_L g7258 ( 
.A(n_6639),
.Y(n_7258)
);

NAND2xp5_ASAP7_75t_L g7259 ( 
.A(n_6231),
.B(n_3687),
.Y(n_7259)
);

AND2x2_ASAP7_75t_L g7260 ( 
.A(n_6650),
.B(n_3688),
.Y(n_7260)
);

NAND3xp33_ASAP7_75t_L g7261 ( 
.A(n_6236),
.B(n_6532),
.C(n_6455),
.Y(n_7261)
);

BUFx6f_ASAP7_75t_L g7262 ( 
.A(n_6330),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_6423),
.Y(n_7263)
);

INVx3_ASAP7_75t_L g7264 ( 
.A(n_6574),
.Y(n_7264)
);

NAND2xp33_ASAP7_75t_SL g7265 ( 
.A(n_6914),
.B(n_3693),
.Y(n_7265)
);

INVx2_ASAP7_75t_L g7266 ( 
.A(n_6522),
.Y(n_7266)
);

BUFx6f_ASAP7_75t_L g7267 ( 
.A(n_6330),
.Y(n_7267)
);

INVx5_ASAP7_75t_L g7268 ( 
.A(n_6398),
.Y(n_7268)
);

INVx2_ASAP7_75t_L g7269 ( 
.A(n_6541),
.Y(n_7269)
);

BUFx8_ASAP7_75t_SL g7270 ( 
.A(n_6858),
.Y(n_7270)
);

INVx2_ASAP7_75t_L g7271 ( 
.A(n_6542),
.Y(n_7271)
);

INVx2_ASAP7_75t_L g7272 ( 
.A(n_6547),
.Y(n_7272)
);

AOI22xp33_ASAP7_75t_L g7273 ( 
.A1(n_6906),
.A2(n_3697),
.B1(n_3698),
.B2(n_3694),
.Y(n_7273)
);

NAND2xp33_ASAP7_75t_L g7274 ( 
.A(n_6923),
.B(n_6926),
.Y(n_7274)
);

INVx2_ASAP7_75t_L g7275 ( 
.A(n_6550),
.Y(n_7275)
);

AOI22xp33_ASAP7_75t_L g7276 ( 
.A1(n_6523),
.A2(n_6694),
.B1(n_6866),
.B2(n_6580),
.Y(n_7276)
);

NAND2xp5_ASAP7_75t_L g7277 ( 
.A(n_6521),
.B(n_3699),
.Y(n_7277)
);

NAND2xp33_ASAP7_75t_L g7278 ( 
.A(n_6477),
.B(n_3700),
.Y(n_7278)
);

INVx2_ASAP7_75t_L g7279 ( 
.A(n_6553),
.Y(n_7279)
);

NAND2xp5_ASAP7_75t_L g7280 ( 
.A(n_6641),
.B(n_3702),
.Y(n_7280)
);

BUFx3_ASAP7_75t_L g7281 ( 
.A(n_6210),
.Y(n_7281)
);

INVx2_ASAP7_75t_L g7282 ( 
.A(n_6556),
.Y(n_7282)
);

NAND2xp5_ASAP7_75t_L g7283 ( 
.A(n_6642),
.B(n_3704),
.Y(n_7283)
);

INVx1_ASAP7_75t_L g7284 ( 
.A(n_6427),
.Y(n_7284)
);

INVx2_ASAP7_75t_L g7285 ( 
.A(n_6563),
.Y(n_7285)
);

AO21x2_ASAP7_75t_L g7286 ( 
.A1(n_6805),
.A2(n_3642),
.B(n_3641),
.Y(n_7286)
);

INVx2_ASAP7_75t_L g7287 ( 
.A(n_6565),
.Y(n_7287)
);

NAND2xp5_ASAP7_75t_SL g7288 ( 
.A(n_6810),
.B(n_6854),
.Y(n_7288)
);

INVx1_ASAP7_75t_L g7289 ( 
.A(n_6429),
.Y(n_7289)
);

INVx2_ASAP7_75t_L g7290 ( 
.A(n_6572),
.Y(n_7290)
);

INVx2_ASAP7_75t_SL g7291 ( 
.A(n_6349),
.Y(n_7291)
);

NAND3xp33_ASAP7_75t_L g7292 ( 
.A(n_6528),
.B(n_3706),
.C(n_3705),
.Y(n_7292)
);

NAND3xp33_ASAP7_75t_L g7293 ( 
.A(n_6911),
.B(n_3711),
.C(n_3708),
.Y(n_7293)
);

NAND2xp5_ASAP7_75t_L g7294 ( 
.A(n_6649),
.B(n_3712),
.Y(n_7294)
);

NAND2xp5_ASAP7_75t_SL g7295 ( 
.A(n_6859),
.B(n_3714),
.Y(n_7295)
);

NAND2xp5_ASAP7_75t_L g7296 ( 
.A(n_6654),
.B(n_3715),
.Y(n_7296)
);

AOI22xp33_ASAP7_75t_L g7297 ( 
.A1(n_6594),
.A2(n_3717),
.B1(n_3718),
.B2(n_3716),
.Y(n_7297)
);

INVx2_ASAP7_75t_L g7298 ( 
.A(n_6577),
.Y(n_7298)
);

CKINVDCx16_ASAP7_75t_R g7299 ( 
.A(n_6890),
.Y(n_7299)
);

NAND2xp5_ASAP7_75t_L g7300 ( 
.A(n_6655),
.B(n_3720),
.Y(n_7300)
);

NAND2xp5_ASAP7_75t_SL g7301 ( 
.A(n_6873),
.B(n_3721),
.Y(n_7301)
);

INVx1_ASAP7_75t_L g7302 ( 
.A(n_6431),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_6434),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_6435),
.Y(n_7304)
);

INVx2_ASAP7_75t_L g7305 ( 
.A(n_6578),
.Y(n_7305)
);

INVx2_ASAP7_75t_L g7306 ( 
.A(n_6579),
.Y(n_7306)
);

INVx2_ASAP7_75t_L g7307 ( 
.A(n_6581),
.Y(n_7307)
);

INVx1_ASAP7_75t_L g7308 ( 
.A(n_6439),
.Y(n_7308)
);

INVx2_ASAP7_75t_SL g7309 ( 
.A(n_6403),
.Y(n_7309)
);

INVx1_ASAP7_75t_L g7310 ( 
.A(n_6440),
.Y(n_7310)
);

AOI22xp33_ASAP7_75t_SL g7311 ( 
.A1(n_6219),
.A2(n_6410),
.B1(n_6882),
.B2(n_6856),
.Y(n_7311)
);

NOR2xp33_ASAP7_75t_L g7312 ( 
.A(n_6801),
.B(n_3724),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_6441),
.Y(n_7313)
);

NOR2xp33_ASAP7_75t_L g7314 ( 
.A(n_6653),
.B(n_3727),
.Y(n_7314)
);

INVxp67_ASAP7_75t_L g7315 ( 
.A(n_6444),
.Y(n_7315)
);

INVx2_ASAP7_75t_SL g7316 ( 
.A(n_6450),
.Y(n_7316)
);

INVx1_ASAP7_75t_L g7317 ( 
.A(n_6443),
.Y(n_7317)
);

INVx3_ASAP7_75t_L g7318 ( 
.A(n_6537),
.Y(n_7318)
);

INVx2_ASAP7_75t_SL g7319 ( 
.A(n_6473),
.Y(n_7319)
);

INVx2_ASAP7_75t_L g7320 ( 
.A(n_6582),
.Y(n_7320)
);

INVx1_ASAP7_75t_L g7321 ( 
.A(n_6447),
.Y(n_7321)
);

NOR2xp33_ASAP7_75t_L g7322 ( 
.A(n_6688),
.B(n_3728),
.Y(n_7322)
);

NAND2xp5_ASAP7_75t_SL g7323 ( 
.A(n_6569),
.B(n_3733),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_6452),
.Y(n_7324)
);

INVx1_ASAP7_75t_L g7325 ( 
.A(n_6453),
.Y(n_7325)
);

NAND3xp33_ASAP7_75t_L g7326 ( 
.A(n_6384),
.B(n_3738),
.C(n_3737),
.Y(n_7326)
);

INVx2_ASAP7_75t_L g7327 ( 
.A(n_6584),
.Y(n_7327)
);

BUFx6f_ASAP7_75t_L g7328 ( 
.A(n_6210),
.Y(n_7328)
);

INVx1_ASAP7_75t_L g7329 ( 
.A(n_6464),
.Y(n_7329)
);

INVx1_ASAP7_75t_L g7330 ( 
.A(n_6465),
.Y(n_7330)
);

NAND2xp5_ASAP7_75t_SL g7331 ( 
.A(n_6551),
.B(n_3739),
.Y(n_7331)
);

CKINVDCx5p33_ASAP7_75t_R g7332 ( 
.A(n_6488),
.Y(n_7332)
);

NAND2xp5_ASAP7_75t_L g7333 ( 
.A(n_6215),
.B(n_3740),
.Y(n_7333)
);

NAND2xp5_ASAP7_75t_SL g7334 ( 
.A(n_6561),
.B(n_3742),
.Y(n_7334)
);

INVx1_ASAP7_75t_L g7335 ( 
.A(n_6466),
.Y(n_7335)
);

INVx1_ASAP7_75t_L g7336 ( 
.A(n_6471),
.Y(n_7336)
);

INVx1_ASAP7_75t_L g7337 ( 
.A(n_6476),
.Y(n_7337)
);

INVx2_ASAP7_75t_L g7338 ( 
.A(n_6585),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_6478),
.Y(n_7339)
);

INVx2_ASAP7_75t_L g7340 ( 
.A(n_6586),
.Y(n_7340)
);

INVx4_ASAP7_75t_L g7341 ( 
.A(n_6750),
.Y(n_7341)
);

INVx2_ASAP7_75t_L g7342 ( 
.A(n_6591),
.Y(n_7342)
);

INVx1_ASAP7_75t_L g7343 ( 
.A(n_6479),
.Y(n_7343)
);

AOI22xp5_ASAP7_75t_L g7344 ( 
.A1(n_6786),
.A2(n_3747),
.B1(n_3748),
.B2(n_3745),
.Y(n_7344)
);

NAND2xp5_ASAP7_75t_SL g7345 ( 
.A(n_6758),
.B(n_3750),
.Y(n_7345)
);

NAND2xp5_ASAP7_75t_SL g7346 ( 
.A(n_6346),
.B(n_3752),
.Y(n_7346)
);

INVx2_ASAP7_75t_L g7347 ( 
.A(n_6593),
.Y(n_7347)
);

INVxp67_ASAP7_75t_SL g7348 ( 
.A(n_6652),
.Y(n_7348)
);

INVx2_ASAP7_75t_L g7349 ( 
.A(n_6597),
.Y(n_7349)
);

NAND3xp33_ASAP7_75t_L g7350 ( 
.A(n_6559),
.B(n_3755),
.C(n_3754),
.Y(n_7350)
);

INVx2_ASAP7_75t_L g7351 ( 
.A(n_6600),
.Y(n_7351)
);

NAND2xp5_ASAP7_75t_SL g7352 ( 
.A(n_6718),
.B(n_3756),
.Y(n_7352)
);

AND2x2_ASAP7_75t_L g7353 ( 
.A(n_6599),
.B(n_6626),
.Y(n_7353)
);

INVx2_ASAP7_75t_SL g7354 ( 
.A(n_6538),
.Y(n_7354)
);

INVx5_ASAP7_75t_L g7355 ( 
.A(n_6398),
.Y(n_7355)
);

INVx1_ASAP7_75t_L g7356 ( 
.A(n_6480),
.Y(n_7356)
);

INVx2_ASAP7_75t_L g7357 ( 
.A(n_6602),
.Y(n_7357)
);

NAND2xp5_ASAP7_75t_L g7358 ( 
.A(n_6723),
.B(n_3757),
.Y(n_7358)
);

INVx1_ASAP7_75t_L g7359 ( 
.A(n_6481),
.Y(n_7359)
);

NAND2xp33_ASAP7_75t_L g7360 ( 
.A(n_6731),
.B(n_3758),
.Y(n_7360)
);

INVx1_ASAP7_75t_L g7361 ( 
.A(n_6486),
.Y(n_7361)
);

AND2x4_ASAP7_75t_L g7362 ( 
.A(n_6332),
.B(n_3645),
.Y(n_7362)
);

BUFx8_ASAP7_75t_SL g7363 ( 
.A(n_6781),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_6490),
.Y(n_7364)
);

NAND2xp5_ASAP7_75t_L g7365 ( 
.A(n_6736),
.B(n_3761),
.Y(n_7365)
);

INVx2_ASAP7_75t_L g7366 ( 
.A(n_6603),
.Y(n_7366)
);

NAND2xp5_ASAP7_75t_SL g7367 ( 
.A(n_6739),
.B(n_3762),
.Y(n_7367)
);

BUFx10_ASAP7_75t_L g7368 ( 
.A(n_6402),
.Y(n_7368)
);

AND2x2_ASAP7_75t_L g7369 ( 
.A(n_6637),
.B(n_3763),
.Y(n_7369)
);

AOI22xp33_ASAP7_75t_L g7370 ( 
.A1(n_6644),
.A2(n_3768),
.B1(n_3772),
.B2(n_3764),
.Y(n_7370)
);

NOR2xp33_ASAP7_75t_L g7371 ( 
.A(n_6915),
.B(n_3773),
.Y(n_7371)
);

NOR2xp33_ASAP7_75t_L g7372 ( 
.A(n_6823),
.B(n_3776),
.Y(n_7372)
);

INVx2_ASAP7_75t_L g7373 ( 
.A(n_6604),
.Y(n_7373)
);

INVx2_ASAP7_75t_L g7374 ( 
.A(n_6646),
.Y(n_7374)
);

NAND2xp5_ASAP7_75t_SL g7375 ( 
.A(n_6740),
.B(n_3777),
.Y(n_7375)
);

BUFx6f_ASAP7_75t_SL g7376 ( 
.A(n_6402),
.Y(n_7376)
);

AO22x2_ASAP7_75t_L g7377 ( 
.A1(n_6878),
.A2(n_3650),
.B1(n_3654),
.B2(n_3648),
.Y(n_7377)
);

BUFx6f_ASAP7_75t_L g7378 ( 
.A(n_6212),
.Y(n_7378)
);

BUFx6f_ASAP7_75t_L g7379 ( 
.A(n_6212),
.Y(n_7379)
);

INVx2_ASAP7_75t_L g7380 ( 
.A(n_6648),
.Y(n_7380)
);

INVx2_ASAP7_75t_L g7381 ( 
.A(n_6662),
.Y(n_7381)
);

INVx1_ASAP7_75t_L g7382 ( 
.A(n_6491),
.Y(n_7382)
);

INVx1_ASAP7_75t_L g7383 ( 
.A(n_6493),
.Y(n_7383)
);

INVx2_ASAP7_75t_L g7384 ( 
.A(n_6667),
.Y(n_7384)
);

AND2x2_ASAP7_75t_SL g7385 ( 
.A(n_6943),
.B(n_3827),
.Y(n_7385)
);

INVx1_ASAP7_75t_L g7386 ( 
.A(n_6494),
.Y(n_7386)
);

NAND2xp5_ASAP7_75t_SL g7387 ( 
.A(n_6744),
.B(n_3778),
.Y(n_7387)
);

INVx1_ASAP7_75t_SL g7388 ( 
.A(n_6566),
.Y(n_7388)
);

AND2x6_ASAP7_75t_L g7389 ( 
.A(n_6855),
.B(n_6856),
.Y(n_7389)
);

NAND2xp5_ASAP7_75t_L g7390 ( 
.A(n_6746),
.B(n_3779),
.Y(n_7390)
);

INVx1_ASAP7_75t_L g7391 ( 
.A(n_6503),
.Y(n_7391)
);

INVx2_ASAP7_75t_L g7392 ( 
.A(n_6673),
.Y(n_7392)
);

INVx1_ASAP7_75t_L g7393 ( 
.A(n_6505),
.Y(n_7393)
);

INVxp33_ASAP7_75t_L g7394 ( 
.A(n_6567),
.Y(n_7394)
);

INVx1_ASAP7_75t_L g7395 ( 
.A(n_6511),
.Y(n_7395)
);

CKINVDCx5p33_ASAP7_75t_R g7396 ( 
.A(n_6555),
.Y(n_7396)
);

NOR2xp33_ASAP7_75t_SL g7397 ( 
.A(n_6770),
.B(n_3780),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_6512),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_6516),
.Y(n_7399)
);

NAND2xp33_ASAP7_75t_SL g7400 ( 
.A(n_6378),
.B(n_3781),
.Y(n_7400)
);

NAND2xp5_ASAP7_75t_SL g7401 ( 
.A(n_6749),
.B(n_3782),
.Y(n_7401)
);

BUFx6f_ASAP7_75t_L g7402 ( 
.A(n_6213),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_6517),
.Y(n_7403)
);

INVx1_ASAP7_75t_L g7404 ( 
.A(n_6703),
.Y(n_7404)
);

INVx2_ASAP7_75t_L g7405 ( 
.A(n_6675),
.Y(n_7405)
);

INVx2_ASAP7_75t_L g7406 ( 
.A(n_6676),
.Y(n_7406)
);

INVx2_ASAP7_75t_L g7407 ( 
.A(n_6682),
.Y(n_7407)
);

CKINVDCx5p33_ASAP7_75t_R g7408 ( 
.A(n_6629),
.Y(n_7408)
);

CKINVDCx5p33_ASAP7_75t_R g7409 ( 
.A(n_6647),
.Y(n_7409)
);

INVx5_ASAP7_75t_L g7410 ( 
.A(n_6483),
.Y(n_7410)
);

INVxp33_ASAP7_75t_L g7411 ( 
.A(n_6576),
.Y(n_7411)
);

AOI22xp33_ASAP7_75t_L g7412 ( 
.A1(n_6894),
.A2(n_3784),
.B1(n_3785),
.B2(n_3783),
.Y(n_7412)
);

BUFx6f_ASAP7_75t_L g7413 ( 
.A(n_6213),
.Y(n_7413)
);

NAND2xp5_ASAP7_75t_SL g7414 ( 
.A(n_6755),
.B(n_3788),
.Y(n_7414)
);

INVx2_ASAP7_75t_L g7415 ( 
.A(n_6683),
.Y(n_7415)
);

BUFx6f_ASAP7_75t_L g7416 ( 
.A(n_6221),
.Y(n_7416)
);

AOI22xp33_ASAP7_75t_L g7417 ( 
.A1(n_6896),
.A2(n_3793),
.B1(n_3795),
.B2(n_3790),
.Y(n_7417)
);

NOR2xp33_ASAP7_75t_L g7418 ( 
.A(n_6828),
.B(n_3797),
.Y(n_7418)
);

INVx2_ASAP7_75t_L g7419 ( 
.A(n_6686),
.Y(n_7419)
);

INVx4_ASAP7_75t_L g7420 ( 
.A(n_6221),
.Y(n_7420)
);

INVxp67_ASAP7_75t_SL g7421 ( 
.A(n_6656),
.Y(n_7421)
);

OAI22xp33_ASAP7_75t_L g7422 ( 
.A1(n_6937),
.A2(n_3803),
.B1(n_3806),
.B2(n_3802),
.Y(n_7422)
);

INVx2_ASAP7_75t_L g7423 ( 
.A(n_6700),
.Y(n_7423)
);

NAND3xp33_ASAP7_75t_L g7424 ( 
.A(n_6867),
.B(n_3809),
.C(n_3807),
.Y(n_7424)
);

AOI22xp5_ASAP7_75t_L g7425 ( 
.A1(n_6658),
.A2(n_3811),
.B1(n_3816),
.B2(n_3810),
.Y(n_7425)
);

INVx2_ASAP7_75t_L g7426 ( 
.A(n_6705),
.Y(n_7426)
);

INVx2_ASAP7_75t_L g7427 ( 
.A(n_6336),
.Y(n_7427)
);

INVx1_ASAP7_75t_SL g7428 ( 
.A(n_6595),
.Y(n_7428)
);

INVx2_ASAP7_75t_L g7429 ( 
.A(n_6339),
.Y(n_7429)
);

BUFx6f_ASAP7_75t_L g7430 ( 
.A(n_6222),
.Y(n_7430)
);

OAI22xp33_ASAP7_75t_L g7431 ( 
.A1(n_6918),
.A2(n_3826),
.B1(n_3828),
.B2(n_3819),
.Y(n_7431)
);

NOR2xp33_ASAP7_75t_L g7432 ( 
.A(n_6851),
.B(n_6868),
.Y(n_7432)
);

INVx2_ASAP7_75t_L g7433 ( 
.A(n_6344),
.Y(n_7433)
);

INVx2_ASAP7_75t_SL g7434 ( 
.A(n_6197),
.Y(n_7434)
);

INVx1_ASAP7_75t_L g7435 ( 
.A(n_6707),
.Y(n_7435)
);

BUFx6f_ASAP7_75t_L g7436 ( 
.A(n_6222),
.Y(n_7436)
);

AOI22xp33_ASAP7_75t_L g7437 ( 
.A1(n_6932),
.A2(n_3830),
.B1(n_3831),
.B2(n_3829),
.Y(n_7437)
);

INVx1_ASAP7_75t_L g7438 ( 
.A(n_6708),
.Y(n_7438)
);

INVx2_ASAP7_75t_L g7439 ( 
.A(n_6347),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_6710),
.Y(n_7440)
);

AOI22xp5_ASAP7_75t_L g7441 ( 
.A1(n_6665),
.A2(n_3834),
.B1(n_3836),
.B2(n_3832),
.Y(n_7441)
);

INVx2_ASAP7_75t_L g7442 ( 
.A(n_6350),
.Y(n_7442)
);

NAND2xp33_ASAP7_75t_L g7443 ( 
.A(n_6757),
.B(n_3838),
.Y(n_7443)
);

INVx2_ASAP7_75t_L g7444 ( 
.A(n_6353),
.Y(n_7444)
);

BUFx6f_ASAP7_75t_SL g7445 ( 
.A(n_6483),
.Y(n_7445)
);

AND2x2_ASAP7_75t_SL g7446 ( 
.A(n_6882),
.B(n_3859),
.Y(n_7446)
);

AND2x2_ASAP7_75t_L g7447 ( 
.A(n_6335),
.B(n_6218),
.Y(n_7447)
);

INVx1_ASAP7_75t_L g7448 ( 
.A(n_6712),
.Y(n_7448)
);

INVx1_ASAP7_75t_L g7449 ( 
.A(n_6713),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_6871),
.Y(n_7450)
);

INVx1_ASAP7_75t_L g7451 ( 
.A(n_6869),
.Y(n_7451)
);

INVx2_ASAP7_75t_L g7452 ( 
.A(n_6361),
.Y(n_7452)
);

NAND2xp5_ASAP7_75t_SL g7453 ( 
.A(n_6759),
.B(n_3839),
.Y(n_7453)
);

INVx2_ASAP7_75t_L g7454 ( 
.A(n_6368),
.Y(n_7454)
);

OR2x2_ASAP7_75t_L g7455 ( 
.A(n_6587),
.B(n_3841),
.Y(n_7455)
);

INVx2_ASAP7_75t_L g7456 ( 
.A(n_6371),
.Y(n_7456)
);

NAND2xp5_ASAP7_75t_L g7457 ( 
.A(n_6766),
.B(n_3842),
.Y(n_7457)
);

NAND2xp5_ASAP7_75t_SL g7458 ( 
.A(n_6669),
.B(n_3847),
.Y(n_7458)
);

NAND2xp5_ASAP7_75t_SL g7459 ( 
.A(n_6259),
.B(n_3850),
.Y(n_7459)
);

INVx5_ASAP7_75t_L g7460 ( 
.A(n_6544),
.Y(n_7460)
);

AOI22xp33_ASAP7_75t_SL g7461 ( 
.A1(n_6900),
.A2(n_3852),
.B1(n_3853),
.B2(n_3851),
.Y(n_7461)
);

NOR2xp33_ASAP7_75t_L g7462 ( 
.A(n_6884),
.B(n_3854),
.Y(n_7462)
);

INVx1_ASAP7_75t_L g7463 ( 
.A(n_6872),
.Y(n_7463)
);

AND2x6_ASAP7_75t_L g7464 ( 
.A(n_6900),
.B(n_3659),
.Y(n_7464)
);

HB1xp67_ASAP7_75t_L g7465 ( 
.A(n_6636),
.Y(n_7465)
);

INVx1_ASAP7_75t_L g7466 ( 
.A(n_6874),
.Y(n_7466)
);

INVx1_ASAP7_75t_L g7467 ( 
.A(n_6373),
.Y(n_7467)
);

BUFx3_ASAP7_75t_L g7468 ( 
.A(n_6227),
.Y(n_7468)
);

NAND2xp5_ASAP7_75t_SL g7469 ( 
.A(n_6199),
.B(n_3855),
.Y(n_7469)
);

INVx2_ASAP7_75t_L g7470 ( 
.A(n_6391),
.Y(n_7470)
);

NAND2xp5_ASAP7_75t_L g7471 ( 
.A(n_6634),
.B(n_6668),
.Y(n_7471)
);

INVxp33_ASAP7_75t_SL g7472 ( 
.A(n_6660),
.Y(n_7472)
);

INVx2_ASAP7_75t_L g7473 ( 
.A(n_6394),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_6714),
.Y(n_7474)
);

INVx3_ASAP7_75t_L g7475 ( 
.A(n_6227),
.Y(n_7475)
);

OAI22xp33_ASAP7_75t_L g7476 ( 
.A1(n_6207),
.A2(n_3857),
.B1(n_3863),
.B2(n_3856),
.Y(n_7476)
);

BUFx6f_ASAP7_75t_SL g7477 ( 
.A(n_6544),
.Y(n_7477)
);

INVx2_ASAP7_75t_L g7478 ( 
.A(n_6715),
.Y(n_7478)
);

INVx2_ASAP7_75t_L g7479 ( 
.A(n_6716),
.Y(n_7479)
);

INVx1_ASAP7_75t_L g7480 ( 
.A(n_6720),
.Y(n_7480)
);

NOR2xp33_ASAP7_75t_L g7481 ( 
.A(n_6892),
.B(n_3864),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_6607),
.Y(n_7482)
);

NAND2xp5_ASAP7_75t_SL g7483 ( 
.A(n_6951),
.B(n_3868),
.Y(n_7483)
);

INVx2_ASAP7_75t_L g7484 ( 
.A(n_6272),
.Y(n_7484)
);

INVx2_ASAP7_75t_SL g7485 ( 
.A(n_6950),
.Y(n_7485)
);

INVx4_ASAP7_75t_L g7486 ( 
.A(n_6234),
.Y(n_7486)
);

NAND2xp5_ASAP7_75t_SL g7487 ( 
.A(n_6401),
.B(n_3869),
.Y(n_7487)
);

INVx2_ASAP7_75t_L g7488 ( 
.A(n_6698),
.Y(n_7488)
);

INVx3_ASAP7_75t_L g7489 ( 
.A(n_6234),
.Y(n_7489)
);

NAND3xp33_ASAP7_75t_L g7490 ( 
.A(n_6835),
.B(n_3875),
.C(n_3872),
.Y(n_7490)
);

INVx3_ASAP7_75t_L g7491 ( 
.A(n_6239),
.Y(n_7491)
);

NAND2xp5_ASAP7_75t_SL g7492 ( 
.A(n_6502),
.B(n_3876),
.Y(n_7492)
);

AND2x2_ASAP7_75t_L g7493 ( 
.A(n_6363),
.B(n_6364),
.Y(n_7493)
);

NOR2xp33_ASAP7_75t_L g7494 ( 
.A(n_6760),
.B(n_3877),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_6889),
.Y(n_7495)
);

INVx2_ASAP7_75t_L g7496 ( 
.A(n_6701),
.Y(n_7496)
);

INVx2_ASAP7_75t_L g7497 ( 
.A(n_6769),
.Y(n_7497)
);

INVx4_ASAP7_75t_L g7498 ( 
.A(n_6239),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_6780),
.Y(n_7499)
);

INVx2_ASAP7_75t_L g7500 ( 
.A(n_6775),
.Y(n_7500)
);

INVx2_ASAP7_75t_SL g7501 ( 
.A(n_6730),
.Y(n_7501)
);

NOR2xp33_ASAP7_75t_L g7502 ( 
.A(n_6771),
.B(n_3878),
.Y(n_7502)
);

INVxp33_ASAP7_75t_L g7503 ( 
.A(n_6806),
.Y(n_7503)
);

INVx2_ASAP7_75t_L g7504 ( 
.A(n_6778),
.Y(n_7504)
);

INVx2_ASAP7_75t_L g7505 ( 
.A(n_6809),
.Y(n_7505)
);

INVx2_ASAP7_75t_L g7506 ( 
.A(n_6812),
.Y(n_7506)
);

INVx1_ASAP7_75t_L g7507 ( 
.A(n_6782),
.Y(n_7507)
);

CKINVDCx5p33_ASAP7_75t_R g7508 ( 
.A(n_6798),
.Y(n_7508)
);

INVx2_ASAP7_75t_L g7509 ( 
.A(n_6816),
.Y(n_7509)
);

NAND2xp5_ASAP7_75t_L g7510 ( 
.A(n_6696),
.B(n_3885),
.Y(n_7510)
);

NAND2xp5_ASAP7_75t_L g7511 ( 
.A(n_6616),
.B(n_3886),
.Y(n_7511)
);

NAND3xp33_ASAP7_75t_L g7512 ( 
.A(n_6725),
.B(n_3888),
.C(n_3887),
.Y(n_7512)
);

AOI22xp5_ASAP7_75t_L g7513 ( 
.A1(n_6825),
.A2(n_3889),
.B1(n_3892),
.B2(n_3890),
.Y(n_7513)
);

AND3x2_ASAP7_75t_L g7514 ( 
.A(n_6913),
.B(n_3979),
.C(n_3861),
.Y(n_7514)
);

INVx5_ASAP7_75t_L g7515 ( 
.A(n_6251),
.Y(n_7515)
);

INVx2_ASAP7_75t_L g7516 ( 
.A(n_6817),
.Y(n_7516)
);

NAND2xp5_ASAP7_75t_L g7517 ( 
.A(n_6619),
.B(n_3893),
.Y(n_7517)
);

OAI22xp33_ASAP7_75t_L g7518 ( 
.A1(n_6870),
.A2(n_6857),
.B1(n_6865),
.B2(n_6830),
.Y(n_7518)
);

BUFx6f_ASAP7_75t_SL g7519 ( 
.A(n_6938),
.Y(n_7519)
);

BUFx3_ASAP7_75t_L g7520 ( 
.A(n_6251),
.Y(n_7520)
);

INVx2_ASAP7_75t_L g7521 ( 
.A(n_6818),
.Y(n_7521)
);

INVx4_ASAP7_75t_L g7522 ( 
.A(n_6948),
.Y(n_7522)
);

NAND2xp5_ASAP7_75t_L g7523 ( 
.A(n_6621),
.B(n_3895),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_6787),
.Y(n_7524)
);

INVx3_ASAP7_75t_L g7525 ( 
.A(n_6948),
.Y(n_7525)
);

INVx8_ASAP7_75t_L g7526 ( 
.A(n_6226),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_6794),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_6795),
.Y(n_7528)
);

INVx1_ASAP7_75t_L g7529 ( 
.A(n_6799),
.Y(n_7529)
);

INVx1_ASAP7_75t_L g7530 ( 
.A(n_6800),
.Y(n_7530)
);

INVx2_ASAP7_75t_L g7531 ( 
.A(n_6820),
.Y(n_7531)
);

INVx2_ASAP7_75t_L g7532 ( 
.A(n_6821),
.Y(n_7532)
);

INVxp33_ASAP7_75t_L g7533 ( 
.A(n_6232),
.Y(n_7533)
);

BUFx2_ASAP7_75t_L g7534 ( 
.A(n_6475),
.Y(n_7534)
);

INVx1_ASAP7_75t_L g7535 ( 
.A(n_6679),
.Y(n_7535)
);

INVx4_ASAP7_75t_L g7536 ( 
.A(n_6273),
.Y(n_7536)
);

INVx2_ASAP7_75t_L g7537 ( 
.A(n_6540),
.Y(n_7537)
);

AOI21x1_ASAP7_75t_L g7538 ( 
.A1(n_6195),
.A2(n_3666),
.B(n_3662),
.Y(n_7538)
);

INVx1_ASAP7_75t_L g7539 ( 
.A(n_6680),
.Y(n_7539)
);

INVx1_ASAP7_75t_L g7540 ( 
.A(n_6690),
.Y(n_7540)
);

NOR3xp33_ASAP7_75t_L g7541 ( 
.A(n_6216),
.B(n_2767),
.C(n_2734),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_6695),
.Y(n_7542)
);

NAND2xp33_ASAP7_75t_L g7543 ( 
.A(n_6625),
.B(n_3896),
.Y(n_7543)
);

INVx2_ASAP7_75t_L g7544 ( 
.A(n_6726),
.Y(n_7544)
);

AOI21x1_ASAP7_75t_L g7545 ( 
.A1(n_6827),
.A2(n_6411),
.B(n_6269),
.Y(n_7545)
);

INVx3_ASAP7_75t_L g7546 ( 
.A(n_6273),
.Y(n_7546)
);

INVx1_ASAP7_75t_L g7547 ( 
.A(n_6853),
.Y(n_7547)
);

INVx2_ASAP7_75t_L g7548 ( 
.A(n_6741),
.Y(n_7548)
);

NAND2xp5_ASAP7_75t_L g7549 ( 
.A(n_6630),
.B(n_3898),
.Y(n_7549)
);

NAND2xp5_ASAP7_75t_L g7550 ( 
.A(n_6496),
.B(n_3902),
.Y(n_7550)
);

INVx1_ASAP7_75t_L g7551 ( 
.A(n_6852),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_6908),
.Y(n_7552)
);

NOR2xp33_ASAP7_75t_L g7553 ( 
.A(n_6260),
.B(n_3905),
.Y(n_7553)
);

INVx5_ASAP7_75t_L g7554 ( 
.A(n_6413),
.Y(n_7554)
);

INVx3_ASAP7_75t_L g7555 ( 
.A(n_6291),
.Y(n_7555)
);

INVx5_ASAP7_75t_L g7556 ( 
.A(n_6291),
.Y(n_7556)
);

BUFx2_ASAP7_75t_L g7557 ( 
.A(n_6643),
.Y(n_7557)
);

NAND2xp5_ASAP7_75t_L g7558 ( 
.A(n_6501),
.B(n_3908),
.Y(n_7558)
);

AND2x6_ASAP7_75t_L g7559 ( 
.A(n_6881),
.B(n_3676),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_6381),
.Y(n_7560)
);

INVx2_ASAP7_75t_L g7561 ( 
.A(n_6557),
.Y(n_7561)
);

BUFx2_ASAP7_75t_L g7562 ( 
.A(n_6358),
.Y(n_7562)
);

INVx2_ASAP7_75t_L g7563 ( 
.A(n_6633),
.Y(n_7563)
);

BUFx2_ASAP7_75t_L g7564 ( 
.A(n_6399),
.Y(n_7564)
);

BUFx10_ASAP7_75t_L g7565 ( 
.A(n_6693),
.Y(n_7565)
);

INVx2_ASAP7_75t_L g7566 ( 
.A(n_6734),
.Y(n_7566)
);

INVx3_ASAP7_75t_L g7567 ( 
.A(n_6722),
.Y(n_7567)
);

INVx2_ASAP7_75t_L g7568 ( 
.A(n_6738),
.Y(n_7568)
);

NAND2xp33_ASAP7_75t_L g7569 ( 
.A(n_6255),
.B(n_3909),
.Y(n_7569)
);

INVx2_ASAP7_75t_SL g7570 ( 
.A(n_6722),
.Y(n_7570)
);

INVxp67_ASAP7_75t_SL g7571 ( 
.A(n_6229),
.Y(n_7571)
);

INVx3_ASAP7_75t_L g7572 ( 
.A(n_6728),
.Y(n_7572)
);

AND2x2_ASAP7_75t_SL g7573 ( 
.A(n_6193),
.B(n_3997),
.Y(n_7573)
);

INVx2_ASAP7_75t_L g7574 ( 
.A(n_6747),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_6314),
.Y(n_7575)
);

INVx2_ASAP7_75t_L g7576 ( 
.A(n_6748),
.Y(n_7576)
);

AND2x2_ASAP7_75t_L g7577 ( 
.A(n_6428),
.B(n_3910),
.Y(n_7577)
);

BUFx6f_ASAP7_75t_SL g7578 ( 
.A(n_6938),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_6337),
.Y(n_7579)
);

NAND2xp5_ASAP7_75t_L g7580 ( 
.A(n_6508),
.B(n_3912),
.Y(n_7580)
);

OR2x6_ASAP7_75t_L g7581 ( 
.A(n_6860),
.B(n_4017),
.Y(n_7581)
);

INVx2_ASAP7_75t_SL g7582 ( 
.A(n_6728),
.Y(n_7582)
);

INVx2_ASAP7_75t_L g7583 ( 
.A(n_6756),
.Y(n_7583)
);

NOR2x1p5_ASAP7_75t_L g7584 ( 
.A(n_6235),
.B(n_3913),
.Y(n_7584)
);

AND2x2_ASAP7_75t_L g7585 ( 
.A(n_6497),
.B(n_3914),
.Y(n_7585)
);

INVx3_ASAP7_75t_L g7586 ( 
.A(n_6729),
.Y(n_7586)
);

AND2x2_ASAP7_75t_L g7587 ( 
.A(n_6499),
.B(n_3917),
.Y(n_7587)
);

INVxp67_ASAP7_75t_SL g7588 ( 
.A(n_6504),
.Y(n_7588)
);

OAI22xp33_ASAP7_75t_SL g7589 ( 
.A1(n_6946),
.A2(n_6208),
.B1(n_6862),
.B2(n_6861),
.Y(n_7589)
);

CKINVDCx20_ASAP7_75t_R g7590 ( 
.A(n_6489),
.Y(n_7590)
);

INVx2_ASAP7_75t_L g7591 ( 
.A(n_6762),
.Y(n_7591)
);

AND2x2_ASAP7_75t_SL g7592 ( 
.A(n_6901),
.B(n_6941),
.Y(n_7592)
);

OR2x6_ASAP7_75t_L g7593 ( 
.A(n_6864),
.B(n_4028),
.Y(n_7593)
);

INVx1_ASAP7_75t_L g7594 ( 
.A(n_6340),
.Y(n_7594)
);

AND2x2_ASAP7_75t_L g7595 ( 
.A(n_6514),
.B(n_3918),
.Y(n_7595)
);

NAND2xp5_ASAP7_75t_L g7596 ( 
.A(n_6510),
.B(n_3919),
.Y(n_7596)
);

INVx4_ASAP7_75t_L g7597 ( 
.A(n_6729),
.Y(n_7597)
);

INVx2_ASAP7_75t_L g7598 ( 
.A(n_6764),
.Y(n_7598)
);

INVx1_ASAP7_75t_L g7599 ( 
.A(n_6342),
.Y(n_7599)
);

OR2x2_ASAP7_75t_L g7600 ( 
.A(n_6724),
.B(n_3921),
.Y(n_7600)
);

AOI22xp33_ASAP7_75t_L g7601 ( 
.A1(n_6763),
.A2(n_3924),
.B1(n_3925),
.B2(n_3922),
.Y(n_7601)
);

INVx3_ASAP7_75t_L g7602 ( 
.A(n_6735),
.Y(n_7602)
);

NOR2xp33_ASAP7_75t_L g7603 ( 
.A(n_6370),
.B(n_3928),
.Y(n_7603)
);

NOR2xp33_ASAP7_75t_SL g7604 ( 
.A(n_6684),
.B(n_3931),
.Y(n_7604)
);

INVx1_ASAP7_75t_L g7605 ( 
.A(n_6348),
.Y(n_7605)
);

AOI22xp33_ASAP7_75t_L g7606 ( 
.A1(n_6888),
.A2(n_3934),
.B1(n_3936),
.B2(n_3932),
.Y(n_7606)
);

INVx1_ASAP7_75t_L g7607 ( 
.A(n_6351),
.Y(n_7607)
);

INVx1_ASAP7_75t_L g7608 ( 
.A(n_6360),
.Y(n_7608)
);

BUFx3_ASAP7_75t_L g7609 ( 
.A(n_6735),
.Y(n_7609)
);

AND2x2_ASAP7_75t_SL g7610 ( 
.A(n_6942),
.B(n_3682),
.Y(n_7610)
);

NAND2xp5_ASAP7_75t_L g7611 ( 
.A(n_6614),
.B(n_3937),
.Y(n_7611)
);

NAND2xp5_ASAP7_75t_L g7612 ( 
.A(n_6313),
.B(n_3939),
.Y(n_7612)
);

AND3x2_ASAP7_75t_L g7613 ( 
.A(n_6699),
.B(n_6709),
.C(n_6811),
.Y(n_7613)
);

INVx2_ASAP7_75t_L g7614 ( 
.A(n_6768),
.Y(n_7614)
);

INVx2_ASAP7_75t_L g7615 ( 
.A(n_6776),
.Y(n_7615)
);

AOI22xp33_ASAP7_75t_L g7616 ( 
.A1(n_6324),
.A2(n_3942),
.B1(n_3943),
.B2(n_3940),
.Y(n_7616)
);

INVx1_ASAP7_75t_L g7617 ( 
.A(n_6372),
.Y(n_7617)
);

INVx2_ASAP7_75t_L g7618 ( 
.A(n_6777),
.Y(n_7618)
);

INVx2_ASAP7_75t_L g7619 ( 
.A(n_6783),
.Y(n_7619)
);

INVx1_ASAP7_75t_L g7620 ( 
.A(n_6386),
.Y(n_7620)
);

AND2x2_ASAP7_75t_L g7621 ( 
.A(n_6319),
.B(n_6224),
.Y(n_7621)
);

INVx1_ASAP7_75t_SL g7622 ( 
.A(n_6808),
.Y(n_7622)
);

NOR2x1p5_ASAP7_75t_L g7623 ( 
.A(n_6832),
.B(n_6311),
.Y(n_7623)
);

INVx2_ASAP7_75t_L g7624 ( 
.A(n_6788),
.Y(n_7624)
);

INVx2_ASAP7_75t_SL g7625 ( 
.A(n_6754),
.Y(n_7625)
);

AND2x2_ASAP7_75t_L g7626 ( 
.A(n_6194),
.B(n_3944),
.Y(n_7626)
);

INVx1_ASAP7_75t_L g7627 ( 
.A(n_6389),
.Y(n_7627)
);

INVx2_ASAP7_75t_SL g7628 ( 
.A(n_6754),
.Y(n_7628)
);

INVx2_ASAP7_75t_L g7629 ( 
.A(n_6791),
.Y(n_7629)
);

INVx2_ASAP7_75t_L g7630 ( 
.A(n_6797),
.Y(n_7630)
);

NOR2xp33_ASAP7_75t_L g7631 ( 
.A(n_6745),
.B(n_3946),
.Y(n_7631)
);

NOR2xp33_ASAP7_75t_L g7632 ( 
.A(n_6753),
.B(n_3947),
.Y(n_7632)
);

INVx3_ASAP7_75t_L g7633 ( 
.A(n_6814),
.Y(n_7633)
);

INVx2_ASAP7_75t_L g7634 ( 
.A(n_6813),
.Y(n_7634)
);

INVx1_ASAP7_75t_L g7635 ( 
.A(n_6415),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_6430),
.Y(n_7636)
);

HB1xp67_ASAP7_75t_L g7637 ( 
.A(n_6456),
.Y(n_7637)
);

INVx2_ASAP7_75t_L g7638 ( 
.A(n_6815),
.Y(n_7638)
);

OR2x2_ASAP7_75t_L g7639 ( 
.A(n_6732),
.B(n_3948),
.Y(n_7639)
);

BUFx3_ASAP7_75t_L g7640 ( 
.A(n_6814),
.Y(n_7640)
);

INVx3_ASAP7_75t_L g7641 ( 
.A(n_6829),
.Y(n_7641)
);

INVx1_ASAP7_75t_L g7642 ( 
.A(n_6457),
.Y(n_7642)
);

INVx2_ASAP7_75t_L g7643 ( 
.A(n_6819),
.Y(n_7643)
);

INVx2_ASAP7_75t_L g7644 ( 
.A(n_6822),
.Y(n_7644)
);

INVx2_ASAP7_75t_SL g7645 ( 
.A(n_6829),
.Y(n_7645)
);

NAND2xp5_ASAP7_75t_L g7646 ( 
.A(n_6458),
.B(n_3949),
.Y(n_7646)
);

BUFx6f_ASAP7_75t_SL g7647 ( 
.A(n_6244),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_6459),
.Y(n_7648)
);

INVx1_ASAP7_75t_L g7649 ( 
.A(n_6462),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_6485),
.Y(n_7650)
);

INVx4_ASAP7_75t_L g7651 ( 
.A(n_6843),
.Y(n_7651)
);

BUFx6f_ASAP7_75t_SL g7652 ( 
.A(n_6256),
.Y(n_7652)
);

AOI22xp33_ASAP7_75t_L g7653 ( 
.A1(n_6886),
.A2(n_3952),
.B1(n_3954),
.B2(n_3951),
.Y(n_7653)
);

INVx2_ASAP7_75t_L g7654 ( 
.A(n_6831),
.Y(n_7654)
);

INVx1_ASAP7_75t_L g7655 ( 
.A(n_6513),
.Y(n_7655)
);

INVx2_ASAP7_75t_L g7656 ( 
.A(n_6834),
.Y(n_7656)
);

INVx1_ASAP7_75t_L g7657 ( 
.A(n_6515),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_6531),
.Y(n_7658)
);

INVx1_ASAP7_75t_L g7659 ( 
.A(n_6539),
.Y(n_7659)
);

INVx2_ASAP7_75t_L g7660 ( 
.A(n_6836),
.Y(n_7660)
);

INVx2_ASAP7_75t_L g7661 ( 
.A(n_6838),
.Y(n_7661)
);

NAND2xp5_ASAP7_75t_L g7662 ( 
.A(n_6742),
.B(n_3956),
.Y(n_7662)
);

NAND2xp5_ASAP7_75t_SL g7663 ( 
.A(n_6323),
.B(n_3958),
.Y(n_7663)
);

BUFx4f_ASAP7_75t_L g7664 ( 
.A(n_6226),
.Y(n_7664)
);

INVx2_ASAP7_75t_L g7665 ( 
.A(n_6845),
.Y(n_7665)
);

NAND2xp5_ASAP7_75t_L g7666 ( 
.A(n_6743),
.B(n_3960),
.Y(n_7666)
);

INVx4_ASAP7_75t_L g7667 ( 
.A(n_6843),
.Y(n_7667)
);

NOR2xp33_ASAP7_75t_L g7668 ( 
.A(n_6850),
.B(n_6844),
.Y(n_7668)
);

INVx2_ASAP7_75t_L g7669 ( 
.A(n_6527),
.Y(n_7669)
);

NOR2xp33_ASAP7_75t_L g7670 ( 
.A(n_6765),
.B(n_6767),
.Y(n_7670)
);

INVx2_ASAP7_75t_L g7671 ( 
.A(n_6833),
.Y(n_7671)
);

CKINVDCx5p33_ASAP7_75t_R g7672 ( 
.A(n_6535),
.Y(n_7672)
);

NAND2xp33_ASAP7_75t_SL g7673 ( 
.A(n_6383),
.B(n_3961),
.Y(n_7673)
);

INVxp33_ASAP7_75t_L g7674 ( 
.A(n_6460),
.Y(n_7674)
);

INVx2_ASAP7_75t_L g7675 ( 
.A(n_6840),
.Y(n_7675)
);

AND2x2_ASAP7_75t_L g7676 ( 
.A(n_6784),
.B(n_3963),
.Y(n_7676)
);

AOI22xp33_ASAP7_75t_L g7677 ( 
.A1(n_6897),
.A2(n_3971),
.B1(n_3973),
.B2(n_3970),
.Y(n_7677)
);

INVx3_ASAP7_75t_L g7678 ( 
.A(n_6717),
.Y(n_7678)
);

INVx1_ASAP7_75t_L g7679 ( 
.A(n_6841),
.Y(n_7679)
);

INVx1_ASAP7_75t_L g7680 ( 
.A(n_6846),
.Y(n_7680)
);

BUFx2_ASAP7_75t_L g7681 ( 
.A(n_6498),
.Y(n_7681)
);

NAND2xp5_ASAP7_75t_L g7682 ( 
.A(n_6226),
.B(n_3976),
.Y(n_7682)
);

INVx2_ASAP7_75t_L g7683 ( 
.A(n_6847),
.Y(n_7683)
);

NAND2xp5_ASAP7_75t_L g7684 ( 
.A(n_6287),
.B(n_3978),
.Y(n_7684)
);

BUFx6f_ASAP7_75t_SL g7685 ( 
.A(n_6387),
.Y(n_7685)
);

NOR2xp33_ASAP7_75t_L g7686 ( 
.A(n_6893),
.B(n_3982),
.Y(n_7686)
);

BUFx3_ASAP7_75t_L g7687 ( 
.A(n_6592),
.Y(n_7687)
);

AND2x2_ASAP7_75t_L g7688 ( 
.A(n_6785),
.B(n_3987),
.Y(n_7688)
);

INVx2_ASAP7_75t_L g7689 ( 
.A(n_6719),
.Y(n_7689)
);

NAND2xp5_ASAP7_75t_SL g7690 ( 
.A(n_6331),
.B(n_3993),
.Y(n_7690)
);

INVx1_ASAP7_75t_L g7691 ( 
.A(n_6711),
.Y(n_7691)
);

INVx2_ASAP7_75t_L g7692 ( 
.A(n_6751),
.Y(n_7692)
);

INVx2_ASAP7_75t_SL g7693 ( 
.A(n_6772),
.Y(n_7693)
);

NOR2xp33_ASAP7_75t_L g7694 ( 
.A(n_6789),
.B(n_3994),
.Y(n_7694)
);

INVx2_ASAP7_75t_L g7695 ( 
.A(n_6752),
.Y(n_7695)
);

NAND2xp5_ASAP7_75t_L g7696 ( 
.A(n_6287),
.B(n_3995),
.Y(n_7696)
);

OAI22xp5_ASAP7_75t_L g7697 ( 
.A1(n_6877),
.A2(n_4003),
.B1(n_4004),
.B2(n_4000),
.Y(n_7697)
);

INVxp67_ASAP7_75t_SL g7698 ( 
.A(n_6520),
.Y(n_7698)
);

NAND2xp5_ASAP7_75t_L g7699 ( 
.A(n_6287),
.B(n_4006),
.Y(n_7699)
);

INVx1_ASAP7_75t_L g7700 ( 
.A(n_6793),
.Y(n_7700)
);

INVx1_ASAP7_75t_L g7701 ( 
.A(n_6826),
.Y(n_7701)
);

INVx1_ASAP7_75t_L g7702 ( 
.A(n_6842),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_6848),
.Y(n_7703)
);

OAI22xp5_ASAP7_75t_L g7704 ( 
.A1(n_6564),
.A2(n_4011),
.B1(n_4013),
.B2(n_4007),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_6568),
.Y(n_7705)
);

INVx2_ASAP7_75t_L g7706 ( 
.A(n_6618),
.Y(n_7706)
);

INVx2_ASAP7_75t_L g7707 ( 
.A(n_6685),
.Y(n_7707)
);

INVx2_ASAP7_75t_L g7708 ( 
.A(n_6687),
.Y(n_7708)
);

INVx1_ASAP7_75t_L g7709 ( 
.A(n_6632),
.Y(n_7709)
);

INVx1_ASAP7_75t_L g7710 ( 
.A(n_6689),
.Y(n_7710)
);

AND2x2_ASAP7_75t_L g7711 ( 
.A(n_6792),
.B(n_6910),
.Y(n_7711)
);

INVx2_ASAP7_75t_SL g7712 ( 
.A(n_6706),
.Y(n_7712)
);

INVx2_ASAP7_75t_L g7713 ( 
.A(n_6849),
.Y(n_7713)
);

INVx2_ASAP7_75t_L g7714 ( 
.A(n_6924),
.Y(n_7714)
);

AND2x6_ASAP7_75t_L g7715 ( 
.A(n_6326),
.B(n_6412),
.Y(n_7715)
);

INVx4_ASAP7_75t_L g7716 ( 
.A(n_6397),
.Y(n_7716)
);

INVx2_ASAP7_75t_L g7717 ( 
.A(n_6529),
.Y(n_7717)
);

INVx3_ASAP7_75t_L g7718 ( 
.A(n_6530),
.Y(n_7718)
);

NAND3xp33_ASAP7_75t_L g7719 ( 
.A(n_6588),
.B(n_4018),
.C(n_4016),
.Y(n_7719)
);

INVx2_ASAP7_75t_L g7720 ( 
.A(n_6925),
.Y(n_7720)
);

INVx2_ASAP7_75t_L g7721 ( 
.A(n_6385),
.Y(n_7721)
);

INVx2_ASAP7_75t_SL g7722 ( 
.A(n_6442),
.Y(n_7722)
);

INVx2_ASAP7_75t_L g7723 ( 
.A(n_6554),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_6558),
.Y(n_7724)
);

NAND2xp5_ASAP7_75t_L g7725 ( 
.A(n_6944),
.B(n_4020),
.Y(n_7725)
);

INVx3_ASAP7_75t_L g7726 ( 
.A(n_6469),
.Y(n_7726)
);

AOI22xp33_ASAP7_75t_L g7727 ( 
.A1(n_6939),
.A2(n_4023),
.B1(n_4025),
.B2(n_4022),
.Y(n_7727)
);

NAND2xp5_ASAP7_75t_L g7728 ( 
.A(n_6261),
.B(n_4026),
.Y(n_7728)
);

INVx1_ASAP7_75t_L g7729 ( 
.A(n_6964),
.Y(n_7729)
);

INVxp67_ASAP7_75t_L g7730 ( 
.A(n_7059),
.Y(n_7730)
);

NOR2xp33_ASAP7_75t_L g7731 ( 
.A(n_6966),
.B(n_4029),
.Y(n_7731)
);

AND2x2_ASAP7_75t_SL g7732 ( 
.A(n_7050),
.B(n_3683),
.Y(n_7732)
);

XOR2xp5_ASAP7_75t_L g7733 ( 
.A(n_7209),
.B(n_4030),
.Y(n_7733)
);

CKINVDCx20_ASAP7_75t_R g7734 ( 
.A(n_7270),
.Y(n_7734)
);

BUFx3_ASAP7_75t_L g7735 ( 
.A(n_7114),
.Y(n_7735)
);

AND2x2_ASAP7_75t_L g7736 ( 
.A(n_7053),
.B(n_4035),
.Y(n_7736)
);

CKINVDCx16_ASAP7_75t_R g7737 ( 
.A(n_7299),
.Y(n_7737)
);

BUFx3_ASAP7_75t_L g7738 ( 
.A(n_7114),
.Y(n_7738)
);

INVxp67_ASAP7_75t_L g7739 ( 
.A(n_7011),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_6975),
.Y(n_7740)
);

INVx3_ASAP7_75t_L g7741 ( 
.A(n_6967),
.Y(n_7741)
);

NAND2xp5_ASAP7_75t_SL g7742 ( 
.A(n_7021),
.B(n_7138),
.Y(n_7742)
);

AOI21x1_ASAP7_75t_L g7743 ( 
.A1(n_7545),
.A2(n_7495),
.B(n_7561),
.Y(n_7743)
);

NOR2xp33_ASAP7_75t_L g7744 ( 
.A(n_7004),
.B(n_4037),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_6977),
.Y(n_7745)
);

XOR2xp5_ASAP7_75t_L g7746 ( 
.A(n_7158),
.B(n_7208),
.Y(n_7746)
);

INVx2_ASAP7_75t_SL g7747 ( 
.A(n_7515),
.Y(n_7747)
);

CKINVDCx5p33_ASAP7_75t_R g7748 ( 
.A(n_7065),
.Y(n_7748)
);

INVx1_ASAP7_75t_L g7749 ( 
.A(n_6984),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_6987),
.Y(n_7750)
);

NAND2xp5_ASAP7_75t_L g7751 ( 
.A(n_7670),
.B(n_4039),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_6993),
.Y(n_7752)
);

INVx2_ASAP7_75t_L g7753 ( 
.A(n_7266),
.Y(n_7753)
);

INVx1_ASAP7_75t_L g7754 ( 
.A(n_7008),
.Y(n_7754)
);

INVx1_ASAP7_75t_L g7755 ( 
.A(n_7009),
.Y(n_7755)
);

INVx1_ASAP7_75t_L g7756 ( 
.A(n_7014),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_7048),
.Y(n_7757)
);

NOR2xp33_ASAP7_75t_L g7758 ( 
.A(n_7174),
.B(n_4040),
.Y(n_7758)
);

INVx1_ASAP7_75t_L g7759 ( 
.A(n_7049),
.Y(n_7759)
);

XOR2xp5_ASAP7_75t_L g7760 ( 
.A(n_7332),
.B(n_7396),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_7052),
.Y(n_7761)
);

NOR2xp67_ASAP7_75t_L g7762 ( 
.A(n_6992),
.B(n_4041),
.Y(n_7762)
);

INVxp33_ASAP7_75t_L g7763 ( 
.A(n_7432),
.Y(n_7763)
);

AND2x2_ASAP7_75t_L g7764 ( 
.A(n_7028),
.B(n_7621),
.Y(n_7764)
);

INVx1_ASAP7_75t_L g7765 ( 
.A(n_7054),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_7055),
.Y(n_7766)
);

XNOR2xp5_ASAP7_75t_L g7767 ( 
.A(n_7573),
.B(n_7133),
.Y(n_7767)
);

INVx1_ASAP7_75t_L g7768 ( 
.A(n_7057),
.Y(n_7768)
);

INVx1_ASAP7_75t_L g7769 ( 
.A(n_7058),
.Y(n_7769)
);

INVx1_ASAP7_75t_L g7770 ( 
.A(n_7069),
.Y(n_7770)
);

XNOR2x2_ASAP7_75t_L g7771 ( 
.A(n_7127),
.B(n_3689),
.Y(n_7771)
);

INVx2_ASAP7_75t_L g7772 ( 
.A(n_7269),
.Y(n_7772)
);

CKINVDCx5p33_ASAP7_75t_R g7773 ( 
.A(n_7025),
.Y(n_7773)
);

AND2x2_ASAP7_75t_L g7774 ( 
.A(n_7371),
.B(n_4042),
.Y(n_7774)
);

NOR2xp33_ASAP7_75t_L g7775 ( 
.A(n_7089),
.B(n_4043),
.Y(n_7775)
);

AOI21xp5_ASAP7_75t_L g7776 ( 
.A1(n_7471),
.A2(n_3004),
.B(n_2998),
.Y(n_7776)
);

INVx1_ASAP7_75t_L g7777 ( 
.A(n_7070),
.Y(n_7777)
);

INVx2_ASAP7_75t_L g7778 ( 
.A(n_7271),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_7073),
.Y(n_7779)
);

BUFx6f_ASAP7_75t_L g7780 ( 
.A(n_6965),
.Y(n_7780)
);

INVxp67_ASAP7_75t_L g7781 ( 
.A(n_7218),
.Y(n_7781)
);

INVx1_ASAP7_75t_L g7782 ( 
.A(n_7084),
.Y(n_7782)
);

NOR2xp33_ASAP7_75t_L g7783 ( 
.A(n_7135),
.B(n_4047),
.Y(n_7783)
);

XOR2xp5_ASAP7_75t_L g7784 ( 
.A(n_7111),
.B(n_7408),
.Y(n_7784)
);

INVx1_ASAP7_75t_L g7785 ( 
.A(n_7088),
.Y(n_7785)
);

INVx2_ASAP7_75t_SL g7786 ( 
.A(n_7515),
.Y(n_7786)
);

INVx1_ASAP7_75t_L g7787 ( 
.A(n_7092),
.Y(n_7787)
);

INVx1_ASAP7_75t_L g7788 ( 
.A(n_7094),
.Y(n_7788)
);

INVx2_ASAP7_75t_L g7789 ( 
.A(n_7272),
.Y(n_7789)
);

INVx1_ASAP7_75t_L g7790 ( 
.A(n_7095),
.Y(n_7790)
);

INVx1_ASAP7_75t_L g7791 ( 
.A(n_7098),
.Y(n_7791)
);

AND2x2_ASAP7_75t_L g7792 ( 
.A(n_7108),
.B(n_4051),
.Y(n_7792)
);

NAND2xp5_ASAP7_75t_L g7793 ( 
.A(n_7221),
.B(n_4054),
.Y(n_7793)
);

INVx1_ASAP7_75t_L g7794 ( 
.A(n_7100),
.Y(n_7794)
);

AND2x2_ASAP7_75t_L g7795 ( 
.A(n_7198),
.B(n_3013),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_7113),
.Y(n_7796)
);

INVx1_ASAP7_75t_L g7797 ( 
.A(n_7119),
.Y(n_7797)
);

INVx1_ASAP7_75t_L g7798 ( 
.A(n_7124),
.Y(n_7798)
);

INVx1_ASAP7_75t_L g7799 ( 
.A(n_7125),
.Y(n_7799)
);

NAND2xp5_ASAP7_75t_L g7800 ( 
.A(n_7225),
.B(n_3054),
.Y(n_7800)
);

NOR2xp33_ASAP7_75t_L g7801 ( 
.A(n_7533),
.B(n_3147),
.Y(n_7801)
);

INVx1_ASAP7_75t_L g7802 ( 
.A(n_7126),
.Y(n_7802)
);

AND2x2_ASAP7_75t_L g7803 ( 
.A(n_7493),
.B(n_3326),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_7128),
.Y(n_7804)
);

CKINVDCx5p33_ASAP7_75t_R g7805 ( 
.A(n_7363),
.Y(n_7805)
);

BUFx2_ASAP7_75t_L g7806 ( 
.A(n_7168),
.Y(n_7806)
);

INVx1_ASAP7_75t_L g7807 ( 
.A(n_7129),
.Y(n_7807)
);

INVx2_ASAP7_75t_L g7808 ( 
.A(n_7275),
.Y(n_7808)
);

INVx1_ASAP7_75t_L g7809 ( 
.A(n_7153),
.Y(n_7809)
);

AND2x2_ASAP7_75t_L g7810 ( 
.A(n_6968),
.B(n_3448),
.Y(n_7810)
);

NOR2xp33_ASAP7_75t_SL g7811 ( 
.A(n_6956),
.B(n_7016),
.Y(n_7811)
);

INVx1_ASAP7_75t_L g7812 ( 
.A(n_7156),
.Y(n_7812)
);

INVx1_ASAP7_75t_L g7813 ( 
.A(n_7162),
.Y(n_7813)
);

INVx1_ASAP7_75t_L g7814 ( 
.A(n_7163),
.Y(n_7814)
);

INVx1_ASAP7_75t_L g7815 ( 
.A(n_7166),
.Y(n_7815)
);

OAI21xp5_ASAP7_75t_L g7816 ( 
.A1(n_7575),
.A2(n_3485),
.B(n_3449),
.Y(n_7816)
);

CKINVDCx20_ASAP7_75t_R g7817 ( 
.A(n_7409),
.Y(n_7817)
);

INVx1_ASAP7_75t_L g7818 ( 
.A(n_7169),
.Y(n_7818)
);

INVx2_ASAP7_75t_L g7819 ( 
.A(n_7279),
.Y(n_7819)
);

CKINVDCx20_ASAP7_75t_R g7820 ( 
.A(n_7118),
.Y(n_7820)
);

INVx2_ASAP7_75t_SL g7821 ( 
.A(n_7556),
.Y(n_7821)
);

AND2x2_ASAP7_75t_L g7822 ( 
.A(n_7446),
.B(n_6973),
.Y(n_7822)
);

NOR2xp33_ASAP7_75t_SL g7823 ( 
.A(n_7137),
.B(n_3692),
.Y(n_7823)
);

BUFx5_ASAP7_75t_L g7824 ( 
.A(n_7389),
.Y(n_7824)
);

INVx1_ASAP7_75t_L g7825 ( 
.A(n_7179),
.Y(n_7825)
);

INVx2_ASAP7_75t_L g7826 ( 
.A(n_7282),
.Y(n_7826)
);

INVx1_ASAP7_75t_L g7827 ( 
.A(n_7180),
.Y(n_7827)
);

XOR2xp5_ASAP7_75t_L g7828 ( 
.A(n_7508),
.B(n_3701),
.Y(n_7828)
);

AND2x2_ASAP7_75t_L g7829 ( 
.A(n_7260),
.B(n_7711),
.Y(n_7829)
);

BUFx5_ASAP7_75t_L g7830 ( 
.A(n_7389),
.Y(n_7830)
);

AND2x2_ASAP7_75t_SL g7831 ( 
.A(n_7664),
.B(n_3710),
.Y(n_7831)
);

NAND2x1p5_ASAP7_75t_L g7832 ( 
.A(n_7556),
.B(n_3719),
.Y(n_7832)
);

INVx1_ASAP7_75t_L g7833 ( 
.A(n_7183),
.Y(n_7833)
);

INVx2_ASAP7_75t_SL g7834 ( 
.A(n_6989),
.Y(n_7834)
);

INVx1_ASAP7_75t_L g7835 ( 
.A(n_7189),
.Y(n_7835)
);

INVx1_ASAP7_75t_L g7836 ( 
.A(n_7192),
.Y(n_7836)
);

INVx1_ASAP7_75t_L g7837 ( 
.A(n_7195),
.Y(n_7837)
);

INVxp67_ASAP7_75t_SL g7838 ( 
.A(n_7248),
.Y(n_7838)
);

NOR2xp33_ASAP7_75t_L g7839 ( 
.A(n_7388),
.B(n_3522),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7199),
.Y(n_7840)
);

AND2x6_ASAP7_75t_L g7841 ( 
.A(n_7726),
.B(n_7447),
.Y(n_7841)
);

NAND2xp5_ASAP7_75t_SL g7842 ( 
.A(n_7604),
.B(n_3735),
.Y(n_7842)
);

AND2x2_ASAP7_75t_L g7843 ( 
.A(n_6981),
.B(n_3804),
.Y(n_7843)
);

INVx2_ASAP7_75t_L g7844 ( 
.A(n_7285),
.Y(n_7844)
);

INVx1_ASAP7_75t_L g7845 ( 
.A(n_7203),
.Y(n_7845)
);

NAND2x1p5_ASAP7_75t_L g7846 ( 
.A(n_7268),
.B(n_3725),
.Y(n_7846)
);

INVx1_ASAP7_75t_L g7847 ( 
.A(n_7206),
.Y(n_7847)
);

INVx2_ASAP7_75t_L g7848 ( 
.A(n_7287),
.Y(n_7848)
);

INVx1_ASAP7_75t_L g7849 ( 
.A(n_7210),
.Y(n_7849)
);

INVx1_ASAP7_75t_L g7850 ( 
.A(n_7212),
.Y(n_7850)
);

CKINVDCx20_ASAP7_75t_R g7851 ( 
.A(n_7229),
.Y(n_7851)
);

INVx1_ASAP7_75t_L g7852 ( 
.A(n_7220),
.Y(n_7852)
);

AND2x2_ASAP7_75t_L g7853 ( 
.A(n_7353),
.B(n_3822),
.Y(n_7853)
);

INVx1_ASAP7_75t_L g7854 ( 
.A(n_7223),
.Y(n_7854)
);

INVx2_ASAP7_75t_L g7855 ( 
.A(n_7290),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_7231),
.Y(n_7856)
);

INVx1_ASAP7_75t_L g7857 ( 
.A(n_7237),
.Y(n_7857)
);

INVx1_ASAP7_75t_L g7858 ( 
.A(n_7240),
.Y(n_7858)
);

CKINVDCx16_ASAP7_75t_R g7859 ( 
.A(n_6989),
.Y(n_7859)
);

AOI21x1_ASAP7_75t_L g7860 ( 
.A1(n_7563),
.A2(n_3729),
.B(n_3726),
.Y(n_7860)
);

AND2x2_ASAP7_75t_L g7861 ( 
.A(n_7577),
.B(n_3957),
.Y(n_7861)
);

INVx1_ASAP7_75t_L g7862 ( 
.A(n_7243),
.Y(n_7862)
);

CKINVDCx20_ASAP7_75t_R g7863 ( 
.A(n_6985),
.Y(n_7863)
);

INVx1_ASAP7_75t_L g7864 ( 
.A(n_7247),
.Y(n_7864)
);

INVx2_ASAP7_75t_L g7865 ( 
.A(n_7298),
.Y(n_7865)
);

XNOR2xp5_ASAP7_75t_L g7866 ( 
.A(n_7472),
.B(n_3730),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_7253),
.Y(n_7867)
);

INVx1_ASAP7_75t_L g7868 ( 
.A(n_7256),
.Y(n_7868)
);

INVx1_ASAP7_75t_L g7869 ( 
.A(n_7263),
.Y(n_7869)
);

AND2x2_ASAP7_75t_L g7870 ( 
.A(n_7585),
.B(n_3974),
.Y(n_7870)
);

BUFx6f_ASAP7_75t_L g7871 ( 
.A(n_6965),
.Y(n_7871)
);

INVxp67_ASAP7_75t_SL g7872 ( 
.A(n_7465),
.Y(n_7872)
);

AND2x2_ASAP7_75t_L g7873 ( 
.A(n_7587),
.B(n_3991),
.Y(n_7873)
);

NOR2xp33_ASAP7_75t_L g7874 ( 
.A(n_7428),
.B(n_7394),
.Y(n_7874)
);

INVx1_ASAP7_75t_L g7875 ( 
.A(n_7284),
.Y(n_7875)
);

INVxp33_ASAP7_75t_L g7876 ( 
.A(n_7312),
.Y(n_7876)
);

INVx1_ASAP7_75t_L g7877 ( 
.A(n_7289),
.Y(n_7877)
);

AOI21xp5_ASAP7_75t_L g7878 ( 
.A1(n_7274),
.A2(n_4049),
.B(n_3743),
.Y(n_7878)
);

CKINVDCx5p33_ASAP7_75t_R g7879 ( 
.A(n_7131),
.Y(n_7879)
);

INVx2_ASAP7_75t_L g7880 ( 
.A(n_7305),
.Y(n_7880)
);

INVx1_ASAP7_75t_L g7881 ( 
.A(n_7302),
.Y(n_7881)
);

BUFx6f_ASAP7_75t_SL g7882 ( 
.A(n_7368),
.Y(n_7882)
);

INVx1_ASAP7_75t_L g7883 ( 
.A(n_7303),
.Y(n_7883)
);

INVx2_ASAP7_75t_SL g7884 ( 
.A(n_7268),
.Y(n_7884)
);

CKINVDCx5p33_ASAP7_75t_R g7885 ( 
.A(n_7376),
.Y(n_7885)
);

NOR2xp33_ASAP7_75t_L g7886 ( 
.A(n_7411),
.B(n_3732),
.Y(n_7886)
);

INVx1_ASAP7_75t_L g7887 ( 
.A(n_7304),
.Y(n_7887)
);

INVx1_ASAP7_75t_L g7888 ( 
.A(n_7308),
.Y(n_7888)
);

INVx1_ASAP7_75t_L g7889 ( 
.A(n_7310),
.Y(n_7889)
);

INVx1_ASAP7_75t_L g7890 ( 
.A(n_7313),
.Y(n_7890)
);

INVx1_ASAP7_75t_L g7891 ( 
.A(n_7317),
.Y(n_7891)
);

AND2x2_ASAP7_75t_L g7892 ( 
.A(n_7595),
.B(n_3749),
.Y(n_7892)
);

INVx1_ASAP7_75t_L g7893 ( 
.A(n_7321),
.Y(n_7893)
);

INVx1_ASAP7_75t_L g7894 ( 
.A(n_7324),
.Y(n_7894)
);

INVx1_ASAP7_75t_L g7895 ( 
.A(n_7325),
.Y(n_7895)
);

NAND2xp33_ASAP7_75t_R g7896 ( 
.A(n_7205),
.B(n_4),
.Y(n_7896)
);

AND2x2_ASAP7_75t_L g7897 ( 
.A(n_7369),
.B(n_3760),
.Y(n_7897)
);

NOR2xp67_ASAP7_75t_L g7898 ( 
.A(n_7261),
.B(n_5),
.Y(n_7898)
);

INVx1_ASAP7_75t_L g7899 ( 
.A(n_7329),
.Y(n_7899)
);

INVx1_ASAP7_75t_L g7900 ( 
.A(n_7330),
.Y(n_7900)
);

INVx1_ASAP7_75t_L g7901 ( 
.A(n_7335),
.Y(n_7901)
);

INVx1_ASAP7_75t_L g7902 ( 
.A(n_7336),
.Y(n_7902)
);

NOR2xp33_ASAP7_75t_L g7903 ( 
.A(n_7674),
.B(n_3765),
.Y(n_7903)
);

XNOR2x2_ASAP7_75t_L g7904 ( 
.A(n_6998),
.B(n_3767),
.Y(n_7904)
);

CKINVDCx16_ASAP7_75t_R g7905 ( 
.A(n_7445),
.Y(n_7905)
);

INVx1_ASAP7_75t_L g7906 ( 
.A(n_7337),
.Y(n_7906)
);

INVx1_ASAP7_75t_L g7907 ( 
.A(n_7339),
.Y(n_7907)
);

NAND2xp5_ASAP7_75t_SL g7908 ( 
.A(n_7190),
.B(n_3261),
.Y(n_7908)
);

NAND2x1p5_ASAP7_75t_L g7909 ( 
.A(n_7355),
.B(n_3769),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_7343),
.Y(n_7910)
);

INVx1_ASAP7_75t_L g7911 ( 
.A(n_7356),
.Y(n_7911)
);

AND2x4_ASAP7_75t_L g7912 ( 
.A(n_6958),
.B(n_3771),
.Y(n_7912)
);

INVx1_ASAP7_75t_L g7913 ( 
.A(n_7359),
.Y(n_7913)
);

NOR2xp33_ASAP7_75t_L g7914 ( 
.A(n_7291),
.B(n_3786),
.Y(n_7914)
);

INVx1_ASAP7_75t_L g7915 ( 
.A(n_7361),
.Y(n_7915)
);

XOR2xp5_ASAP7_75t_L g7916 ( 
.A(n_7590),
.B(n_3787),
.Y(n_7916)
);

AND2x2_ASAP7_75t_L g7917 ( 
.A(n_7698),
.B(n_3791),
.Y(n_7917)
);

INVxp33_ASAP7_75t_SL g7918 ( 
.A(n_7672),
.Y(n_7918)
);

INVx1_ASAP7_75t_L g7919 ( 
.A(n_7364),
.Y(n_7919)
);

INVx1_ASAP7_75t_L g7920 ( 
.A(n_7382),
.Y(n_7920)
);

CKINVDCx5p33_ASAP7_75t_R g7921 ( 
.A(n_7477),
.Y(n_7921)
);

INVx1_ASAP7_75t_L g7922 ( 
.A(n_7383),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_7386),
.Y(n_7923)
);

INVx1_ASAP7_75t_L g7924 ( 
.A(n_7391),
.Y(n_7924)
);

NOR2xp33_ASAP7_75t_L g7925 ( 
.A(n_7309),
.B(n_3794),
.Y(n_7925)
);

INVx1_ASAP7_75t_L g7926 ( 
.A(n_7393),
.Y(n_7926)
);

INVx1_ASAP7_75t_L g7927 ( 
.A(n_7395),
.Y(n_7927)
);

BUFx6f_ASAP7_75t_L g7928 ( 
.A(n_6990),
.Y(n_7928)
);

NOR2xp33_ASAP7_75t_L g7929 ( 
.A(n_7230),
.B(n_3796),
.Y(n_7929)
);

CKINVDCx20_ASAP7_75t_R g7930 ( 
.A(n_6996),
.Y(n_7930)
);

AND2x2_ASAP7_75t_L g7931 ( 
.A(n_7626),
.B(n_3799),
.Y(n_7931)
);

NOR2xp33_ASAP7_75t_L g7932 ( 
.A(n_7236),
.B(n_3814),
.Y(n_7932)
);

INVx1_ASAP7_75t_L g7933 ( 
.A(n_7398),
.Y(n_7933)
);

INVx1_ASAP7_75t_L g7934 ( 
.A(n_7399),
.Y(n_7934)
);

AND2x2_ASAP7_75t_L g7935 ( 
.A(n_7322),
.B(n_3818),
.Y(n_7935)
);

XNOR2xp5_ASAP7_75t_L g7936 ( 
.A(n_7501),
.B(n_3820),
.Y(n_7936)
);

INVx1_ASAP7_75t_L g7937 ( 
.A(n_7403),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_7404),
.Y(n_7938)
);

AND2x4_ASAP7_75t_L g7939 ( 
.A(n_6969),
.B(n_3823),
.Y(n_7939)
);

INVx2_ASAP7_75t_L g7940 ( 
.A(n_7306),
.Y(n_7940)
);

XOR2xp5_ASAP7_75t_L g7941 ( 
.A(n_7311),
.B(n_3835),
.Y(n_7941)
);

AND2x2_ASAP7_75t_L g7942 ( 
.A(n_7705),
.B(n_3843),
.Y(n_7942)
);

INVx1_ASAP7_75t_L g7943 ( 
.A(n_7435),
.Y(n_7943)
);

NOR2xp33_ASAP7_75t_L g7944 ( 
.A(n_7579),
.B(n_3846),
.Y(n_7944)
);

INVx1_ASAP7_75t_L g7945 ( 
.A(n_7438),
.Y(n_7945)
);

NAND2x1p5_ASAP7_75t_L g7946 ( 
.A(n_7355),
.B(n_3848),
.Y(n_7946)
);

INVx1_ASAP7_75t_L g7947 ( 
.A(n_7440),
.Y(n_7947)
);

NAND2xp5_ASAP7_75t_L g7948 ( 
.A(n_7728),
.B(n_3860),
.Y(n_7948)
);

NAND2xp5_ASAP7_75t_L g7949 ( 
.A(n_6994),
.B(n_3862),
.Y(n_7949)
);

INVx2_ASAP7_75t_L g7950 ( 
.A(n_7307),
.Y(n_7950)
);

AND2x4_ASAP7_75t_L g7951 ( 
.A(n_7015),
.B(n_3867),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_7448),
.Y(n_7952)
);

INVx1_ASAP7_75t_L g7953 ( 
.A(n_7449),
.Y(n_7953)
);

CKINVDCx20_ASAP7_75t_R g7954 ( 
.A(n_6996),
.Y(n_7954)
);

INVx2_ASAP7_75t_L g7955 ( 
.A(n_7320),
.Y(n_7955)
);

NAND2xp5_ASAP7_75t_SL g7956 ( 
.A(n_7316),
.B(n_3871),
.Y(n_7956)
);

AND2x2_ASAP7_75t_L g7957 ( 
.A(n_7709),
.B(n_7676),
.Y(n_7957)
);

INVx1_ASAP7_75t_L g7958 ( 
.A(n_7451),
.Y(n_7958)
);

INVx2_ASAP7_75t_SL g7959 ( 
.A(n_7410),
.Y(n_7959)
);

INVx1_ASAP7_75t_L g7960 ( 
.A(n_7463),
.Y(n_7960)
);

INVx1_ASAP7_75t_L g7961 ( 
.A(n_7466),
.Y(n_7961)
);

INVx1_ASAP7_75t_L g7962 ( 
.A(n_7720),
.Y(n_7962)
);

NOR2xp33_ASAP7_75t_L g7963 ( 
.A(n_7594),
.B(n_3874),
.Y(n_7963)
);

NOR2xp33_ASAP7_75t_L g7964 ( 
.A(n_7599),
.B(n_3879),
.Y(n_7964)
);

AND2x2_ASAP7_75t_L g7965 ( 
.A(n_7688),
.B(n_3880),
.Y(n_7965)
);

AND2x2_ASAP7_75t_L g7966 ( 
.A(n_7557),
.B(n_3881),
.Y(n_7966)
);

NAND2xp5_ASAP7_75t_L g7967 ( 
.A(n_6970),
.B(n_3891),
.Y(n_7967)
);

INVx1_ASAP7_75t_L g7968 ( 
.A(n_7450),
.Y(n_7968)
);

AND2x2_ASAP7_75t_L g7969 ( 
.A(n_7562),
.B(n_3897),
.Y(n_7969)
);

NAND2xp5_ASAP7_75t_L g7970 ( 
.A(n_7622),
.B(n_7035),
.Y(n_7970)
);

INVx2_ASAP7_75t_L g7971 ( 
.A(n_7327),
.Y(n_7971)
);

XOR2xp5_ASAP7_75t_L g7972 ( 
.A(n_6990),
.B(n_3899),
.Y(n_7972)
);

NAND2xp5_ASAP7_75t_L g7973 ( 
.A(n_7694),
.B(n_3900),
.Y(n_7973)
);

BUFx6f_ASAP7_75t_L g7974 ( 
.A(n_7001),
.Y(n_7974)
);

INVxp33_ASAP7_75t_SL g7975 ( 
.A(n_7397),
.Y(n_7975)
);

XOR2xp5_ASAP7_75t_L g7976 ( 
.A(n_7534),
.B(n_3901),
.Y(n_7976)
);

BUFx8_ASAP7_75t_L g7977 ( 
.A(n_7519),
.Y(n_7977)
);

INVx1_ASAP7_75t_L g7978 ( 
.A(n_7338),
.Y(n_7978)
);

INVx1_ASAP7_75t_L g7979 ( 
.A(n_7340),
.Y(n_7979)
);

OR2x2_ASAP7_75t_L g7980 ( 
.A(n_7018),
.B(n_7564),
.Y(n_7980)
);

NAND2xp5_ASAP7_75t_L g7981 ( 
.A(n_7605),
.B(n_3904),
.Y(n_7981)
);

INVx1_ASAP7_75t_L g7982 ( 
.A(n_7342),
.Y(n_7982)
);

NAND2xp5_ASAP7_75t_SL g7983 ( 
.A(n_7319),
.B(n_3911),
.Y(n_7983)
);

INVx1_ASAP7_75t_L g7984 ( 
.A(n_7347),
.Y(n_7984)
);

NOR2xp33_ASAP7_75t_L g7985 ( 
.A(n_7607),
.B(n_3915),
.Y(n_7985)
);

BUFx6f_ASAP7_75t_L g7986 ( 
.A(n_7001),
.Y(n_7986)
);

INVx1_ASAP7_75t_L g7987 ( 
.A(n_7349),
.Y(n_7987)
);

INVxp33_ASAP7_75t_L g7988 ( 
.A(n_7242),
.Y(n_7988)
);

AND2x4_ASAP7_75t_L g7989 ( 
.A(n_7226),
.B(n_3920),
.Y(n_7989)
);

NOR2xp33_ASAP7_75t_L g7990 ( 
.A(n_7608),
.B(n_3923),
.Y(n_7990)
);

INVx1_ASAP7_75t_L g7991 ( 
.A(n_7351),
.Y(n_7991)
);

NOR2xp33_ASAP7_75t_SL g7992 ( 
.A(n_6983),
.B(n_7023),
.Y(n_7992)
);

AND2x2_ASAP7_75t_L g7993 ( 
.A(n_7372),
.B(n_3929),
.Y(n_7993)
);

AND2x2_ASAP7_75t_L g7994 ( 
.A(n_7418),
.B(n_3930),
.Y(n_7994)
);

INVx1_ASAP7_75t_L g7995 ( 
.A(n_7357),
.Y(n_7995)
);

INVx1_ASAP7_75t_L g7996 ( 
.A(n_7366),
.Y(n_7996)
);

INVxp33_ASAP7_75t_L g7997 ( 
.A(n_7637),
.Y(n_7997)
);

INVx2_ASAP7_75t_L g7998 ( 
.A(n_7373),
.Y(n_7998)
);

BUFx3_ASAP7_75t_L g7999 ( 
.A(n_7045),
.Y(n_7999)
);

INVxp67_ASAP7_75t_SL g8000 ( 
.A(n_6961),
.Y(n_8000)
);

XOR2xp5_ASAP7_75t_L g8001 ( 
.A(n_7006),
.B(n_3933),
.Y(n_8001)
);

CKINVDCx20_ASAP7_75t_R g8002 ( 
.A(n_7023),
.Y(n_8002)
);

AND2x2_ASAP7_75t_L g8003 ( 
.A(n_7462),
.B(n_3935),
.Y(n_8003)
);

NOR2xp33_ASAP7_75t_L g8004 ( 
.A(n_7617),
.B(n_3950),
.Y(n_8004)
);

XOR2xp5_ASAP7_75t_L g8005 ( 
.A(n_7106),
.B(n_3953),
.Y(n_8005)
);

INVx1_ASAP7_75t_L g8006 ( 
.A(n_7374),
.Y(n_8006)
);

AOI21xp5_ASAP7_75t_L g8007 ( 
.A1(n_7620),
.A2(n_3962),
.B(n_3959),
.Y(n_8007)
);

INVx1_ASAP7_75t_L g8008 ( 
.A(n_7380),
.Y(n_8008)
);

NOR2x1_ASAP7_75t_L g8009 ( 
.A(n_7420),
.B(n_3967),
.Y(n_8009)
);

INVx1_ASAP7_75t_L g8010 ( 
.A(n_7381),
.Y(n_8010)
);

INVx2_ASAP7_75t_L g8011 ( 
.A(n_7384),
.Y(n_8011)
);

XOR2xp5_ASAP7_75t_L g8012 ( 
.A(n_7122),
.B(n_3969),
.Y(n_8012)
);

AND2x4_ASAP7_75t_L g8013 ( 
.A(n_7716),
.B(n_3984),
.Y(n_8013)
);

AND2x2_ASAP7_75t_L g8014 ( 
.A(n_7481),
.B(n_3985),
.Y(n_8014)
);

INVx2_ASAP7_75t_L g8015 ( 
.A(n_7392),
.Y(n_8015)
);

INVx2_ASAP7_75t_L g8016 ( 
.A(n_7405),
.Y(n_8016)
);

INVx1_ASAP7_75t_L g8017 ( 
.A(n_7406),
.Y(n_8017)
);

INVx1_ASAP7_75t_L g8018 ( 
.A(n_7407),
.Y(n_8018)
);

INVxp67_ASAP7_75t_L g8019 ( 
.A(n_7348),
.Y(n_8019)
);

AND2x4_ASAP7_75t_L g8020 ( 
.A(n_7281),
.B(n_3986),
.Y(n_8020)
);

INVx1_ASAP7_75t_L g8021 ( 
.A(n_7415),
.Y(n_8021)
);

INVx1_ASAP7_75t_L g8022 ( 
.A(n_7419),
.Y(n_8022)
);

INVx1_ASAP7_75t_L g8023 ( 
.A(n_7423),
.Y(n_8023)
);

NOR2xp67_ASAP7_75t_L g8024 ( 
.A(n_7227),
.B(n_5),
.Y(n_8024)
);

INVx1_ASAP7_75t_L g8025 ( 
.A(n_7426),
.Y(n_8025)
);

CKINVDCx20_ASAP7_75t_R g8026 ( 
.A(n_7213),
.Y(n_8026)
);

XOR2xp5_ASAP7_75t_L g8027 ( 
.A(n_7007),
.B(n_3988),
.Y(n_8027)
);

INVx1_ASAP7_75t_L g8028 ( 
.A(n_6952),
.Y(n_8028)
);

INVx1_ASAP7_75t_L g8029 ( 
.A(n_6955),
.Y(n_8029)
);

CKINVDCx5p33_ASAP7_75t_R g8030 ( 
.A(n_7578),
.Y(n_8030)
);

INVx1_ASAP7_75t_L g8031 ( 
.A(n_6957),
.Y(n_8031)
);

NAND2xp5_ASAP7_75t_L g8032 ( 
.A(n_7627),
.B(n_3990),
.Y(n_8032)
);

XNOR2xp5_ASAP7_75t_L g8033 ( 
.A(n_7051),
.B(n_3992),
.Y(n_8033)
);

BUFx3_ASAP7_75t_L g8034 ( 
.A(n_7005),
.Y(n_8034)
);

INVx1_ASAP7_75t_L g8035 ( 
.A(n_6960),
.Y(n_8035)
);

AND2x2_ASAP7_75t_L g8036 ( 
.A(n_7033),
.B(n_7040),
.Y(n_8036)
);

INVx2_ASAP7_75t_L g8037 ( 
.A(n_6962),
.Y(n_8037)
);

NOR2xp33_ASAP7_75t_L g8038 ( 
.A(n_7635),
.B(n_4005),
.Y(n_8038)
);

INVxp33_ASAP7_75t_L g8039 ( 
.A(n_7681),
.Y(n_8039)
);

INVx1_ASAP7_75t_SL g8040 ( 
.A(n_7565),
.Y(n_8040)
);

AND2x2_ASAP7_75t_L g8041 ( 
.A(n_7043),
.B(n_4014),
.Y(n_8041)
);

XNOR2x2_ASAP7_75t_L g8042 ( 
.A(n_7165),
.B(n_4021),
.Y(n_8042)
);

INVx1_ASAP7_75t_L g8043 ( 
.A(n_6971),
.Y(n_8043)
);

INVx1_ASAP7_75t_L g8044 ( 
.A(n_6978),
.Y(n_8044)
);

INVx1_ASAP7_75t_L g8045 ( 
.A(n_6979),
.Y(n_8045)
);

INVxp67_ASAP7_75t_SL g8046 ( 
.A(n_7315),
.Y(n_8046)
);

INVx1_ASAP7_75t_L g8047 ( 
.A(n_6980),
.Y(n_8047)
);

INVxp33_ASAP7_75t_L g8048 ( 
.A(n_7494),
.Y(n_8048)
);

AND2x4_ASAP7_75t_L g8049 ( 
.A(n_7468),
.B(n_4024),
.Y(n_8049)
);

AND2x2_ASAP7_75t_L g8050 ( 
.A(n_7112),
.B(n_5),
.Y(n_8050)
);

CKINVDCx5p33_ASAP7_75t_R g8051 ( 
.A(n_7213),
.Y(n_8051)
);

XOR2xp5_ASAP7_75t_L g8052 ( 
.A(n_7120),
.B(n_6),
.Y(n_8052)
);

BUFx2_ASAP7_75t_L g8053 ( 
.A(n_7715),
.Y(n_8053)
);

BUFx6f_ASAP7_75t_L g8054 ( 
.A(n_7005),
.Y(n_8054)
);

INVx1_ASAP7_75t_L g8055 ( 
.A(n_6982),
.Y(n_8055)
);

INVx2_ASAP7_75t_L g8056 ( 
.A(n_6988),
.Y(n_8056)
);

NOR2xp33_ASAP7_75t_L g8057 ( 
.A(n_7636),
.B(n_2453),
.Y(n_8057)
);

AND2x4_ASAP7_75t_L g8058 ( 
.A(n_7520),
.B(n_6),
.Y(n_8058)
);

INVx2_ASAP7_75t_L g8059 ( 
.A(n_6995),
.Y(n_8059)
);

INVx1_ASAP7_75t_L g8060 ( 
.A(n_6997),
.Y(n_8060)
);

INVxp67_ASAP7_75t_L g8061 ( 
.A(n_7421),
.Y(n_8061)
);

NOR2xp33_ASAP7_75t_L g8062 ( 
.A(n_7642),
.B(n_2453),
.Y(n_8062)
);

INVx2_ASAP7_75t_SL g8063 ( 
.A(n_7410),
.Y(n_8063)
);

OR2x2_ASAP7_75t_L g8064 ( 
.A(n_7080),
.B(n_7117),
.Y(n_8064)
);

NAND2xp5_ASAP7_75t_L g8065 ( 
.A(n_7648),
.B(n_6),
.Y(n_8065)
);

INVx4_ASAP7_75t_L g8066 ( 
.A(n_7460),
.Y(n_8066)
);

INVx1_ASAP7_75t_L g8067 ( 
.A(n_7002),
.Y(n_8067)
);

INVx2_ASAP7_75t_L g8068 ( 
.A(n_7013),
.Y(n_8068)
);

BUFx5_ASAP7_75t_L g8069 ( 
.A(n_7389),
.Y(n_8069)
);

XOR2xp5_ASAP7_75t_L g8070 ( 
.A(n_7024),
.B(n_7),
.Y(n_8070)
);

INVx1_ASAP7_75t_L g8071 ( 
.A(n_7020),
.Y(n_8071)
);

CKINVDCx20_ASAP7_75t_R g8072 ( 
.A(n_7460),
.Y(n_8072)
);

NOR2xp33_ASAP7_75t_L g8073 ( 
.A(n_7649),
.B(n_2454),
.Y(n_8073)
);

INVx1_ASAP7_75t_L g8074 ( 
.A(n_7026),
.Y(n_8074)
);

AND2x2_ASAP7_75t_L g8075 ( 
.A(n_7139),
.B(n_7),
.Y(n_8075)
);

INVx2_ASAP7_75t_L g8076 ( 
.A(n_7029),
.Y(n_8076)
);

INVx1_ASAP7_75t_L g8077 ( 
.A(n_7032),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_7036),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_7038),
.Y(n_8079)
);

BUFx3_ASAP7_75t_L g8080 ( 
.A(n_7024),
.Y(n_8080)
);

INVx1_ASAP7_75t_L g8081 ( 
.A(n_7041),
.Y(n_8081)
);

BUFx2_ASAP7_75t_L g8082 ( 
.A(n_7715),
.Y(n_8082)
);

INVx1_ASAP7_75t_L g8083 ( 
.A(n_7042),
.Y(n_8083)
);

CKINVDCx20_ASAP7_75t_R g8084 ( 
.A(n_7193),
.Y(n_8084)
);

INVx1_ASAP7_75t_L g8085 ( 
.A(n_7047),
.Y(n_8085)
);

INVx1_ASAP7_75t_L g8086 ( 
.A(n_7062),
.Y(n_8086)
);

INVx1_ASAP7_75t_L g8087 ( 
.A(n_7066),
.Y(n_8087)
);

INVx1_ASAP7_75t_L g8088 ( 
.A(n_7076),
.Y(n_8088)
);

OAI21xp5_ASAP7_75t_L g8089 ( 
.A1(n_7650),
.A2(n_7259),
.B(n_7333),
.Y(n_8089)
);

AND2x2_ASAP7_75t_L g8090 ( 
.A(n_7502),
.B(n_7),
.Y(n_8090)
);

CKINVDCx20_ASAP7_75t_R g8091 ( 
.A(n_7219),
.Y(n_8091)
);

INVx1_ASAP7_75t_L g8092 ( 
.A(n_7079),
.Y(n_8092)
);

AND2x2_ASAP7_75t_L g8093 ( 
.A(n_7154),
.B(n_7714),
.Y(n_8093)
);

INVx1_ASAP7_75t_L g8094 ( 
.A(n_7081),
.Y(n_8094)
);

INVx1_ASAP7_75t_L g8095 ( 
.A(n_7082),
.Y(n_8095)
);

INVx1_ASAP7_75t_L g8096 ( 
.A(n_7083),
.Y(n_8096)
);

XNOR2xp5_ASAP7_75t_L g8097 ( 
.A(n_7514),
.B(n_8),
.Y(n_8097)
);

NOR2xp33_ASAP7_75t_SL g8098 ( 
.A(n_6986),
.B(n_8),
.Y(n_8098)
);

INVx1_ASAP7_75t_L g8099 ( 
.A(n_7091),
.Y(n_8099)
);

NAND2xp5_ASAP7_75t_L g8100 ( 
.A(n_7039),
.B(n_8),
.Y(n_8100)
);

INVx1_ASAP7_75t_L g8101 ( 
.A(n_7093),
.Y(n_8101)
);

CKINVDCx5p33_ASAP7_75t_R g8102 ( 
.A(n_7233),
.Y(n_8102)
);

INVx1_ASAP7_75t_L g8103 ( 
.A(n_7103),
.Y(n_8103)
);

INVx1_ASAP7_75t_L g8104 ( 
.A(n_7105),
.Y(n_8104)
);

INVx2_ASAP7_75t_L g8105 ( 
.A(n_7110),
.Y(n_8105)
);

INVx1_ASAP7_75t_L g8106 ( 
.A(n_7116),
.Y(n_8106)
);

CKINVDCx20_ASAP7_75t_R g8107 ( 
.A(n_7207),
.Y(n_8107)
);

INVx1_ASAP7_75t_L g8108 ( 
.A(n_7123),
.Y(n_8108)
);

INVx1_ASAP7_75t_L g8109 ( 
.A(n_7132),
.Y(n_8109)
);

INVx1_ASAP7_75t_L g8110 ( 
.A(n_7141),
.Y(n_8110)
);

INVx2_ASAP7_75t_L g8111 ( 
.A(n_7142),
.Y(n_8111)
);

XNOR2xp5_ASAP7_75t_L g8112 ( 
.A(n_7012),
.B(n_9),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_7145),
.Y(n_8113)
);

INVx2_ASAP7_75t_SL g8114 ( 
.A(n_7554),
.Y(n_8114)
);

INVxp33_ASAP7_75t_L g8115 ( 
.A(n_7314),
.Y(n_8115)
);

INVx1_ASAP7_75t_L g8116 ( 
.A(n_7146),
.Y(n_8116)
);

INVx1_ASAP7_75t_L g8117 ( 
.A(n_7148),
.Y(n_8117)
);

INVx1_ASAP7_75t_L g8118 ( 
.A(n_7151),
.Y(n_8118)
);

INVx2_ASAP7_75t_SL g8119 ( 
.A(n_7554),
.Y(n_8119)
);

INVx1_ASAP7_75t_L g8120 ( 
.A(n_7152),
.Y(n_8120)
);

INVx1_ASAP7_75t_L g8121 ( 
.A(n_7159),
.Y(n_8121)
);

INVx2_ASAP7_75t_SL g8122 ( 
.A(n_7090),
.Y(n_8122)
);

INVx1_ASAP7_75t_L g8123 ( 
.A(n_7161),
.Y(n_8123)
);

INVx4_ASAP7_75t_SL g8124 ( 
.A(n_7715),
.Y(n_8124)
);

INVx1_ASAP7_75t_L g8125 ( 
.A(n_7171),
.Y(n_8125)
);

INVx1_ASAP7_75t_L g8126 ( 
.A(n_7172),
.Y(n_8126)
);

NOR2xp33_ASAP7_75t_L g8127 ( 
.A(n_7655),
.B(n_2455),
.Y(n_8127)
);

INVx4_ASAP7_75t_SL g8128 ( 
.A(n_7647),
.Y(n_8128)
);

NOR2xp33_ASAP7_75t_L g8129 ( 
.A(n_7657),
.B(n_2455),
.Y(n_8129)
);

AOI21xp5_ASAP7_75t_L g8130 ( 
.A1(n_6953),
.A2(n_2457),
.B(n_2456),
.Y(n_8130)
);

INVx1_ASAP7_75t_L g8131 ( 
.A(n_7175),
.Y(n_8131)
);

INVx2_ASAP7_75t_SL g8132 ( 
.A(n_7090),
.Y(n_8132)
);

AND2x4_ASAP7_75t_L g8133 ( 
.A(n_7609),
.B(n_9),
.Y(n_8133)
);

BUFx6f_ASAP7_75t_L g8134 ( 
.A(n_7134),
.Y(n_8134)
);

AND2x2_ASAP7_75t_L g8135 ( 
.A(n_7691),
.B(n_9),
.Y(n_8135)
);

INVx2_ASAP7_75t_L g8136 ( 
.A(n_7176),
.Y(n_8136)
);

CKINVDCx5p33_ASAP7_75t_R g8137 ( 
.A(n_7652),
.Y(n_8137)
);

INVx1_ASAP7_75t_L g8138 ( 
.A(n_7177),
.Y(n_8138)
);

INVx2_ASAP7_75t_L g8139 ( 
.A(n_7181),
.Y(n_8139)
);

INVx1_ASAP7_75t_L g8140 ( 
.A(n_7187),
.Y(n_8140)
);

AND2x6_ASAP7_75t_L g8141 ( 
.A(n_7552),
.B(n_10),
.Y(n_8141)
);

AND2x2_ASAP7_75t_L g8142 ( 
.A(n_7718),
.B(n_10),
.Y(n_8142)
);

INVx1_ASAP7_75t_L g8143 ( 
.A(n_7191),
.Y(n_8143)
);

INVx1_ASAP7_75t_L g8144 ( 
.A(n_7196),
.Y(n_8144)
);

XNOR2x2_ASAP7_75t_SL g8145 ( 
.A(n_7425),
.B(n_10),
.Y(n_8145)
);

OAI21xp5_ASAP7_75t_L g8146 ( 
.A1(n_7658),
.A2(n_2457),
.B(n_2456),
.Y(n_8146)
);

NOR2xp33_ASAP7_75t_L g8147 ( 
.A(n_7659),
.B(n_2459),
.Y(n_8147)
);

INVx2_ASAP7_75t_L g8148 ( 
.A(n_7197),
.Y(n_8148)
);

INVx1_ASAP7_75t_L g8149 ( 
.A(n_7200),
.Y(n_8149)
);

INVx1_ASAP7_75t_L g8150 ( 
.A(n_7204),
.Y(n_8150)
);

INVx1_ASAP7_75t_L g8151 ( 
.A(n_7238),
.Y(n_8151)
);

INVx1_ASAP7_75t_L g8152 ( 
.A(n_7239),
.Y(n_8152)
);

INVx1_ASAP7_75t_L g8153 ( 
.A(n_7467),
.Y(n_8153)
);

NOR2xp33_ASAP7_75t_L g8154 ( 
.A(n_6972),
.B(n_2460),
.Y(n_8154)
);

BUFx6f_ASAP7_75t_L g8155 ( 
.A(n_7134),
.Y(n_8155)
);

INVxp33_ASAP7_75t_L g8156 ( 
.A(n_7328),
.Y(n_8156)
);

INVx1_ASAP7_75t_L g8157 ( 
.A(n_7499),
.Y(n_8157)
);

CKINVDCx20_ASAP7_75t_R g8158 ( 
.A(n_7640),
.Y(n_8158)
);

XNOR2x2_ASAP7_75t_L g8159 ( 
.A(n_7377),
.B(n_11),
.Y(n_8159)
);

INVx1_ASAP7_75t_L g8160 ( 
.A(n_7507),
.Y(n_8160)
);

INVx2_ASAP7_75t_L g8161 ( 
.A(n_7245),
.Y(n_8161)
);

INVx1_ASAP7_75t_L g8162 ( 
.A(n_7524),
.Y(n_8162)
);

XOR2xp5_ASAP7_75t_L g8163 ( 
.A(n_7234),
.B(n_11),
.Y(n_8163)
);

CKINVDCx5p33_ASAP7_75t_R g8164 ( 
.A(n_7685),
.Y(n_8164)
);

INVxp67_ASAP7_75t_L g8165 ( 
.A(n_7354),
.Y(n_8165)
);

INVx2_ASAP7_75t_L g8166 ( 
.A(n_7249),
.Y(n_8166)
);

INVx2_ASAP7_75t_L g8167 ( 
.A(n_7254),
.Y(n_8167)
);

INVx2_ASAP7_75t_L g8168 ( 
.A(n_7257),
.Y(n_8168)
);

INVx1_ASAP7_75t_L g8169 ( 
.A(n_7527),
.Y(n_8169)
);

BUFx6f_ASAP7_75t_L g8170 ( 
.A(n_7234),
.Y(n_8170)
);

AND2x2_ASAP7_75t_L g8171 ( 
.A(n_7224),
.B(n_11),
.Y(n_8171)
);

INVx1_ASAP7_75t_L g8172 ( 
.A(n_7528),
.Y(n_8172)
);

AND2x2_ASAP7_75t_L g8173 ( 
.A(n_7693),
.B(n_12),
.Y(n_8173)
);

INVx1_ASAP7_75t_L g8174 ( 
.A(n_7529),
.Y(n_8174)
);

NAND2xp33_ASAP7_75t_R g8175 ( 
.A(n_7264),
.B(n_12),
.Y(n_8175)
);

AND2x2_ASAP7_75t_L g8176 ( 
.A(n_7717),
.B(n_12),
.Y(n_8176)
);

NOR2xp33_ASAP7_75t_L g8177 ( 
.A(n_7518),
.B(n_2460),
.Y(n_8177)
);

INVx1_ASAP7_75t_L g8178 ( 
.A(n_7530),
.Y(n_8178)
);

INVx1_ASAP7_75t_L g8179 ( 
.A(n_7258),
.Y(n_8179)
);

BUFx3_ASAP7_75t_L g8180 ( 
.A(n_7235),
.Y(n_8180)
);

INVx1_ASAP7_75t_L g8181 ( 
.A(n_7474),
.Y(n_8181)
);

INVx1_ASAP7_75t_L g8182 ( 
.A(n_7480),
.Y(n_8182)
);

INVx1_ASAP7_75t_L g8183 ( 
.A(n_7482),
.Y(n_8183)
);

INVx1_ASAP7_75t_L g8184 ( 
.A(n_7427),
.Y(n_8184)
);

INVx4_ASAP7_75t_L g8185 ( 
.A(n_7235),
.Y(n_8185)
);

NAND2xp5_ASAP7_75t_L g8186 ( 
.A(n_7276),
.B(n_13),
.Y(n_8186)
);

INVx1_ASAP7_75t_L g8187 ( 
.A(n_7429),
.Y(n_8187)
);

INVx1_ASAP7_75t_L g8188 ( 
.A(n_7433),
.Y(n_8188)
);

INVx2_ASAP7_75t_L g8189 ( 
.A(n_7484),
.Y(n_8189)
);

CKINVDCx20_ASAP7_75t_R g8190 ( 
.A(n_7244),
.Y(n_8190)
);

INVx1_ASAP7_75t_L g8191 ( 
.A(n_7439),
.Y(n_8191)
);

INVx1_ASAP7_75t_L g8192 ( 
.A(n_7442),
.Y(n_8192)
);

XOR2xp5_ASAP7_75t_L g8193 ( 
.A(n_7244),
.B(n_14),
.Y(n_8193)
);

INVx1_ASAP7_75t_L g8194 ( 
.A(n_7444),
.Y(n_8194)
);

AND2x2_ASAP7_75t_L g8195 ( 
.A(n_7610),
.B(n_14),
.Y(n_8195)
);

INVx1_ASAP7_75t_L g8196 ( 
.A(n_7452),
.Y(n_8196)
);

INVx1_ASAP7_75t_L g8197 ( 
.A(n_7454),
.Y(n_8197)
);

INVx1_ASAP7_75t_L g8198 ( 
.A(n_7456),
.Y(n_8198)
);

INVx1_ASAP7_75t_L g8199 ( 
.A(n_7470),
.Y(n_8199)
);

INVx2_ASAP7_75t_SL g8200 ( 
.A(n_7262),
.Y(n_8200)
);

NOR2xp33_ASAP7_75t_L g8201 ( 
.A(n_7511),
.B(n_2461),
.Y(n_8201)
);

INVx2_ASAP7_75t_L g8202 ( 
.A(n_7473),
.Y(n_8202)
);

INVx1_ASAP7_75t_L g8203 ( 
.A(n_7478),
.Y(n_8203)
);

INVx1_ASAP7_75t_L g8204 ( 
.A(n_7479),
.Y(n_8204)
);

INVx1_ASAP7_75t_L g8205 ( 
.A(n_7535),
.Y(n_8205)
);

NOR2xp33_ASAP7_75t_L g8206 ( 
.A(n_7517),
.B(n_2461),
.Y(n_8206)
);

INVx1_ASAP7_75t_L g8207 ( 
.A(n_7539),
.Y(n_8207)
);

INVx2_ASAP7_75t_L g8208 ( 
.A(n_7488),
.Y(n_8208)
);

INVx2_ASAP7_75t_L g8209 ( 
.A(n_7496),
.Y(n_8209)
);

INVx1_ASAP7_75t_L g8210 ( 
.A(n_7540),
.Y(n_8210)
);

NOR2xp33_ASAP7_75t_L g8211 ( 
.A(n_7523),
.B(n_2462),
.Y(n_8211)
);

BUFx5_ASAP7_75t_L g8212 ( 
.A(n_7542),
.Y(n_8212)
);

XNOR2xp5_ASAP7_75t_L g8213 ( 
.A(n_7592),
.B(n_15),
.Y(n_8213)
);

INVx1_ASAP7_75t_L g8214 ( 
.A(n_7551),
.Y(n_8214)
);

INVx1_ASAP7_75t_L g8215 ( 
.A(n_7547),
.Y(n_8215)
);

NOR2xp67_ASAP7_75t_L g8216 ( 
.A(n_7318),
.B(n_15),
.Y(n_8216)
);

INVx2_ASAP7_75t_L g8217 ( 
.A(n_7505),
.Y(n_8217)
);

INVx1_ASAP7_75t_L g8218 ( 
.A(n_7497),
.Y(n_8218)
);

INVx1_ASAP7_75t_L g8219 ( 
.A(n_7500),
.Y(n_8219)
);

INVx1_ASAP7_75t_L g8220 ( 
.A(n_7504),
.Y(n_8220)
);

INVx1_ASAP7_75t_L g8221 ( 
.A(n_7679),
.Y(n_8221)
);

NOR2xp33_ASAP7_75t_L g8222 ( 
.A(n_7549),
.B(n_2462),
.Y(n_8222)
);

AND2x2_ASAP7_75t_L g8223 ( 
.A(n_7455),
.B(n_16),
.Y(n_8223)
);

BUFx2_ASAP7_75t_L g8224 ( 
.A(n_7046),
.Y(n_8224)
);

INVx1_ASAP7_75t_L g8225 ( 
.A(n_7680),
.Y(n_8225)
);

INVx1_ASAP7_75t_L g8226 ( 
.A(n_7506),
.Y(n_8226)
);

INVxp67_ASAP7_75t_SL g8227 ( 
.A(n_7288),
.Y(n_8227)
);

INVx1_ASAP7_75t_L g8228 ( 
.A(n_7509),
.Y(n_8228)
);

OR2x2_ASAP7_75t_SL g8229 ( 
.A(n_7350),
.B(n_16),
.Y(n_8229)
);

INVx1_ASAP7_75t_L g8230 ( 
.A(n_7516),
.Y(n_8230)
);

INVx1_ASAP7_75t_L g8231 ( 
.A(n_7521),
.Y(n_8231)
);

INVx1_ASAP7_75t_L g8232 ( 
.A(n_7531),
.Y(n_8232)
);

INVx2_ASAP7_75t_L g8233 ( 
.A(n_7532),
.Y(n_8233)
);

INVx1_ASAP7_75t_L g8234 ( 
.A(n_7173),
.Y(n_8234)
);

INVx2_ASAP7_75t_L g8235 ( 
.A(n_7566),
.Y(n_8235)
);

INVx1_ASAP7_75t_L g8236 ( 
.A(n_7671),
.Y(n_8236)
);

INVxp67_ASAP7_75t_SL g8237 ( 
.A(n_7328),
.Y(n_8237)
);

INVx1_ASAP7_75t_L g8238 ( 
.A(n_7675),
.Y(n_8238)
);

XNOR2x2_ASAP7_75t_L g8239 ( 
.A(n_7344),
.B(n_7441),
.Y(n_8239)
);

AND2x2_ASAP7_75t_L g8240 ( 
.A(n_7581),
.B(n_16),
.Y(n_8240)
);

AND2x2_ASAP7_75t_L g8241 ( 
.A(n_7581),
.B(n_17),
.Y(n_8241)
);

CKINVDCx5p33_ASAP7_75t_R g8242 ( 
.A(n_7262),
.Y(n_8242)
);

INVx1_ASAP7_75t_L g8243 ( 
.A(n_7683),
.Y(n_8243)
);

INVx1_ASAP7_75t_L g8244 ( 
.A(n_7072),
.Y(n_8244)
);

INVx1_ASAP7_75t_L g8245 ( 
.A(n_7107),
.Y(n_8245)
);

NAND2xp5_ASAP7_75t_L g8246 ( 
.A(n_7034),
.B(n_17),
.Y(n_8246)
);

AND2x2_ASAP7_75t_L g8247 ( 
.A(n_7593),
.B(n_18),
.Y(n_8247)
);

CKINVDCx20_ASAP7_75t_R g8248 ( 
.A(n_7267),
.Y(n_8248)
);

INVx1_ASAP7_75t_L g8249 ( 
.A(n_7164),
.Y(n_8249)
);

INVx2_ASAP7_75t_L g8250 ( 
.A(n_7568),
.Y(n_8250)
);

NAND2x1p5_ASAP7_75t_L g8251 ( 
.A(n_7030),
.B(n_19),
.Y(n_8251)
);

CKINVDCx16_ASAP7_75t_R g8252 ( 
.A(n_7046),
.Y(n_8252)
);

INVxp33_ASAP7_75t_L g8253 ( 
.A(n_7378),
.Y(n_8253)
);

INVx1_ASAP7_75t_L g8254 ( 
.A(n_7286),
.Y(n_8254)
);

NOR2xp33_ASAP7_75t_L g8255 ( 
.A(n_7215),
.B(n_2463),
.Y(n_8255)
);

INVx1_ASAP7_75t_L g8256 ( 
.A(n_7574),
.Y(n_8256)
);

INVx1_ASAP7_75t_L g8257 ( 
.A(n_7576),
.Y(n_8257)
);

NOR2x1_ASAP7_75t_L g8258 ( 
.A(n_7486),
.B(n_19),
.Y(n_8258)
);

XOR2xp5_ASAP7_75t_L g8259 ( 
.A(n_7267),
.B(n_19),
.Y(n_8259)
);

INVx1_ASAP7_75t_L g8260 ( 
.A(n_7583),
.Y(n_8260)
);

XOR2xp5_ASAP7_75t_L g8261 ( 
.A(n_7461),
.B(n_7378),
.Y(n_8261)
);

INVx1_ASAP7_75t_L g8262 ( 
.A(n_7591),
.Y(n_8262)
);

INVx1_ASAP7_75t_L g8263 ( 
.A(n_7598),
.Y(n_8263)
);

INVx1_ASAP7_75t_L g8264 ( 
.A(n_7614),
.Y(n_8264)
);

AOI21xp5_ASAP7_75t_L g8265 ( 
.A1(n_7459),
.A2(n_2464),
.B(n_2463),
.Y(n_8265)
);

INVx1_ASAP7_75t_L g8266 ( 
.A(n_7615),
.Y(n_8266)
);

BUFx6f_ASAP7_75t_L g8267 ( 
.A(n_7379),
.Y(n_8267)
);

INVx2_ASAP7_75t_L g8268 ( 
.A(n_7618),
.Y(n_8268)
);

NAND2xp5_ASAP7_75t_SL g8269 ( 
.A(n_7379),
.B(n_2464),
.Y(n_8269)
);

INVx1_ASAP7_75t_L g8270 ( 
.A(n_7619),
.Y(n_8270)
);

NAND2xp5_ASAP7_75t_L g8271 ( 
.A(n_7222),
.B(n_20),
.Y(n_8271)
);

INVx1_ASAP7_75t_L g8272 ( 
.A(n_7624),
.Y(n_8272)
);

INVx1_ASAP7_75t_L g8273 ( 
.A(n_7629),
.Y(n_8273)
);

NOR2xp33_ASAP7_75t_L g8274 ( 
.A(n_7510),
.B(n_2465),
.Y(n_8274)
);

NAND2xp5_ASAP7_75t_L g8275 ( 
.A(n_7085),
.B(n_20),
.Y(n_8275)
);

AND2x2_ASAP7_75t_L g8276 ( 
.A(n_7593),
.B(n_21),
.Y(n_8276)
);

BUFx5_ASAP7_75t_L g8277 ( 
.A(n_7019),
.Y(n_8277)
);

INVx1_ASAP7_75t_L g8278 ( 
.A(n_7630),
.Y(n_8278)
);

OAI21xp5_ASAP7_75t_L g8279 ( 
.A1(n_7550),
.A2(n_2466),
.B(n_2465),
.Y(n_8279)
);

INVx1_ASAP7_75t_L g8280 ( 
.A(n_7634),
.Y(n_8280)
);

INVx1_ASAP7_75t_L g8281 ( 
.A(n_7638),
.Y(n_8281)
);

INVxp33_ASAP7_75t_L g8282 ( 
.A(n_7402),
.Y(n_8282)
);

INVx1_ASAP7_75t_L g8283 ( 
.A(n_7643),
.Y(n_8283)
);

XOR2xp5_ASAP7_75t_L g8284 ( 
.A(n_7402),
.B(n_21),
.Y(n_8284)
);

AND2x2_ASAP7_75t_L g8285 ( 
.A(n_7385),
.B(n_21),
.Y(n_8285)
);

XNOR2x2_ASAP7_75t_L g8286 ( 
.A(n_7424),
.B(n_23),
.Y(n_8286)
);

INVx1_ASAP7_75t_SL g8287 ( 
.A(n_7075),
.Y(n_8287)
);

INVx1_ASAP7_75t_L g8288 ( 
.A(n_7644),
.Y(n_8288)
);

INVx1_ASAP7_75t_L g8289 ( 
.A(n_7654),
.Y(n_8289)
);

INVx1_ASAP7_75t_SL g8290 ( 
.A(n_7075),
.Y(n_8290)
);

INVx1_ASAP7_75t_L g8291 ( 
.A(n_7656),
.Y(n_8291)
);

AND2x2_ASAP7_75t_L g8292 ( 
.A(n_7211),
.B(n_23),
.Y(n_8292)
);

NAND2xp5_ASAP7_75t_L g8293 ( 
.A(n_7109),
.B(n_23),
.Y(n_8293)
);

AND2x2_ASAP7_75t_L g8294 ( 
.A(n_7087),
.B(n_7101),
.Y(n_8294)
);

BUFx6f_ASAP7_75t_L g8295 ( 
.A(n_7413),
.Y(n_8295)
);

INVx2_ASAP7_75t_L g8296 ( 
.A(n_7660),
.Y(n_8296)
);

INVx1_ASAP7_75t_L g8297 ( 
.A(n_7661),
.Y(n_8297)
);

INVx2_ASAP7_75t_L g8298 ( 
.A(n_7665),
.Y(n_8298)
);

INVx1_ASAP7_75t_L g8299 ( 
.A(n_7713),
.Y(n_8299)
);

AND2x2_ASAP7_75t_L g8300 ( 
.A(n_7087),
.B(n_24),
.Y(n_8300)
);

INVx1_ASAP7_75t_L g8301 ( 
.A(n_7538),
.Y(n_8301)
);

INVx1_ASAP7_75t_L g8302 ( 
.A(n_7077),
.Y(n_8302)
);

INVx1_ASAP7_75t_L g8303 ( 
.A(n_7170),
.Y(n_8303)
);

NAND2xp5_ASAP7_75t_L g8304 ( 
.A(n_6999),
.B(n_24),
.Y(n_8304)
);

INVx2_ASAP7_75t_L g8305 ( 
.A(n_7537),
.Y(n_8305)
);

INVx1_ASAP7_75t_L g8306 ( 
.A(n_7182),
.Y(n_8306)
);

INVxp67_ASAP7_75t_L g8307 ( 
.A(n_7413),
.Y(n_8307)
);

INVxp67_ASAP7_75t_SL g8308 ( 
.A(n_7416),
.Y(n_8308)
);

NOR2xp33_ASAP7_75t_L g8309 ( 
.A(n_7360),
.B(n_2467),
.Y(n_8309)
);

NAND2xp5_ASAP7_75t_SL g8310 ( 
.A(n_7416),
.B(n_2467),
.Y(n_8310)
);

AND2x2_ASAP7_75t_L g8311 ( 
.A(n_7101),
.B(n_7102),
.Y(n_8311)
);

INVx1_ASAP7_75t_L g8312 ( 
.A(n_7185),
.Y(n_8312)
);

INVx1_ASAP7_75t_L g8313 ( 
.A(n_7194),
.Y(n_8313)
);

NOR2xp33_ASAP7_75t_L g8314 ( 
.A(n_7443),
.B(n_2468),
.Y(n_8314)
);

INVx1_ASAP7_75t_L g8315 ( 
.A(n_7251),
.Y(n_8315)
);

NOR2xp33_ASAP7_75t_L g8316 ( 
.A(n_7558),
.B(n_2468),
.Y(n_8316)
);

INVx5_ASAP7_75t_L g8317 ( 
.A(n_7019),
.Y(n_8317)
);

AND2x2_ASAP7_75t_L g8318 ( 
.A(n_7102),
.B(n_24),
.Y(n_8318)
);

INVxp33_ASAP7_75t_L g8319 ( 
.A(n_7430),
.Y(n_8319)
);

INVx1_ASAP7_75t_L g8320 ( 
.A(n_7277),
.Y(n_8320)
);

INVx4_ASAP7_75t_SL g8321 ( 
.A(n_7464),
.Y(n_8321)
);

INVx1_ASAP7_75t_L g8322 ( 
.A(n_7280),
.Y(n_8322)
);

INVx1_ASAP7_75t_L g8323 ( 
.A(n_7283),
.Y(n_8323)
);

NAND2xp5_ASAP7_75t_L g8324 ( 
.A(n_7294),
.B(n_25),
.Y(n_8324)
);

INVx1_ASAP7_75t_L g8325 ( 
.A(n_7296),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_7300),
.Y(n_8326)
);

CKINVDCx20_ASAP7_75t_R g8327 ( 
.A(n_7068),
.Y(n_8327)
);

AND2x4_ASAP7_75t_L g8328 ( 
.A(n_7687),
.B(n_25),
.Y(n_8328)
);

INVx1_ASAP7_75t_L g8329 ( 
.A(n_7588),
.Y(n_8329)
);

INVx1_ASAP7_75t_L g8330 ( 
.A(n_7571),
.Y(n_8330)
);

INVx1_ASAP7_75t_L g8331 ( 
.A(n_7358),
.Y(n_8331)
);

XNOR2x2_ASAP7_75t_L g8332 ( 
.A(n_7293),
.B(n_25),
.Y(n_8332)
);

AND2x2_ASAP7_75t_L g8333 ( 
.A(n_7104),
.B(n_26),
.Y(n_8333)
);

INVx2_ASAP7_75t_L g8334 ( 
.A(n_7544),
.Y(n_8334)
);

INVx1_ASAP7_75t_L g8335 ( 
.A(n_7365),
.Y(n_8335)
);

INVx1_ASAP7_75t_L g8336 ( 
.A(n_7390),
.Y(n_8336)
);

NOR2xp33_ASAP7_75t_SL g8337 ( 
.A(n_7130),
.B(n_7140),
.Y(n_8337)
);

INVx1_ASAP7_75t_L g8338 ( 
.A(n_7457),
.Y(n_8338)
);

NOR2xp33_ASAP7_75t_L g8339 ( 
.A(n_7580),
.B(n_2470),
.Y(n_8339)
);

INVx1_ASAP7_75t_L g8340 ( 
.A(n_7559),
.Y(n_8340)
);

INVxp33_ASAP7_75t_SL g8341 ( 
.A(n_7241),
.Y(n_8341)
);

INVx1_ASAP7_75t_L g8342 ( 
.A(n_7559),
.Y(n_8342)
);

INVx1_ASAP7_75t_L g8343 ( 
.A(n_7559),
.Y(n_8343)
);

XNOR2xp5_ASAP7_75t_L g8344 ( 
.A(n_7584),
.B(n_26),
.Y(n_8344)
);

INVx1_ASAP7_75t_L g8345 ( 
.A(n_7706),
.Y(n_8345)
);

INVx1_ASAP7_75t_L g8346 ( 
.A(n_7707),
.Y(n_8346)
);

NOR2xp33_ASAP7_75t_L g8347 ( 
.A(n_7596),
.B(n_2470),
.Y(n_8347)
);

NAND2xp5_ASAP7_75t_L g8348 ( 
.A(n_7246),
.B(n_26),
.Y(n_8348)
);

NAND2x1p5_ASAP7_75t_L g8349 ( 
.A(n_7143),
.B(n_27),
.Y(n_8349)
);

INVx1_ASAP7_75t_L g8350 ( 
.A(n_7708),
.Y(n_8350)
);

NAND2xp33_ASAP7_75t_SL g8351 ( 
.A(n_7722),
.B(n_7724),
.Y(n_8351)
);

INVx1_ASAP7_75t_L g8352 ( 
.A(n_7689),
.Y(n_8352)
);

INVx2_ASAP7_75t_L g8353 ( 
.A(n_7548),
.Y(n_8353)
);

INVx1_ASAP7_75t_L g8354 ( 
.A(n_7692),
.Y(n_8354)
);

INVx1_ASAP7_75t_L g8355 ( 
.A(n_7695),
.Y(n_8355)
);

INVx1_ASAP7_75t_L g8356 ( 
.A(n_7710),
.Y(n_8356)
);

INVx4_ASAP7_75t_L g8357 ( 
.A(n_7430),
.Y(n_8357)
);

INVx2_ASAP7_75t_L g8358 ( 
.A(n_7560),
.Y(n_8358)
);

NOR2xp67_ASAP7_75t_L g8359 ( 
.A(n_7498),
.B(n_27),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_7097),
.Y(n_8360)
);

NOR2xp33_ASAP7_75t_L g8361 ( 
.A(n_7022),
.B(n_2471),
.Y(n_8361)
);

INVx1_ASAP7_75t_L g8362 ( 
.A(n_7136),
.Y(n_8362)
);

INVx1_ASAP7_75t_L g8363 ( 
.A(n_7149),
.Y(n_8363)
);

XNOR2xp5_ASAP7_75t_L g8364 ( 
.A(n_7613),
.B(n_27),
.Y(n_8364)
);

AND2x2_ASAP7_75t_L g8365 ( 
.A(n_7104),
.B(n_28),
.Y(n_8365)
);

INVx1_ASAP7_75t_L g8366 ( 
.A(n_7160),
.Y(n_8366)
);

INVx1_ASAP7_75t_L g8367 ( 
.A(n_7700),
.Y(n_8367)
);

INVx1_ASAP7_75t_SL g8368 ( 
.A(n_7155),
.Y(n_8368)
);

INVx1_ASAP7_75t_L g8369 ( 
.A(n_7701),
.Y(n_8369)
);

NOR2xp33_ASAP7_75t_L g8370 ( 
.A(n_7611),
.B(n_2471),
.Y(n_8370)
);

INVxp67_ASAP7_75t_L g8371 ( 
.A(n_7436),
.Y(n_8371)
);

NAND2x1p5_ASAP7_75t_L g8372 ( 
.A(n_7250),
.B(n_28),
.Y(n_8372)
);

XNOR2xp5_ASAP7_75t_L g8373 ( 
.A(n_7155),
.B(n_28),
.Y(n_8373)
);

NOR2xp67_ASAP7_75t_L g8374 ( 
.A(n_7522),
.B(n_29),
.Y(n_8374)
);

NAND2xp5_ASAP7_75t_SL g8375 ( 
.A(n_7436),
.B(n_2472),
.Y(n_8375)
);

INVx1_ASAP7_75t_L g8376 ( 
.A(n_7702),
.Y(n_8376)
);

INVx1_ASAP7_75t_L g8377 ( 
.A(n_7703),
.Y(n_8377)
);

INVx3_ASAP7_75t_L g8378 ( 
.A(n_7341),
.Y(n_8378)
);

HB1xp67_ASAP7_75t_L g8379 ( 
.A(n_7096),
.Y(n_8379)
);

AND2x2_ASAP7_75t_L g8380 ( 
.A(n_7362),
.B(n_29),
.Y(n_8380)
);

AND2x4_ASAP7_75t_L g8381 ( 
.A(n_7536),
.B(n_29),
.Y(n_8381)
);

CKINVDCx16_ASAP7_75t_R g8382 ( 
.A(n_7019),
.Y(n_8382)
);

INVx1_ASAP7_75t_L g8383 ( 
.A(n_7188),
.Y(n_8383)
);

INVx1_ASAP7_75t_L g8384 ( 
.A(n_7216),
.Y(n_8384)
);

INVx1_ASAP7_75t_L g8385 ( 
.A(n_7228),
.Y(n_8385)
);

AND2x4_ASAP7_75t_L g8386 ( 
.A(n_7570),
.B(n_30),
.Y(n_8386)
);

INVx1_ASAP7_75t_L g8387 ( 
.A(n_7232),
.Y(n_8387)
);

INVx1_ASAP7_75t_L g8388 ( 
.A(n_7255),
.Y(n_8388)
);

INVx1_ASAP7_75t_L g8389 ( 
.A(n_7721),
.Y(n_8389)
);

INVx1_ASAP7_75t_L g8390 ( 
.A(n_7723),
.Y(n_8390)
);

INVx1_ASAP7_75t_L g8391 ( 
.A(n_7589),
.Y(n_8391)
);

XOR2xp5_ASAP7_75t_L g8392 ( 
.A(n_7503),
.B(n_31),
.Y(n_8392)
);

NOR2xp33_ASAP7_75t_L g8393 ( 
.A(n_6959),
.B(n_2473),
.Y(n_8393)
);

INVx1_ASAP7_75t_L g8394 ( 
.A(n_7214),
.Y(n_8394)
);

INVx1_ASAP7_75t_L g8395 ( 
.A(n_6963),
.Y(n_8395)
);

AND2x2_ASAP7_75t_L g8396 ( 
.A(n_7612),
.B(n_31),
.Y(n_8396)
);

INVx1_ASAP7_75t_L g8397 ( 
.A(n_7352),
.Y(n_8397)
);

XNOR2x2_ASAP7_75t_L g8398 ( 
.A(n_7513),
.B(n_32),
.Y(n_8398)
);

INVx1_ASAP7_75t_L g8399 ( 
.A(n_7367),
.Y(n_8399)
);

AND2x2_ASAP7_75t_L g8400 ( 
.A(n_7273),
.B(n_32),
.Y(n_8400)
);

INVx1_ASAP7_75t_L g8401 ( 
.A(n_7375),
.Y(n_8401)
);

AND2x2_ASAP7_75t_L g8402 ( 
.A(n_7297),
.B(n_33),
.Y(n_8402)
);

INVx1_ASAP7_75t_L g8403 ( 
.A(n_7387),
.Y(n_8403)
);

INVx1_ASAP7_75t_L g8404 ( 
.A(n_7401),
.Y(n_8404)
);

AOI21xp5_ASAP7_75t_L g8405 ( 
.A1(n_7469),
.A2(n_2474),
.B(n_2473),
.Y(n_8405)
);

INVx1_ASAP7_75t_L g8406 ( 
.A(n_7414),
.Y(n_8406)
);

INVxp33_ASAP7_75t_L g8407 ( 
.A(n_7553),
.Y(n_8407)
);

AND2x2_ASAP7_75t_L g8408 ( 
.A(n_7201),
.B(n_33),
.Y(n_8408)
);

INVx1_ASAP7_75t_L g8409 ( 
.A(n_7453),
.Y(n_8409)
);

INVx1_ASAP7_75t_L g8410 ( 
.A(n_7962),
.Y(n_8410)
);

BUFx6f_ASAP7_75t_L g8411 ( 
.A(n_7735),
.Y(n_8411)
);

CKINVDCx5p33_ASAP7_75t_R g8412 ( 
.A(n_7734),
.Y(n_8412)
);

INVx2_ASAP7_75t_SL g8413 ( 
.A(n_7738),
.Y(n_8413)
);

INVx1_ASAP7_75t_L g8414 ( 
.A(n_7729),
.Y(n_8414)
);

NAND2xp5_ASAP7_75t_L g8415 ( 
.A(n_8036),
.B(n_7464),
.Y(n_8415)
);

INVx2_ASAP7_75t_L g8416 ( 
.A(n_7753),
.Y(n_8416)
);

INVx2_ASAP7_75t_L g8417 ( 
.A(n_7772),
.Y(n_8417)
);

AND2x2_ASAP7_75t_L g8418 ( 
.A(n_7829),
.B(n_7616),
.Y(n_8418)
);

NAND2xp5_ASAP7_75t_L g8419 ( 
.A(n_7731),
.B(n_7744),
.Y(n_8419)
);

NAND2xp5_ASAP7_75t_SL g8420 ( 
.A(n_7763),
.B(n_7017),
.Y(n_8420)
);

NAND2xp5_ASAP7_75t_L g8421 ( 
.A(n_8341),
.B(n_7464),
.Y(n_8421)
);

NAND2xp5_ASAP7_75t_L g8422 ( 
.A(n_7935),
.B(n_7060),
.Y(n_8422)
);

INVx2_ASAP7_75t_L g8423 ( 
.A(n_7778),
.Y(n_8423)
);

AOI22xp33_ASAP7_75t_L g8424 ( 
.A1(n_7732),
.A2(n_7904),
.B1(n_7774),
.B2(n_7941),
.Y(n_8424)
);

INVx2_ASAP7_75t_L g8425 ( 
.A(n_7789),
.Y(n_8425)
);

AO221x1_ASAP7_75t_L g8426 ( 
.A1(n_8145),
.A2(n_7252),
.B1(n_7422),
.B2(n_7431),
.C(n_7476),
.Y(n_8426)
);

NOR2xp33_ASAP7_75t_L g8427 ( 
.A(n_7876),
.B(n_7292),
.Y(n_8427)
);

INVx2_ASAP7_75t_L g8428 ( 
.A(n_7808),
.Y(n_8428)
);

BUFx3_ASAP7_75t_L g8429 ( 
.A(n_8190),
.Y(n_8429)
);

NOR2xp33_ASAP7_75t_L g8430 ( 
.A(n_7988),
.B(n_7326),
.Y(n_8430)
);

BUFx12f_ASAP7_75t_L g8431 ( 
.A(n_7977),
.Y(n_8431)
);

AND2x4_ASAP7_75t_SL g8432 ( 
.A(n_7820),
.B(n_7597),
.Y(n_8432)
);

A2O1A1Ixp33_ASAP7_75t_L g8433 ( 
.A1(n_8201),
.A2(n_7686),
.B(n_7061),
.C(n_7632),
.Y(n_8433)
);

AND2x4_ASAP7_75t_L g8434 ( 
.A(n_8124),
.B(n_7010),
.Y(n_8434)
);

INVx2_ASAP7_75t_L g8435 ( 
.A(n_7819),
.Y(n_8435)
);

NAND2xp5_ASAP7_75t_SL g8436 ( 
.A(n_7823),
.B(n_7074),
.Y(n_8436)
);

A2O1A1Ixp33_ASAP7_75t_L g8437 ( 
.A1(n_8206),
.A2(n_7631),
.B(n_7603),
.C(n_7490),
.Y(n_8437)
);

INVx2_ASAP7_75t_L g8438 ( 
.A(n_7826),
.Y(n_8438)
);

INVx1_ASAP7_75t_L g8439 ( 
.A(n_7740),
.Y(n_8439)
);

NOR2xp33_ASAP7_75t_L g8440 ( 
.A(n_8048),
.B(n_7027),
.Y(n_8440)
);

INVx1_ASAP7_75t_L g8441 ( 
.A(n_7745),
.Y(n_8441)
);

AND2x6_ASAP7_75t_SL g8442 ( 
.A(n_7874),
.B(n_7121),
.Y(n_8442)
);

NAND2xp5_ASAP7_75t_L g8443 ( 
.A(n_8000),
.B(n_7475),
.Y(n_8443)
);

AOI22xp5_ASAP7_75t_L g8444 ( 
.A1(n_8255),
.A2(n_7278),
.B1(n_7569),
.B2(n_7458),
.Y(n_8444)
);

NAND2xp5_ASAP7_75t_L g8445 ( 
.A(n_7736),
.B(n_7489),
.Y(n_8445)
);

NAND2xp5_ASAP7_75t_L g8446 ( 
.A(n_8093),
.B(n_7491),
.Y(n_8446)
);

NAND2xp5_ASAP7_75t_L g8447 ( 
.A(n_7764),
.B(n_7525),
.Y(n_8447)
);

INVx4_ASAP7_75t_L g8448 ( 
.A(n_8051),
.Y(n_8448)
);

INVx2_ASAP7_75t_L g8449 ( 
.A(n_7844),
.Y(n_8449)
);

NAND2xp5_ASAP7_75t_SL g8450 ( 
.A(n_8317),
.B(n_7031),
.Y(n_8450)
);

AND2x2_ASAP7_75t_SL g8451 ( 
.A(n_8382),
.B(n_7543),
.Y(n_8451)
);

INVx2_ASAP7_75t_L g8452 ( 
.A(n_7848),
.Y(n_8452)
);

INVx2_ASAP7_75t_SL g8453 ( 
.A(n_7859),
.Y(n_8453)
);

INVx2_ASAP7_75t_SL g8454 ( 
.A(n_8242),
.Y(n_8454)
);

NAND2xp5_ASAP7_75t_L g8455 ( 
.A(n_7751),
.B(n_7546),
.Y(n_8455)
);

NOR2xp67_ASAP7_75t_L g8456 ( 
.A(n_7834),
.B(n_7651),
.Y(n_8456)
);

NAND2xp5_ASAP7_75t_L g8457 ( 
.A(n_8302),
.B(n_7555),
.Y(n_8457)
);

INVx1_ASAP7_75t_L g8458 ( 
.A(n_7749),
.Y(n_8458)
);

NOR2xp33_ASAP7_75t_L g8459 ( 
.A(n_8115),
.B(n_8407),
.Y(n_8459)
);

INVx2_ASAP7_75t_L g8460 ( 
.A(n_7855),
.Y(n_8460)
);

INVx1_ASAP7_75t_L g8461 ( 
.A(n_7750),
.Y(n_8461)
);

INVx1_ASAP7_75t_L g8462 ( 
.A(n_7752),
.Y(n_8462)
);

NAND2xp5_ASAP7_75t_L g8463 ( 
.A(n_8303),
.B(n_7037),
.Y(n_8463)
);

NOR2x1p5_ASAP7_75t_L g8464 ( 
.A(n_7885),
.B(n_7044),
.Y(n_8464)
);

NAND2xp5_ASAP7_75t_SL g8465 ( 
.A(n_8317),
.B(n_7086),
.Y(n_8465)
);

INVx1_ASAP7_75t_L g8466 ( 
.A(n_7754),
.Y(n_8466)
);

NOR3xp33_ASAP7_75t_L g8467 ( 
.A(n_8100),
.B(n_8177),
.C(n_7742),
.Y(n_8467)
);

AOI22xp5_ASAP7_75t_L g8468 ( 
.A1(n_8309),
.A2(n_7346),
.B1(n_7345),
.B2(n_7115),
.Y(n_8468)
);

INVx2_ASAP7_75t_L g8469 ( 
.A(n_7865),
.Y(n_8469)
);

INVx2_ASAP7_75t_L g8470 ( 
.A(n_7880),
.Y(n_8470)
);

INVx1_ASAP7_75t_L g8471 ( 
.A(n_7755),
.Y(n_8471)
);

INVx2_ASAP7_75t_L g8472 ( 
.A(n_7940),
.Y(n_8472)
);

NAND2xp5_ASAP7_75t_L g8473 ( 
.A(n_8306),
.B(n_7099),
.Y(n_8473)
);

INVx4_ASAP7_75t_L g8474 ( 
.A(n_7921),
.Y(n_8474)
);

NOR2xp33_ASAP7_75t_L g8475 ( 
.A(n_7822),
.B(n_7071),
.Y(n_8475)
);

INVxp67_ASAP7_75t_SL g8476 ( 
.A(n_8019),
.Y(n_8476)
);

NOR2xp33_ASAP7_75t_L g8477 ( 
.A(n_7918),
.B(n_7483),
.Y(n_8477)
);

AOI22xp5_ASAP7_75t_L g8478 ( 
.A1(n_8314),
.A2(n_7144),
.B1(n_7150),
.B2(n_7331),
.Y(n_8478)
);

NAND2xp5_ASAP7_75t_L g8479 ( 
.A(n_8312),
.B(n_7147),
.Y(n_8479)
);

INVx1_ASAP7_75t_L g8480 ( 
.A(n_7756),
.Y(n_8480)
);

AOI21xp5_ASAP7_75t_L g8481 ( 
.A1(n_8089),
.A2(n_7669),
.B(n_6976),
.Y(n_8481)
);

INVx2_ASAP7_75t_L g8482 ( 
.A(n_7950),
.Y(n_8482)
);

INVx2_ASAP7_75t_L g8483 ( 
.A(n_7955),
.Y(n_8483)
);

AOI22x1_ASAP7_75t_L g8484 ( 
.A1(n_8279),
.A2(n_7623),
.B1(n_7639),
.B2(n_7600),
.Y(n_8484)
);

INVx1_ASAP7_75t_L g8485 ( 
.A(n_7757),
.Y(n_8485)
);

INVx1_ASAP7_75t_L g8486 ( 
.A(n_7759),
.Y(n_8486)
);

NOR2xp33_ASAP7_75t_L g8487 ( 
.A(n_7730),
.B(n_7157),
.Y(n_8487)
);

INVx2_ASAP7_75t_L g8488 ( 
.A(n_7971),
.Y(n_8488)
);

NAND2xp5_ASAP7_75t_L g8489 ( 
.A(n_8313),
.B(n_8315),
.Y(n_8489)
);

NAND2xp5_ASAP7_75t_L g8490 ( 
.A(n_8320),
.B(n_7167),
.Y(n_8490)
);

A2O1A1Ixp33_ASAP7_75t_L g8491 ( 
.A1(n_8211),
.A2(n_7512),
.B(n_7646),
.C(n_7400),
.Y(n_8491)
);

NAND2xp5_ASAP7_75t_SL g8492 ( 
.A(n_8317),
.B(n_7582),
.Y(n_8492)
);

INVx1_ASAP7_75t_L g8493 ( 
.A(n_7761),
.Y(n_8493)
);

INVx2_ASAP7_75t_L g8494 ( 
.A(n_7998),
.Y(n_8494)
);

NOR2xp33_ASAP7_75t_L g8495 ( 
.A(n_7773),
.B(n_7334),
.Y(n_8495)
);

NAND2xp5_ASAP7_75t_L g8496 ( 
.A(n_8322),
.B(n_7625),
.Y(n_8496)
);

NOR2xp33_ASAP7_75t_L g8497 ( 
.A(n_7739),
.B(n_7667),
.Y(n_8497)
);

INVx1_ASAP7_75t_L g8498 ( 
.A(n_7765),
.Y(n_8498)
);

NAND2xp5_ASAP7_75t_L g8499 ( 
.A(n_8323),
.B(n_8325),
.Y(n_8499)
);

INVx2_ASAP7_75t_L g8500 ( 
.A(n_8011),
.Y(n_8500)
);

A2O1A1Ixp33_ASAP7_75t_L g8501 ( 
.A1(n_8222),
.A2(n_8316),
.B(n_8339),
.C(n_8274),
.Y(n_8501)
);

NAND3xp33_ASAP7_75t_L g8502 ( 
.A(n_7758),
.B(n_7417),
.C(n_7412),
.Y(n_8502)
);

NAND2xp5_ASAP7_75t_L g8503 ( 
.A(n_8326),
.B(n_7628),
.Y(n_8503)
);

INVx2_ASAP7_75t_L g8504 ( 
.A(n_8015),
.Y(n_8504)
);

NAND2xp5_ASAP7_75t_L g8505 ( 
.A(n_8331),
.B(n_7645),
.Y(n_8505)
);

NAND2xp5_ASAP7_75t_L g8506 ( 
.A(n_8335),
.B(n_8336),
.Y(n_8506)
);

NAND2xp5_ASAP7_75t_L g8507 ( 
.A(n_8338),
.B(n_7567),
.Y(n_8507)
);

OAI22xp33_ASAP7_75t_L g8508 ( 
.A1(n_8098),
.A2(n_7684),
.B1(n_7696),
.B2(n_7682),
.Y(n_8508)
);

HB1xp67_ASAP7_75t_L g8509 ( 
.A(n_7781),
.Y(n_8509)
);

INVx2_ASAP7_75t_L g8510 ( 
.A(n_8016),
.Y(n_8510)
);

INVx1_ASAP7_75t_L g8511 ( 
.A(n_7766),
.Y(n_8511)
);

OR2x2_ASAP7_75t_L g8512 ( 
.A(n_8064),
.B(n_7699),
.Y(n_8512)
);

AND2x6_ASAP7_75t_L g8513 ( 
.A(n_8391),
.B(n_7668),
.Y(n_8513)
);

NAND2xp5_ASAP7_75t_L g8514 ( 
.A(n_7993),
.B(n_7572),
.Y(n_8514)
);

INVx1_ASAP7_75t_L g8515 ( 
.A(n_7768),
.Y(n_8515)
);

NAND2xp5_ASAP7_75t_SL g8516 ( 
.A(n_8061),
.B(n_7697),
.Y(n_8516)
);

INVx1_ASAP7_75t_SL g8517 ( 
.A(n_7980),
.Y(n_8517)
);

NAND2xp5_ASAP7_75t_L g8518 ( 
.A(n_7994),
.B(n_8003),
.Y(n_8518)
);

NAND2xp5_ASAP7_75t_L g8519 ( 
.A(n_8014),
.B(n_7838),
.Y(n_8519)
);

NOR2xp67_ASAP7_75t_L g8520 ( 
.A(n_8165),
.B(n_7586),
.Y(n_8520)
);

NAND2xp5_ASAP7_75t_L g8521 ( 
.A(n_7872),
.B(n_7602),
.Y(n_8521)
);

NOR2xp33_ASAP7_75t_L g8522 ( 
.A(n_7806),
.B(n_7186),
.Y(n_8522)
);

NOR2xp33_ASAP7_75t_L g8523 ( 
.A(n_7733),
.B(n_7633),
.Y(n_8523)
);

NAND2xp5_ASAP7_75t_SL g8524 ( 
.A(n_8212),
.B(n_7641),
.Y(n_8524)
);

NAND2xp5_ASAP7_75t_L g8525 ( 
.A(n_8041),
.B(n_7662),
.Y(n_8525)
);

NAND2xp5_ASAP7_75t_L g8526 ( 
.A(n_7897),
.B(n_7666),
.Y(n_8526)
);

AND2x2_ASAP7_75t_L g8527 ( 
.A(n_7957),
.B(n_7601),
.Y(n_8527)
);

INVx2_ASAP7_75t_L g8528 ( 
.A(n_7978),
.Y(n_8528)
);

INVx1_ASAP7_75t_L g8529 ( 
.A(n_7769),
.Y(n_8529)
);

INVx2_ASAP7_75t_L g8530 ( 
.A(n_7979),
.Y(n_8530)
);

AOI22xp33_ASAP7_75t_L g8531 ( 
.A1(n_8027),
.A2(n_7063),
.B1(n_7541),
.B2(n_7184),
.Y(n_8531)
);

INVx2_ASAP7_75t_L g8532 ( 
.A(n_7982),
.Y(n_8532)
);

NOR2xp67_ASAP7_75t_L g8533 ( 
.A(n_8378),
.B(n_7748),
.Y(n_8533)
);

O2A1O1Ixp33_ASAP7_75t_L g8534 ( 
.A1(n_7973),
.A2(n_7178),
.B(n_6974),
.C(n_7000),
.Y(n_8534)
);

NAND2xp5_ASAP7_75t_L g8535 ( 
.A(n_7892),
.B(n_7653),
.Y(n_8535)
);

NAND2xp5_ASAP7_75t_L g8536 ( 
.A(n_8046),
.B(n_7677),
.Y(n_8536)
);

NAND2xp5_ASAP7_75t_L g8537 ( 
.A(n_7931),
.B(n_7965),
.Y(n_8537)
);

NAND2xp5_ASAP7_75t_L g8538 ( 
.A(n_7803),
.B(n_6954),
.Y(n_8538)
);

NAND2xp33_ASAP7_75t_L g8539 ( 
.A(n_8212),
.B(n_7719),
.Y(n_8539)
);

NOR3xp33_ASAP7_75t_L g8540 ( 
.A(n_8347),
.B(n_8370),
.C(n_8154),
.Y(n_8540)
);

NAND2xp5_ASAP7_75t_SL g8541 ( 
.A(n_8212),
.B(n_7712),
.Y(n_8541)
);

NOR2x1p5_ASAP7_75t_L g8542 ( 
.A(n_7805),
.B(n_7678),
.Y(n_8542)
);

A2O1A1Ixp33_ASAP7_75t_L g8543 ( 
.A1(n_8057),
.A2(n_7673),
.B(n_7003),
.C(n_6991),
.Y(n_8543)
);

NOR2xp33_ASAP7_75t_L g8544 ( 
.A(n_7842),
.B(n_7725),
.Y(n_8544)
);

O2A1O1Ixp33_ASAP7_75t_L g8545 ( 
.A1(n_8361),
.A2(n_7704),
.B(n_7056),
.C(n_7323),
.Y(n_8545)
);

INVx3_ASAP7_75t_L g8546 ( 
.A(n_8066),
.Y(n_8546)
);

NAND2xp5_ASAP7_75t_L g8547 ( 
.A(n_7917),
.B(n_7727),
.Y(n_8547)
);

NOR2xp33_ASAP7_75t_L g8548 ( 
.A(n_7775),
.B(n_7526),
.Y(n_8548)
);

NOR2xp33_ASAP7_75t_L g8549 ( 
.A(n_7783),
.B(n_7526),
.Y(n_8549)
);

NOR2xp33_ASAP7_75t_L g8550 ( 
.A(n_7975),
.B(n_7434),
.Y(n_8550)
);

NOR2xp33_ASAP7_75t_L g8551 ( 
.A(n_7976),
.B(n_7485),
.Y(n_8551)
);

INVx1_ASAP7_75t_L g8552 ( 
.A(n_7770),
.Y(n_8552)
);

AND2x2_ASAP7_75t_L g8553 ( 
.A(n_7831),
.B(n_7217),
.Y(n_8553)
);

NAND2xp5_ASAP7_75t_L g8554 ( 
.A(n_7853),
.B(n_7370),
.Y(n_8554)
);

NAND2xp5_ASAP7_75t_L g8555 ( 
.A(n_7792),
.B(n_7606),
.Y(n_8555)
);

INVx1_ASAP7_75t_L g8556 ( 
.A(n_7777),
.Y(n_8556)
);

INVx2_ASAP7_75t_L g8557 ( 
.A(n_7984),
.Y(n_8557)
);

NAND2xp5_ASAP7_75t_SL g8558 ( 
.A(n_8212),
.B(n_7265),
.Y(n_8558)
);

INVx2_ASAP7_75t_L g8559 ( 
.A(n_7987),
.Y(n_8559)
);

NOR2xp33_ASAP7_75t_L g8560 ( 
.A(n_7784),
.B(n_7078),
.Y(n_8560)
);

NAND2xp5_ASAP7_75t_L g8561 ( 
.A(n_7810),
.B(n_7437),
.Y(n_8561)
);

NAND2xp5_ASAP7_75t_SL g8562 ( 
.A(n_8277),
.B(n_7064),
.Y(n_8562)
);

NAND2xp5_ASAP7_75t_SL g8563 ( 
.A(n_8277),
.B(n_7067),
.Y(n_8563)
);

NOR2xp33_ASAP7_75t_L g8564 ( 
.A(n_8039),
.B(n_7295),
.Y(n_8564)
);

NAND2xp5_ASAP7_75t_L g8565 ( 
.A(n_7843),
.B(n_7301),
.Y(n_8565)
);

INVx1_ASAP7_75t_L g8566 ( 
.A(n_7779),
.Y(n_8566)
);

INVx1_ASAP7_75t_L g8567 ( 
.A(n_7782),
.Y(n_8567)
);

NAND2xp5_ASAP7_75t_L g8568 ( 
.A(n_7861),
.B(n_7487),
.Y(n_8568)
);

INVx2_ASAP7_75t_L g8569 ( 
.A(n_7991),
.Y(n_8569)
);

NAND2xp5_ASAP7_75t_SL g8570 ( 
.A(n_8277),
.B(n_7492),
.Y(n_8570)
);

NOR2xp33_ASAP7_75t_R g8571 ( 
.A(n_7817),
.B(n_2474),
.Y(n_8571)
);

NOR2xp33_ASAP7_75t_L g8572 ( 
.A(n_8248),
.B(n_7663),
.Y(n_8572)
);

INVx1_ASAP7_75t_L g8573 ( 
.A(n_7785),
.Y(n_8573)
);

INVx1_ASAP7_75t_L g8574 ( 
.A(n_7787),
.Y(n_8574)
);

BUFx2_ASAP7_75t_L g8575 ( 
.A(n_8158),
.Y(n_8575)
);

NAND2xp5_ASAP7_75t_L g8576 ( 
.A(n_7870),
.B(n_7690),
.Y(n_8576)
);

INVx2_ASAP7_75t_L g8577 ( 
.A(n_7995),
.Y(n_8577)
);

NAND2xp5_ASAP7_75t_L g8578 ( 
.A(n_7873),
.B(n_7202),
.Y(n_8578)
);

INVx2_ASAP7_75t_L g8579 ( 
.A(n_7996),
.Y(n_8579)
);

OR2x6_ASAP7_75t_L g8580 ( 
.A(n_8053),
.B(n_34),
.Y(n_8580)
);

INVx1_ASAP7_75t_L g8581 ( 
.A(n_7788),
.Y(n_8581)
);

NAND2xp5_ASAP7_75t_L g8582 ( 
.A(n_7795),
.B(n_34),
.Y(n_8582)
);

NAND2xp5_ASAP7_75t_L g8583 ( 
.A(n_7944),
.B(n_34),
.Y(n_8583)
);

INVx2_ASAP7_75t_L g8584 ( 
.A(n_8218),
.Y(n_8584)
);

AND2x6_ASAP7_75t_SL g8585 ( 
.A(n_7839),
.B(n_35),
.Y(n_8585)
);

NOR2x1p5_ASAP7_75t_L g8586 ( 
.A(n_8137),
.B(n_2475),
.Y(n_8586)
);

AND2x2_ASAP7_75t_L g8587 ( 
.A(n_7966),
.B(n_2476),
.Y(n_8587)
);

NAND2xp5_ASAP7_75t_L g8588 ( 
.A(n_7963),
.B(n_7964),
.Y(n_8588)
);

NAND2xp5_ASAP7_75t_SL g8589 ( 
.A(n_8277),
.B(n_8252),
.Y(n_8589)
);

INVx1_ASAP7_75t_L g8590 ( 
.A(n_7790),
.Y(n_8590)
);

NAND2xp5_ASAP7_75t_L g8591 ( 
.A(n_7985),
.B(n_35),
.Y(n_8591)
);

INVx2_ASAP7_75t_L g8592 ( 
.A(n_8219),
.Y(n_8592)
);

NOR2xp33_ASAP7_75t_L g8593 ( 
.A(n_8156),
.B(n_2476),
.Y(n_8593)
);

NAND2xp5_ASAP7_75t_L g8594 ( 
.A(n_7990),
.B(n_8004),
.Y(n_8594)
);

AOI22xp5_ASAP7_75t_L g8595 ( 
.A1(n_8107),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_8595)
);

BUFx3_ASAP7_75t_L g8596 ( 
.A(n_8084),
.Y(n_8596)
);

INVx1_ASAP7_75t_L g8597 ( 
.A(n_7791),
.Y(n_8597)
);

CKINVDCx5p33_ASAP7_75t_R g8598 ( 
.A(n_7905),
.Y(n_8598)
);

INVx2_ASAP7_75t_L g8599 ( 
.A(n_8220),
.Y(n_8599)
);

INVx2_ASAP7_75t_L g8600 ( 
.A(n_8215),
.Y(n_8600)
);

NOR2xp67_ASAP7_75t_SL g8601 ( 
.A(n_7737),
.B(n_2477),
.Y(n_8601)
);

NOR2xp67_ASAP7_75t_L g8602 ( 
.A(n_7741),
.B(n_36),
.Y(n_8602)
);

INVx1_ASAP7_75t_L g8603 ( 
.A(n_7794),
.Y(n_8603)
);

AND2x6_ASAP7_75t_L g8604 ( 
.A(n_8124),
.B(n_36),
.Y(n_8604)
);

OAI22xp5_ASAP7_75t_L g8605 ( 
.A1(n_7793),
.A2(n_2478),
.B1(n_2479),
.B2(n_2477),
.Y(n_8605)
);

NAND2xp5_ASAP7_75t_L g8606 ( 
.A(n_8038),
.B(n_38),
.Y(n_8606)
);

NAND2xp5_ASAP7_75t_SL g8607 ( 
.A(n_7898),
.B(n_8351),
.Y(n_8607)
);

NAND2xp5_ASAP7_75t_L g8608 ( 
.A(n_7969),
.B(n_38),
.Y(n_8608)
);

NOR2xp33_ASAP7_75t_L g8609 ( 
.A(n_8253),
.B(n_2480),
.Y(n_8609)
);

AOI22xp33_ASAP7_75t_L g8610 ( 
.A1(n_7771),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_8610)
);

INVx1_ASAP7_75t_L g8611 ( 
.A(n_7796),
.Y(n_8611)
);

INVx1_ASAP7_75t_L g8612 ( 
.A(n_7797),
.Y(n_8612)
);

AND2x2_ASAP7_75t_L g8613 ( 
.A(n_8195),
.B(n_2480),
.Y(n_8613)
);

NAND2xp5_ASAP7_75t_SL g8614 ( 
.A(n_7816),
.B(n_2482),
.Y(n_8614)
);

NAND2xp5_ASAP7_75t_L g8615 ( 
.A(n_7841),
.B(n_39),
.Y(n_8615)
);

A2O1A1Ixp33_ASAP7_75t_L g8616 ( 
.A1(n_8062),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_8616)
);

INVx1_ASAP7_75t_L g8617 ( 
.A(n_7798),
.Y(n_8617)
);

AND2x2_ASAP7_75t_L g8618 ( 
.A(n_8380),
.B(n_2483),
.Y(n_8618)
);

NOR2xp67_ASAP7_75t_L g8619 ( 
.A(n_8357),
.B(n_41),
.Y(n_8619)
);

AND2x2_ASAP7_75t_SL g8620 ( 
.A(n_8082),
.B(n_41),
.Y(n_8620)
);

NAND2xp33_ASAP7_75t_L g8621 ( 
.A(n_7824),
.B(n_2484),
.Y(n_8621)
);

BUFx3_ASAP7_75t_L g8622 ( 
.A(n_8091),
.Y(n_8622)
);

NAND2xp5_ASAP7_75t_SL g8623 ( 
.A(n_8330),
.B(n_2484),
.Y(n_8623)
);

NAND2xp5_ASAP7_75t_L g8624 ( 
.A(n_7841),
.B(n_42),
.Y(n_8624)
);

AOI22xp33_ASAP7_75t_L g8625 ( 
.A1(n_8042),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_8625)
);

NOR2xp33_ASAP7_75t_L g8626 ( 
.A(n_8282),
.B(n_2485),
.Y(n_8626)
);

NAND2xp5_ASAP7_75t_SL g8627 ( 
.A(n_8329),
.B(n_2487),
.Y(n_8627)
);

NAND2xp5_ASAP7_75t_L g8628 ( 
.A(n_7841),
.B(n_43),
.Y(n_8628)
);

NAND2xp5_ASAP7_75t_L g8629 ( 
.A(n_7970),
.B(n_44),
.Y(n_8629)
);

NAND2xp5_ASAP7_75t_L g8630 ( 
.A(n_7914),
.B(n_44),
.Y(n_8630)
);

NAND2xp5_ASAP7_75t_L g8631 ( 
.A(n_7925),
.B(n_45),
.Y(n_8631)
);

OAI22xp5_ASAP7_75t_L g8632 ( 
.A1(n_8348),
.A2(n_2488),
.B1(n_2489),
.B2(n_2487),
.Y(n_8632)
);

AOI22xp33_ASAP7_75t_L g8633 ( 
.A1(n_8398),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_8633)
);

XOR2x2_ASAP7_75t_L g8634 ( 
.A(n_7767),
.B(n_46),
.Y(n_8634)
);

NAND2xp5_ASAP7_75t_L g8635 ( 
.A(n_7903),
.B(n_47),
.Y(n_8635)
);

NOR2xp33_ASAP7_75t_L g8636 ( 
.A(n_8319),
.B(n_2488),
.Y(n_8636)
);

NAND2xp5_ASAP7_75t_L g8637 ( 
.A(n_7929),
.B(n_48),
.Y(n_8637)
);

NAND3xp33_ASAP7_75t_L g8638 ( 
.A(n_8393),
.B(n_48),
.C(n_49),
.Y(n_8638)
);

NOR2xp67_ASAP7_75t_L g8639 ( 
.A(n_8122),
.B(n_8132),
.Y(n_8639)
);

NAND2xp5_ASAP7_75t_L g8640 ( 
.A(n_7932),
.B(n_7801),
.Y(n_8640)
);

NAND2xp5_ASAP7_75t_L g8641 ( 
.A(n_7942),
.B(n_49),
.Y(n_8641)
);

NAND2xp5_ASAP7_75t_L g8642 ( 
.A(n_7800),
.B(n_50),
.Y(n_8642)
);

INVx1_ASAP7_75t_L g8643 ( 
.A(n_7799),
.Y(n_8643)
);

INVx2_ASAP7_75t_SL g8644 ( 
.A(n_7780),
.Y(n_8644)
);

NAND2xp5_ASAP7_75t_L g8645 ( 
.A(n_7802),
.B(n_50),
.Y(n_8645)
);

INVx3_ASAP7_75t_L g8646 ( 
.A(n_7780),
.Y(n_8646)
);

INVxp67_ASAP7_75t_L g8647 ( 
.A(n_8379),
.Y(n_8647)
);

NOR2xp33_ASAP7_75t_L g8648 ( 
.A(n_7866),
.B(n_2490),
.Y(n_8648)
);

O2A1O1Ixp5_ASAP7_75t_L g8649 ( 
.A1(n_8146),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_8649)
);

AOI21xp5_ASAP7_75t_L g8650 ( 
.A1(n_7948),
.A2(n_2491),
.B(n_2490),
.Y(n_8650)
);

BUFx3_ASAP7_75t_L g8651 ( 
.A(n_8072),
.Y(n_8651)
);

NAND2xp5_ASAP7_75t_L g8652 ( 
.A(n_7804),
.B(n_51),
.Y(n_8652)
);

INVx2_ASAP7_75t_L g8653 ( 
.A(n_8006),
.Y(n_8653)
);

BUFx4f_ASAP7_75t_L g8654 ( 
.A(n_7871),
.Y(n_8654)
);

INVx2_ASAP7_75t_L g8655 ( 
.A(n_8008),
.Y(n_8655)
);

INVx1_ASAP7_75t_L g8656 ( 
.A(n_7807),
.Y(n_8656)
);

NOR2xp33_ASAP7_75t_L g8657 ( 
.A(n_8239),
.B(n_8001),
.Y(n_8657)
);

NAND2xp5_ASAP7_75t_SL g8658 ( 
.A(n_7992),
.B(n_2491),
.Y(n_8658)
);

NAND2xp5_ASAP7_75t_L g8659 ( 
.A(n_7809),
.B(n_51),
.Y(n_8659)
);

NOR2xp33_ASAP7_75t_L g8660 ( 
.A(n_8005),
.B(n_2492),
.Y(n_8660)
);

OAI221xp5_ASAP7_75t_L g8661 ( 
.A1(n_8052),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.C(n_55),
.Y(n_8661)
);

NAND2xp5_ASAP7_75t_L g8662 ( 
.A(n_7812),
.B(n_54),
.Y(n_8662)
);

NAND2xp5_ASAP7_75t_L g8663 ( 
.A(n_7813),
.B(n_54),
.Y(n_8663)
);

NAND2xp5_ASAP7_75t_L g8664 ( 
.A(n_7814),
.B(n_55),
.Y(n_8664)
);

INVx1_ASAP7_75t_L g8665 ( 
.A(n_7815),
.Y(n_8665)
);

NOR2xp33_ASAP7_75t_L g8666 ( 
.A(n_8012),
.B(n_2492),
.Y(n_8666)
);

NAND2xp33_ASAP7_75t_SL g8667 ( 
.A(n_8050),
.B(n_2493),
.Y(n_8667)
);

O2A1O1Ixp33_ASAP7_75t_L g8668 ( 
.A1(n_8304),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_8668)
);

NAND2xp5_ASAP7_75t_SL g8669 ( 
.A(n_7824),
.B(n_2494),
.Y(n_8669)
);

INVx1_ASAP7_75t_L g8670 ( 
.A(n_7818),
.Y(n_8670)
);

INVx2_ASAP7_75t_SL g8671 ( 
.A(n_7871),
.Y(n_8671)
);

NOR3xp33_ASAP7_75t_L g8672 ( 
.A(n_8271),
.B(n_56),
.C(n_57),
.Y(n_8672)
);

INVx2_ASAP7_75t_L g8673 ( 
.A(n_8010),
.Y(n_8673)
);

NAND2xp5_ASAP7_75t_L g8674 ( 
.A(n_7825),
.B(n_56),
.Y(n_8674)
);

OAI22xp5_ASAP7_75t_L g8675 ( 
.A1(n_8246),
.A2(n_2496),
.B1(n_2498),
.B2(n_2495),
.Y(n_8675)
);

NOR2xp33_ASAP7_75t_L g8676 ( 
.A(n_8073),
.B(n_2495),
.Y(n_8676)
);

INVx3_ASAP7_75t_L g8677 ( 
.A(n_7928),
.Y(n_8677)
);

NAND2xp5_ASAP7_75t_SL g8678 ( 
.A(n_7824),
.B(n_2496),
.Y(n_8678)
);

NOR3xp33_ASAP7_75t_L g8679 ( 
.A(n_8075),
.B(n_57),
.C(n_58),
.Y(n_8679)
);

INVx2_ASAP7_75t_L g8680 ( 
.A(n_8017),
.Y(n_8680)
);

NOR2xp33_ASAP7_75t_L g8681 ( 
.A(n_8127),
.B(n_2499),
.Y(n_8681)
);

INVx2_ASAP7_75t_L g8682 ( 
.A(n_8018),
.Y(n_8682)
);

NOR2xp67_ASAP7_75t_L g8683 ( 
.A(n_8307),
.B(n_8371),
.Y(n_8683)
);

INVx1_ASAP7_75t_L g8684 ( 
.A(n_7827),
.Y(n_8684)
);

NOR2xp33_ASAP7_75t_SL g8685 ( 
.A(n_7811),
.B(n_58),
.Y(n_8685)
);

INVx2_ASAP7_75t_SL g8686 ( 
.A(n_7928),
.Y(n_8686)
);

NAND2xp5_ASAP7_75t_SL g8687 ( 
.A(n_7824),
.B(n_2500),
.Y(n_8687)
);

NAND2xp5_ASAP7_75t_L g8688 ( 
.A(n_7833),
.B(n_59),
.Y(n_8688)
);

INVx2_ASAP7_75t_L g8689 ( 
.A(n_8021),
.Y(n_8689)
);

NAND2xp5_ASAP7_75t_L g8690 ( 
.A(n_7835),
.B(n_7836),
.Y(n_8690)
);

NAND2xp5_ASAP7_75t_SL g8691 ( 
.A(n_7830),
.B(n_2500),
.Y(n_8691)
);

NAND2xp5_ASAP7_75t_L g8692 ( 
.A(n_7837),
.B(n_59),
.Y(n_8692)
);

BUFx6f_ASAP7_75t_SL g8693 ( 
.A(n_7999),
.Y(n_8693)
);

NAND2xp5_ASAP7_75t_SL g8694 ( 
.A(n_7830),
.B(n_2501),
.Y(n_8694)
);

OAI22xp33_ASAP7_75t_L g8695 ( 
.A1(n_8175),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_8695)
);

NAND2xp5_ASAP7_75t_SL g8696 ( 
.A(n_7830),
.B(n_2502),
.Y(n_8696)
);

OR2x2_ASAP7_75t_L g8697 ( 
.A(n_8287),
.B(n_60),
.Y(n_8697)
);

NAND2xp5_ASAP7_75t_L g8698 ( 
.A(n_7840),
.B(n_60),
.Y(n_8698)
);

NAND2xp5_ASAP7_75t_L g8699 ( 
.A(n_7845),
.B(n_61),
.Y(n_8699)
);

INVx8_ASAP7_75t_L g8700 ( 
.A(n_7851),
.Y(n_8700)
);

NOR2xp33_ASAP7_75t_L g8701 ( 
.A(n_8129),
.B(n_2502),
.Y(n_8701)
);

INVx4_ASAP7_75t_L g8702 ( 
.A(n_8164),
.Y(n_8702)
);

NOR3xp33_ASAP7_75t_L g8703 ( 
.A(n_8090),
.B(n_61),
.C(n_62),
.Y(n_8703)
);

NAND2xp5_ASAP7_75t_L g8704 ( 
.A(n_7847),
.B(n_62),
.Y(n_8704)
);

NOR2x1p5_ASAP7_75t_L g8705 ( 
.A(n_8030),
.B(n_2503),
.Y(n_8705)
);

INVx1_ASAP7_75t_L g8706 ( 
.A(n_7849),
.Y(n_8706)
);

NOR2xp33_ASAP7_75t_L g8707 ( 
.A(n_8147),
.B(n_2504),
.Y(n_8707)
);

NAND2xp5_ASAP7_75t_SL g8708 ( 
.A(n_7830),
.B(n_2506),
.Y(n_8708)
);

OAI21xp5_ASAP7_75t_L g8709 ( 
.A1(n_7949),
.A2(n_8293),
.B(n_8275),
.Y(n_8709)
);

OAI22xp33_ASAP7_75t_L g8710 ( 
.A1(n_7896),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_8710)
);

OAI22xp5_ASAP7_75t_L g8711 ( 
.A1(n_8324),
.A2(n_2507),
.B1(n_2508),
.B2(n_2506),
.Y(n_8711)
);

NAND2xp5_ASAP7_75t_SL g8712 ( 
.A(n_8069),
.B(n_2508),
.Y(n_8712)
);

NOR2xp33_ASAP7_75t_L g8713 ( 
.A(n_8261),
.B(n_2509),
.Y(n_8713)
);

AND2x2_ASAP7_75t_L g8714 ( 
.A(n_8223),
.B(n_2509),
.Y(n_8714)
);

INVx1_ASAP7_75t_L g8715 ( 
.A(n_7850),
.Y(n_8715)
);

NOR2xp33_ASAP7_75t_L g8716 ( 
.A(n_8170),
.B(n_2510),
.Y(n_8716)
);

NAND2xp5_ASAP7_75t_L g8717 ( 
.A(n_7852),
.B(n_63),
.Y(n_8717)
);

NAND2xp5_ASAP7_75t_SL g8718 ( 
.A(n_8069),
.B(n_2510),
.Y(n_8718)
);

NAND2xp5_ASAP7_75t_SL g8719 ( 
.A(n_8069),
.B(n_2511),
.Y(n_8719)
);

NAND2xp5_ASAP7_75t_SL g8720 ( 
.A(n_8069),
.B(n_2511),
.Y(n_8720)
);

INVx2_ASAP7_75t_L g8721 ( 
.A(n_8022),
.Y(n_8721)
);

NOR2xp33_ASAP7_75t_L g8722 ( 
.A(n_8170),
.B(n_2513),
.Y(n_8722)
);

INVx2_ASAP7_75t_L g8723 ( 
.A(n_8023),
.Y(n_8723)
);

INVx1_ASAP7_75t_L g8724 ( 
.A(n_7854),
.Y(n_8724)
);

NAND2xp5_ASAP7_75t_L g8725 ( 
.A(n_7856),
.B(n_64),
.Y(n_8725)
);

NAND2xp5_ASAP7_75t_L g8726 ( 
.A(n_7857),
.B(n_7858),
.Y(n_8726)
);

OAI22xp5_ASAP7_75t_L g8727 ( 
.A1(n_8292),
.A2(n_2515),
.B1(n_2516),
.B2(n_2513),
.Y(n_8727)
);

NAND2xp5_ASAP7_75t_L g8728 ( 
.A(n_7862),
.B(n_64),
.Y(n_8728)
);

AOI21xp5_ASAP7_75t_L g8729 ( 
.A1(n_8301),
.A2(n_2517),
.B(n_2516),
.Y(n_8729)
);

NAND2xp5_ASAP7_75t_L g8730 ( 
.A(n_7864),
.B(n_7867),
.Y(n_8730)
);

AND2x2_ASAP7_75t_L g8731 ( 
.A(n_8300),
.B(n_2517),
.Y(n_8731)
);

INVx2_ASAP7_75t_L g8732 ( 
.A(n_8025),
.Y(n_8732)
);

AO22x1_ASAP7_75t_L g8733 ( 
.A1(n_8102),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_8733)
);

NAND2xp5_ASAP7_75t_L g8734 ( 
.A(n_7868),
.B(n_65),
.Y(n_8734)
);

INVx2_ASAP7_75t_SL g8735 ( 
.A(n_7974),
.Y(n_8735)
);

NAND2xp5_ASAP7_75t_L g8736 ( 
.A(n_7869),
.B(n_66),
.Y(n_8736)
);

AND2x2_ASAP7_75t_L g8737 ( 
.A(n_8318),
.B(n_2518),
.Y(n_8737)
);

INVx1_ASAP7_75t_L g8738 ( 
.A(n_7875),
.Y(n_8738)
);

INVx1_ASAP7_75t_L g8739 ( 
.A(n_7877),
.Y(n_8739)
);

INVx1_ASAP7_75t_L g8740 ( 
.A(n_7881),
.Y(n_8740)
);

INVx1_ASAP7_75t_L g8741 ( 
.A(n_7883),
.Y(n_8741)
);

NAND2xp5_ASAP7_75t_SL g8742 ( 
.A(n_8224),
.B(n_7832),
.Y(n_8742)
);

INVx1_ASAP7_75t_L g8743 ( 
.A(n_7887),
.Y(n_8743)
);

INVx2_ASAP7_75t_SL g8744 ( 
.A(n_7974),
.Y(n_8744)
);

NAND2xp5_ASAP7_75t_L g8745 ( 
.A(n_7888),
.B(n_67),
.Y(n_8745)
);

INVx2_ASAP7_75t_L g8746 ( 
.A(n_8037),
.Y(n_8746)
);

AOI22xp33_ASAP7_75t_L g8747 ( 
.A1(n_8400),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_8747)
);

NAND2xp5_ASAP7_75t_L g8748 ( 
.A(n_7889),
.B(n_7890),
.Y(n_8748)
);

BUFx5_ASAP7_75t_L g8749 ( 
.A(n_8141),
.Y(n_8749)
);

INVx2_ASAP7_75t_SL g8750 ( 
.A(n_7986),
.Y(n_8750)
);

NAND3xp33_ASAP7_75t_L g8751 ( 
.A(n_8130),
.B(n_68),
.C(n_69),
.Y(n_8751)
);

INVx3_ASAP7_75t_L g8752 ( 
.A(n_7986),
.Y(n_8752)
);

NAND2xp5_ASAP7_75t_L g8753 ( 
.A(n_7891),
.B(n_68),
.Y(n_8753)
);

INVx2_ASAP7_75t_SL g8754 ( 
.A(n_8054),
.Y(n_8754)
);

NAND2xp5_ASAP7_75t_SL g8755 ( 
.A(n_8294),
.B(n_2518),
.Y(n_8755)
);

AND2x2_ASAP7_75t_L g8756 ( 
.A(n_8333),
.B(n_2519),
.Y(n_8756)
);

O2A1O1Ixp33_ASAP7_75t_L g8757 ( 
.A1(n_8171),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_8757)
);

NAND2xp5_ASAP7_75t_SL g8758 ( 
.A(n_8311),
.B(n_2519),
.Y(n_8758)
);

BUFx6f_ASAP7_75t_L g8759 ( 
.A(n_8054),
.Y(n_8759)
);

INVx1_ASAP7_75t_L g8760 ( 
.A(n_7893),
.Y(n_8760)
);

NAND2xp5_ASAP7_75t_L g8761 ( 
.A(n_7894),
.B(n_71),
.Y(n_8761)
);

INVx2_ASAP7_75t_L g8762 ( 
.A(n_8056),
.Y(n_8762)
);

CKINVDCx5p33_ASAP7_75t_R g8763 ( 
.A(n_7879),
.Y(n_8763)
);

INVx1_ASAP7_75t_L g8764 ( 
.A(n_7895),
.Y(n_8764)
);

OAI22xp5_ASAP7_75t_L g8765 ( 
.A1(n_8383),
.A2(n_8394),
.B1(n_8399),
.B2(n_8397),
.Y(n_8765)
);

NAND2xp5_ASAP7_75t_L g8766 ( 
.A(n_7899),
.B(n_71),
.Y(n_8766)
);

AND2x2_ASAP7_75t_SL g8767 ( 
.A(n_8285),
.B(n_72),
.Y(n_8767)
);

AOI22xp5_ASAP7_75t_L g8768 ( 
.A1(n_8213),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_8768)
);

NAND2xp5_ASAP7_75t_L g8769 ( 
.A(n_7900),
.B(n_73),
.Y(n_8769)
);

NOR3xp33_ASAP7_75t_L g8770 ( 
.A(n_8269),
.B(n_73),
.C(n_74),
.Y(n_8770)
);

OAI21xp5_ASAP7_75t_L g8771 ( 
.A1(n_7776),
.A2(n_74),
.B(n_76),
.Y(n_8771)
);

NAND2xp5_ASAP7_75t_L g8772 ( 
.A(n_7901),
.B(n_76),
.Y(n_8772)
);

NAND2xp5_ASAP7_75t_L g8773 ( 
.A(n_7902),
.B(n_77),
.Y(n_8773)
);

NAND2xp5_ASAP7_75t_SL g8774 ( 
.A(n_8134),
.B(n_2520),
.Y(n_8774)
);

INVxp67_ASAP7_75t_L g8775 ( 
.A(n_8134),
.Y(n_8775)
);

NAND2xp5_ASAP7_75t_SL g8776 ( 
.A(n_8155),
.B(n_2522),
.Y(n_8776)
);

NOR2x1p5_ASAP7_75t_L g8777 ( 
.A(n_8180),
.B(n_2524),
.Y(n_8777)
);

NAND2xp5_ASAP7_75t_L g8778 ( 
.A(n_7906),
.B(n_77),
.Y(n_8778)
);

INVx1_ASAP7_75t_L g8779 ( 
.A(n_7907),
.Y(n_8779)
);

OAI22xp5_ASAP7_75t_L g8780 ( 
.A1(n_8401),
.A2(n_2525),
.B1(n_2526),
.B2(n_2524),
.Y(n_8780)
);

AOI22xp5_ASAP7_75t_L g8781 ( 
.A1(n_8327),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_8781)
);

AOI22xp5_ASAP7_75t_L g8782 ( 
.A1(n_8402),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_8782)
);

AOI22xp5_ASAP7_75t_L g8783 ( 
.A1(n_8408),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_8783)
);

NAND2xp5_ASAP7_75t_SL g8784 ( 
.A(n_8155),
.B(n_2525),
.Y(n_8784)
);

NOR2xp33_ASAP7_75t_L g8785 ( 
.A(n_8395),
.B(n_2527),
.Y(n_8785)
);

NOR3xp33_ASAP7_75t_L g8786 ( 
.A(n_8310),
.B(n_80),
.C(n_81),
.Y(n_8786)
);

AOI21xp5_ASAP7_75t_L g8787 ( 
.A1(n_8065),
.A2(n_2531),
.B(n_2527),
.Y(n_8787)
);

NAND2xp5_ASAP7_75t_L g8788 ( 
.A(n_7910),
.B(n_7911),
.Y(n_8788)
);

INVx1_ASAP7_75t_L g8789 ( 
.A(n_7913),
.Y(n_8789)
);

INVxp67_ASAP7_75t_L g8790 ( 
.A(n_8267),
.Y(n_8790)
);

NAND2xp5_ASAP7_75t_L g8791 ( 
.A(n_7915),
.B(n_81),
.Y(n_8791)
);

INVx1_ASAP7_75t_L g8792 ( 
.A(n_7919),
.Y(n_8792)
);

AOI22xp5_ASAP7_75t_L g8793 ( 
.A1(n_8337),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_8793)
);

NOR2xp33_ASAP7_75t_L g8794 ( 
.A(n_8267),
.B(n_2531),
.Y(n_8794)
);

NAND2xp5_ASAP7_75t_SL g8795 ( 
.A(n_8295),
.B(n_2532),
.Y(n_8795)
);

NAND2xp5_ASAP7_75t_L g8796 ( 
.A(n_7920),
.B(n_83),
.Y(n_8796)
);

NAND2xp5_ASAP7_75t_L g8797 ( 
.A(n_7922),
.B(n_83),
.Y(n_8797)
);

AND2x2_ASAP7_75t_L g8798 ( 
.A(n_8365),
.B(n_2533),
.Y(n_8798)
);

OAI22xp5_ASAP7_75t_L g8799 ( 
.A1(n_8403),
.A2(n_8406),
.B1(n_8409),
.B2(n_8404),
.Y(n_8799)
);

AOI22xp5_ASAP7_75t_L g8800 ( 
.A1(n_8290),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_8800)
);

OR2x2_ASAP7_75t_L g8801 ( 
.A(n_8368),
.B(n_84),
.Y(n_8801)
);

NAND2xp5_ASAP7_75t_L g8802 ( 
.A(n_7923),
.B(n_85),
.Y(n_8802)
);

NAND2xp5_ASAP7_75t_L g8803 ( 
.A(n_7924),
.B(n_85),
.Y(n_8803)
);

INVx1_ASAP7_75t_L g8804 ( 
.A(n_7926),
.Y(n_8804)
);

NAND2xp5_ASAP7_75t_L g8805 ( 
.A(n_7927),
.B(n_86),
.Y(n_8805)
);

INVx6_ASAP7_75t_L g8806 ( 
.A(n_8128),
.Y(n_8806)
);

INVx1_ASAP7_75t_L g8807 ( 
.A(n_7933),
.Y(n_8807)
);

NAND2xp5_ASAP7_75t_L g8808 ( 
.A(n_7934),
.B(n_87),
.Y(n_8808)
);

NAND2xp5_ASAP7_75t_L g8809 ( 
.A(n_7937),
.B(n_87),
.Y(n_8809)
);

NAND2xp5_ASAP7_75t_SL g8810 ( 
.A(n_8295),
.B(n_7846),
.Y(n_8810)
);

AND2x2_ASAP7_75t_L g8811 ( 
.A(n_8240),
.B(n_2533),
.Y(n_8811)
);

INVx2_ASAP7_75t_L g8812 ( 
.A(n_8059),
.Y(n_8812)
);

NAND2xp5_ASAP7_75t_L g8813 ( 
.A(n_7938),
.B(n_7943),
.Y(n_8813)
);

AND2x4_ASAP7_75t_L g8814 ( 
.A(n_8034),
.B(n_8080),
.Y(n_8814)
);

OAI22xp5_ASAP7_75t_L g8815 ( 
.A1(n_8186),
.A2(n_2535),
.B1(n_2536),
.B2(n_2534),
.Y(n_8815)
);

INVx1_ASAP7_75t_L g8816 ( 
.A(n_7945),
.Y(n_8816)
);

NAND2xp5_ASAP7_75t_L g8817 ( 
.A(n_7947),
.B(n_88),
.Y(n_8817)
);

AO221x1_ASAP7_75t_L g8818 ( 
.A1(n_8159),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.C(n_91),
.Y(n_8818)
);

NOR2xp33_ASAP7_75t_L g8819 ( 
.A(n_8384),
.B(n_2535),
.Y(n_8819)
);

NAND2xp5_ASAP7_75t_SL g8820 ( 
.A(n_7909),
.B(n_2537),
.Y(n_8820)
);

INVx1_ASAP7_75t_L g8821 ( 
.A(n_7952),
.Y(n_8821)
);

AOI22xp5_ASAP7_75t_L g8822 ( 
.A1(n_8227),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_8822)
);

AND2x6_ASAP7_75t_SL g8823 ( 
.A(n_7886),
.B(n_90),
.Y(n_8823)
);

INVxp67_ASAP7_75t_L g8824 ( 
.A(n_8237),
.Y(n_8824)
);

NAND2xp5_ASAP7_75t_SL g8825 ( 
.A(n_7946),
.B(n_2537),
.Y(n_8825)
);

NAND3xp33_ASAP7_75t_SL g8826 ( 
.A(n_7930),
.B(n_91),
.C(n_92),
.Y(n_8826)
);

OAI22xp33_ASAP7_75t_L g8827 ( 
.A1(n_7967),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_8827)
);

NAND2xp5_ASAP7_75t_SL g8828 ( 
.A(n_8321),
.B(n_2538),
.Y(n_8828)
);

INVxp67_ASAP7_75t_L g8829 ( 
.A(n_8308),
.Y(n_8829)
);

INVx2_ASAP7_75t_L g8830 ( 
.A(n_8068),
.Y(n_8830)
);

NOR2xp33_ASAP7_75t_L g8831 ( 
.A(n_8385),
.B(n_2538),
.Y(n_8831)
);

NAND2xp5_ASAP7_75t_L g8832 ( 
.A(n_7953),
.B(n_93),
.Y(n_8832)
);

NOR2xp33_ASAP7_75t_L g8833 ( 
.A(n_8387),
.B(n_2539),
.Y(n_8833)
);

INVxp67_ASAP7_75t_SL g8834 ( 
.A(n_8205),
.Y(n_8834)
);

NAND2xp5_ASAP7_75t_SL g8835 ( 
.A(n_8321),
.B(n_2540),
.Y(n_8835)
);

NAND2xp5_ASAP7_75t_L g8836 ( 
.A(n_7981),
.B(n_93),
.Y(n_8836)
);

NOR2xp33_ASAP7_75t_L g8837 ( 
.A(n_8388),
.B(n_2541),
.Y(n_8837)
);

INVx1_ASAP7_75t_L g8838 ( 
.A(n_8157),
.Y(n_8838)
);

AND2x4_ASAP7_75t_L g8839 ( 
.A(n_8128),
.B(n_94),
.Y(n_8839)
);

NOR2xp33_ASAP7_75t_L g8840 ( 
.A(n_7997),
.B(n_2543),
.Y(n_8840)
);

NOR2x1p5_ASAP7_75t_L g8841 ( 
.A(n_8185),
.B(n_2543),
.Y(n_8841)
);

NOR2xp33_ASAP7_75t_L g8842 ( 
.A(n_7956),
.B(n_2545),
.Y(n_8842)
);

NAND2xp5_ASAP7_75t_L g8843 ( 
.A(n_8032),
.B(n_94),
.Y(n_8843)
);

AOI22xp5_ASAP7_75t_L g8844 ( 
.A1(n_7983),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_8844)
);

BUFx3_ASAP7_75t_L g8845 ( 
.A(n_7954),
.Y(n_8845)
);

AOI22xp5_ASAP7_75t_L g8846 ( 
.A1(n_8373),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_8846)
);

INVx2_ASAP7_75t_L g8847 ( 
.A(n_8076),
.Y(n_8847)
);

INVxp67_ASAP7_75t_SL g8848 ( 
.A(n_8207),
.Y(n_8848)
);

AND2x2_ASAP7_75t_L g8849 ( 
.A(n_8241),
.B(n_2545),
.Y(n_8849)
);

NAND2xp5_ASAP7_75t_SL g8850 ( 
.A(n_8340),
.B(n_8342),
.Y(n_8850)
);

AOI21xp5_ASAP7_75t_L g8851 ( 
.A1(n_8234),
.A2(n_2547),
.B(n_2546),
.Y(n_8851)
);

OAI22xp5_ASAP7_75t_L g8852 ( 
.A1(n_8360),
.A2(n_2548),
.B1(n_2549),
.B2(n_2547),
.Y(n_8852)
);

INVx2_ASAP7_75t_L g8853 ( 
.A(n_8105),
.Y(n_8853)
);

AOI22xp33_ASAP7_75t_SL g8854 ( 
.A1(n_8286),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_8854)
);

HB1xp67_ASAP7_75t_L g8855 ( 
.A(n_8200),
.Y(n_8855)
);

INVx2_ASAP7_75t_L g8856 ( 
.A(n_8111),
.Y(n_8856)
);

INVx2_ASAP7_75t_L g8857 ( 
.A(n_8136),
.Y(n_8857)
);

INVx1_ASAP7_75t_L g8858 ( 
.A(n_8160),
.Y(n_8858)
);

INVx2_ASAP7_75t_SL g8859 ( 
.A(n_7884),
.Y(n_8859)
);

NOR2xp67_ASAP7_75t_L g8860 ( 
.A(n_7747),
.B(n_98),
.Y(n_8860)
);

NAND2xp5_ASAP7_75t_L g8861 ( 
.A(n_7958),
.B(n_98),
.Y(n_8861)
);

NAND2xp5_ASAP7_75t_SL g8862 ( 
.A(n_8343),
.B(n_2548),
.Y(n_8862)
);

INVx2_ASAP7_75t_L g8863 ( 
.A(n_8139),
.Y(n_8863)
);

NAND2xp5_ASAP7_75t_L g8864 ( 
.A(n_7960),
.B(n_98),
.Y(n_8864)
);

INVx2_ASAP7_75t_L g8865 ( 
.A(n_8148),
.Y(n_8865)
);

AOI22xp5_ASAP7_75t_L g8866 ( 
.A1(n_8141),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_8866)
);

AND2x4_ASAP7_75t_L g8867 ( 
.A(n_8040),
.B(n_99),
.Y(n_8867)
);

INVx2_ASAP7_75t_L g8868 ( 
.A(n_8161),
.Y(n_8868)
);

AOI22xp33_ASAP7_75t_L g8869 ( 
.A1(n_8332),
.A2(n_8141),
.B1(n_7989),
.B2(n_8112),
.Y(n_8869)
);

INVx2_ASAP7_75t_L g8870 ( 
.A(n_8166),
.Y(n_8870)
);

AND2x2_ASAP7_75t_L g8871 ( 
.A(n_8247),
.B(n_2550),
.Y(n_8871)
);

AOI22xp5_ASAP7_75t_L g8872 ( 
.A1(n_8013),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_8872)
);

NAND2xp5_ASAP7_75t_L g8873 ( 
.A(n_7961),
.B(n_100),
.Y(n_8873)
);

NAND2xp5_ASAP7_75t_L g8874 ( 
.A(n_8221),
.B(n_101),
.Y(n_8874)
);

NAND2xp5_ASAP7_75t_L g8875 ( 
.A(n_8225),
.B(n_102),
.Y(n_8875)
);

NAND2xp5_ASAP7_75t_L g8876 ( 
.A(n_8162),
.B(n_102),
.Y(n_8876)
);

AND3x1_ASAP7_75t_L g8877 ( 
.A(n_8276),
.B(n_102),
.C(n_103),
.Y(n_8877)
);

NAND2xp5_ASAP7_75t_L g8878 ( 
.A(n_8169),
.B(n_103),
.Y(n_8878)
);

NOR2xp33_ASAP7_75t_L g8879 ( 
.A(n_7746),
.B(n_2550),
.Y(n_8879)
);

NAND2xp5_ASAP7_75t_L g8880 ( 
.A(n_8172),
.B(n_103),
.Y(n_8880)
);

BUFx6f_ASAP7_75t_L g8881 ( 
.A(n_7959),
.Y(n_8881)
);

INVxp67_ASAP7_75t_L g8882 ( 
.A(n_8345),
.Y(n_8882)
);

NOR2x1p5_ASAP7_75t_L g8883 ( 
.A(n_8362),
.B(n_2551),
.Y(n_8883)
);

NOR2xp33_ASAP7_75t_L g8884 ( 
.A(n_8363),
.B(n_2552),
.Y(n_8884)
);

INVx5_ASAP7_75t_L g8885 ( 
.A(n_8063),
.Y(n_8885)
);

AOI22xp33_ASAP7_75t_L g8886 ( 
.A1(n_8396),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_8886)
);

INVx2_ASAP7_75t_L g8887 ( 
.A(n_8167),
.Y(n_8887)
);

AND2x6_ASAP7_75t_SL g8888 ( 
.A(n_7912),
.B(n_104),
.Y(n_8888)
);

O2A1O1Ixp5_ASAP7_75t_L g8889 ( 
.A1(n_7878),
.A2(n_107),
.B(n_105),
.C(n_106),
.Y(n_8889)
);

INVx1_ASAP7_75t_L g8890 ( 
.A(n_8174),
.Y(n_8890)
);

INVx2_ASAP7_75t_L g8891 ( 
.A(n_8168),
.Y(n_8891)
);

NAND2xp5_ASAP7_75t_SL g8892 ( 
.A(n_8009),
.B(n_2552),
.Y(n_8892)
);

NAND2xp5_ASAP7_75t_L g8893 ( 
.A(n_8178),
.B(n_106),
.Y(n_8893)
);

INVxp67_ASAP7_75t_L g8894 ( 
.A(n_8346),
.Y(n_8894)
);

NOR2xp33_ASAP7_75t_L g8895 ( 
.A(n_8366),
.B(n_2553),
.Y(n_8895)
);

INVx2_ASAP7_75t_SL g8896 ( 
.A(n_7786),
.Y(n_8896)
);

INVxp67_ASAP7_75t_L g8897 ( 
.A(n_8350),
.Y(n_8897)
);

NAND2xp5_ASAP7_75t_L g8898 ( 
.A(n_8183),
.B(n_107),
.Y(n_8898)
);

AND2x2_ASAP7_75t_SL g8899 ( 
.A(n_8386),
.B(n_107),
.Y(n_8899)
);

HB1xp67_ASAP7_75t_L g8900 ( 
.A(n_8352),
.Y(n_8900)
);

NOR2xp33_ASAP7_75t_L g8901 ( 
.A(n_8229),
.B(n_2553),
.Y(n_8901)
);

INVx2_ASAP7_75t_L g8902 ( 
.A(n_8202),
.Y(n_8902)
);

INVx4_ASAP7_75t_L g8903 ( 
.A(n_7882),
.Y(n_8903)
);

INVx1_ASAP7_75t_L g8904 ( 
.A(n_7968),
.Y(n_8904)
);

NAND2xp5_ASAP7_75t_L g8905 ( 
.A(n_8210),
.B(n_108),
.Y(n_8905)
);

INVx1_ASAP7_75t_L g8906 ( 
.A(n_8153),
.Y(n_8906)
);

AOI22xp33_ASAP7_75t_L g8907 ( 
.A1(n_7972),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_8907)
);

INVx2_ASAP7_75t_L g8908 ( 
.A(n_8208),
.Y(n_8908)
);

NOR2xp33_ASAP7_75t_SL g8909 ( 
.A(n_7863),
.B(n_109),
.Y(n_8909)
);

NOR2xp33_ASAP7_75t_L g8910 ( 
.A(n_7908),
.B(n_109),
.Y(n_8910)
);

AND2x4_ASAP7_75t_L g8911 ( 
.A(n_7821),
.B(n_110),
.Y(n_8911)
);

INVx2_ASAP7_75t_L g8912 ( 
.A(n_8209),
.Y(n_8912)
);

NAND2xp5_ASAP7_75t_SL g8913 ( 
.A(n_8214),
.B(n_111),
.Y(n_8913)
);

NAND2xp5_ASAP7_75t_L g8914 ( 
.A(n_8226),
.B(n_111),
.Y(n_8914)
);

NOR2xp33_ASAP7_75t_R g8915 ( 
.A(n_8002),
.B(n_111),
.Y(n_8915)
);

NAND2xp5_ASAP7_75t_L g8916 ( 
.A(n_8228),
.B(n_112),
.Y(n_8916)
);

NOR2xp67_ASAP7_75t_SL g8917 ( 
.A(n_8114),
.B(n_113),
.Y(n_8917)
);

INVx1_ASAP7_75t_L g8918 ( 
.A(n_8181),
.Y(n_8918)
);

NAND2xp5_ASAP7_75t_SL g8919 ( 
.A(n_8216),
.B(n_8024),
.Y(n_8919)
);

AND2x4_ASAP7_75t_L g8920 ( 
.A(n_8119),
.B(n_113),
.Y(n_8920)
);

HB1xp67_ASAP7_75t_L g8921 ( 
.A(n_8354),
.Y(n_8921)
);

NAND2xp5_ASAP7_75t_SL g8922 ( 
.A(n_7762),
.B(n_114),
.Y(n_8922)
);

NAND2xp5_ASAP7_75t_L g8923 ( 
.A(n_8230),
.B(n_115),
.Y(n_8923)
);

NAND2xp5_ASAP7_75t_L g8924 ( 
.A(n_8231),
.B(n_115),
.Y(n_8924)
);

NAND2xp5_ASAP7_75t_L g8925 ( 
.A(n_8232),
.B(n_115),
.Y(n_8925)
);

INVxp67_ASAP7_75t_L g8926 ( 
.A(n_8355),
.Y(n_8926)
);

AOI22xp33_ASAP7_75t_L g8927 ( 
.A1(n_8235),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_8927)
);

INVx2_ASAP7_75t_SL g8928 ( 
.A(n_8026),
.Y(n_8928)
);

INVx1_ASAP7_75t_L g8929 ( 
.A(n_8182),
.Y(n_8929)
);

INVx1_ASAP7_75t_L g8930 ( 
.A(n_8217),
.Y(n_8930)
);

NAND2xp5_ASAP7_75t_L g8931 ( 
.A(n_8236),
.B(n_116),
.Y(n_8931)
);

NAND2xp5_ASAP7_75t_L g8932 ( 
.A(n_8238),
.B(n_117),
.Y(n_8932)
);

INVx1_ASAP7_75t_L g8933 ( 
.A(n_8233),
.Y(n_8933)
);

INVx2_ASAP7_75t_L g8934 ( 
.A(n_8189),
.Y(n_8934)
);

NAND2xp5_ASAP7_75t_SL g8935 ( 
.A(n_8359),
.B(n_117),
.Y(n_8935)
);

INVxp67_ASAP7_75t_SL g8936 ( 
.A(n_8243),
.Y(n_8936)
);

NAND2xp5_ASAP7_75t_SL g8937 ( 
.A(n_8374),
.B(n_8356),
.Y(n_8937)
);

NAND2xp5_ASAP7_75t_SL g8938 ( 
.A(n_8367),
.B(n_118),
.Y(n_8938)
);

NAND2xp5_ASAP7_75t_SL g8939 ( 
.A(n_8369),
.B(n_118),
.Y(n_8939)
);

NAND2xp5_ASAP7_75t_SL g8940 ( 
.A(n_8376),
.B(n_119),
.Y(n_8940)
);

NAND2xp5_ASAP7_75t_L g8941 ( 
.A(n_8007),
.B(n_119),
.Y(n_8941)
);

INVx2_ASAP7_75t_L g8942 ( 
.A(n_8028),
.Y(n_8942)
);

INVx1_ASAP7_75t_L g8943 ( 
.A(n_8029),
.Y(n_8943)
);

INVx2_ASAP7_75t_L g8944 ( 
.A(n_8031),
.Y(n_8944)
);

INVx1_ASAP7_75t_L g8945 ( 
.A(n_8035),
.Y(n_8945)
);

HB1xp67_ASAP7_75t_L g8946 ( 
.A(n_8142),
.Y(n_8946)
);

NAND2xp5_ASAP7_75t_L g8947 ( 
.A(n_8389),
.B(n_120),
.Y(n_8947)
);

INVx1_ASAP7_75t_L g8948 ( 
.A(n_8043),
.Y(n_8948)
);

NAND2xp5_ASAP7_75t_L g8949 ( 
.A(n_8390),
.B(n_120),
.Y(n_8949)
);

BUFx8_ASAP7_75t_L g8950 ( 
.A(n_8328),
.Y(n_8950)
);

AND2x2_ASAP7_75t_L g8951 ( 
.A(n_8176),
.B(n_8135),
.Y(n_8951)
);

NAND2xp5_ASAP7_75t_SL g8952 ( 
.A(n_8377),
.B(n_121),
.Y(n_8952)
);

INVx2_ASAP7_75t_L g8953 ( 
.A(n_8044),
.Y(n_8953)
);

NAND2xp5_ASAP7_75t_L g8954 ( 
.A(n_8045),
.B(n_121),
.Y(n_8954)
);

INVx5_ASAP7_75t_L g8955 ( 
.A(n_8381),
.Y(n_8955)
);

NOR2xp33_ASAP7_75t_L g8956 ( 
.A(n_8344),
.B(n_121),
.Y(n_8956)
);

NOR2xp33_ASAP7_75t_L g8957 ( 
.A(n_7916),
.B(n_122),
.Y(n_8957)
);

NAND2xp5_ASAP7_75t_L g8958 ( 
.A(n_8047),
.B(n_122),
.Y(n_8958)
);

OR2x6_ASAP7_75t_L g8959 ( 
.A(n_8251),
.B(n_122),
.Y(n_8959)
);

NAND2xp5_ASAP7_75t_SL g8960 ( 
.A(n_8058),
.B(n_123),
.Y(n_8960)
);

NAND2xp5_ASAP7_75t_SL g8961 ( 
.A(n_8133),
.B(n_123),
.Y(n_8961)
);

INVx2_ASAP7_75t_L g8962 ( 
.A(n_8055),
.Y(n_8962)
);

HB1xp67_ASAP7_75t_L g8963 ( 
.A(n_8173),
.Y(n_8963)
);

NAND2xp5_ASAP7_75t_L g8964 ( 
.A(n_8060),
.B(n_123),
.Y(n_8964)
);

INVx1_ASAP7_75t_L g8965 ( 
.A(n_8067),
.Y(n_8965)
);

NAND2xp5_ASAP7_75t_L g8966 ( 
.A(n_8071),
.B(n_124),
.Y(n_8966)
);

INVx2_ASAP7_75t_L g8967 ( 
.A(n_8074),
.Y(n_8967)
);

NOR2xp33_ASAP7_75t_L g8968 ( 
.A(n_8163),
.B(n_124),
.Y(n_8968)
);

NAND2xp5_ASAP7_75t_L g8969 ( 
.A(n_8077),
.B(n_124),
.Y(n_8969)
);

OR2x2_ASAP7_75t_L g8970 ( 
.A(n_8299),
.B(n_125),
.Y(n_8970)
);

NAND2xp5_ASAP7_75t_SL g8971 ( 
.A(n_8020),
.B(n_125),
.Y(n_8971)
);

NOR2xp33_ASAP7_75t_L g8972 ( 
.A(n_8193),
.B(n_125),
.Y(n_8972)
);

BUFx6f_ASAP7_75t_L g8973 ( 
.A(n_7939),
.Y(n_8973)
);

NAND3xp33_ASAP7_75t_L g8974 ( 
.A(n_8265),
.B(n_126),
.C(n_127),
.Y(n_8974)
);

NAND2xp5_ASAP7_75t_L g8975 ( 
.A(n_8078),
.B(n_126),
.Y(n_8975)
);

NAND2xp5_ASAP7_75t_L g8976 ( 
.A(n_8079),
.B(n_126),
.Y(n_8976)
);

NOR2xp33_ASAP7_75t_L g8977 ( 
.A(n_8259),
.B(n_127),
.Y(n_8977)
);

NAND2xp5_ASAP7_75t_L g8978 ( 
.A(n_8081),
.B(n_127),
.Y(n_8978)
);

INVx2_ASAP7_75t_L g8979 ( 
.A(n_8083),
.Y(n_8979)
);

HB1xp67_ASAP7_75t_L g8980 ( 
.A(n_8049),
.Y(n_8980)
);

O2A1O1Ixp5_ASAP7_75t_L g8981 ( 
.A1(n_7860),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_8981)
);

INVx1_ASAP7_75t_L g8982 ( 
.A(n_8085),
.Y(n_8982)
);

NAND2xp5_ASAP7_75t_L g8983 ( 
.A(n_8086),
.B(n_128),
.Y(n_8983)
);

OAI22xp5_ASAP7_75t_L g8984 ( 
.A1(n_8405),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_8984)
);

NAND2xp5_ASAP7_75t_SL g8985 ( 
.A(n_8258),
.B(n_129),
.Y(n_8985)
);

INVx2_ASAP7_75t_L g8986 ( 
.A(n_8087),
.Y(n_8986)
);

NOR2xp33_ASAP7_75t_L g8987 ( 
.A(n_8070),
.B(n_130),
.Y(n_8987)
);

AOI22xp33_ASAP7_75t_L g8988 ( 
.A1(n_8250),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_8988)
);

OR2x2_ASAP7_75t_L g8989 ( 
.A(n_8088),
.B(n_132),
.Y(n_8989)
);

NOR2xp33_ASAP7_75t_L g8990 ( 
.A(n_8284),
.B(n_133),
.Y(n_8990)
);

NAND2xp5_ASAP7_75t_SL g8991 ( 
.A(n_7951),
.B(n_133),
.Y(n_8991)
);

AOI22xp5_ASAP7_75t_L g8992 ( 
.A1(n_8097),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_8992)
);

INVx2_ASAP7_75t_L g8993 ( 
.A(n_8092),
.Y(n_8993)
);

NAND2xp5_ASAP7_75t_L g8994 ( 
.A(n_8094),
.B(n_134),
.Y(n_8994)
);

AOI22xp33_ASAP7_75t_L g8995 ( 
.A1(n_8268),
.A2(n_137),
.B1(n_134),
.B2(n_136),
.Y(n_8995)
);

AND2x6_ASAP7_75t_SL g8996 ( 
.A(n_7760),
.B(n_137),
.Y(n_8996)
);

NAND2xp5_ASAP7_75t_L g8997 ( 
.A(n_8095),
.B(n_138),
.Y(n_8997)
);

INVx1_ASAP7_75t_L g8998 ( 
.A(n_8096),
.Y(n_8998)
);

INVx2_ASAP7_75t_L g8999 ( 
.A(n_8099),
.Y(n_8999)
);

HB1xp67_ASAP7_75t_L g9000 ( 
.A(n_8256),
.Y(n_9000)
);

NOR2xp33_ASAP7_75t_L g9001 ( 
.A(n_8392),
.B(n_7828),
.Y(n_9001)
);

NOR2xp33_ASAP7_75t_L g9002 ( 
.A(n_8375),
.B(n_138),
.Y(n_9002)
);

INVx2_ASAP7_75t_SL g9003 ( 
.A(n_8296),
.Y(n_9003)
);

AOI22xp33_ASAP7_75t_L g9004 ( 
.A1(n_8298),
.A2(n_8260),
.B1(n_8262),
.B2(n_8257),
.Y(n_9004)
);

NAND2xp5_ASAP7_75t_SL g9005 ( 
.A(n_8364),
.B(n_138),
.Y(n_9005)
);

INVxp67_ASAP7_75t_L g9006 ( 
.A(n_8263),
.Y(n_9006)
);

AND2x2_ASAP7_75t_L g9007 ( 
.A(n_8033),
.B(n_139),
.Y(n_9007)
);

CKINVDCx5p33_ASAP7_75t_R g9008 ( 
.A(n_7936),
.Y(n_9008)
);

INVx2_ASAP7_75t_L g9009 ( 
.A(n_8101),
.Y(n_9009)
);

INVx2_ASAP7_75t_SL g9010 ( 
.A(n_8264),
.Y(n_9010)
);

NAND2xp5_ASAP7_75t_L g9011 ( 
.A(n_8103),
.B(n_139),
.Y(n_9011)
);

INVx1_ASAP7_75t_L g9012 ( 
.A(n_8104),
.Y(n_9012)
);

NAND2xp5_ASAP7_75t_L g9013 ( 
.A(n_8106),
.B(n_139),
.Y(n_9013)
);

NAND2xp5_ASAP7_75t_SL g9014 ( 
.A(n_8372),
.B(n_140),
.Y(n_9014)
);

INVx4_ASAP7_75t_L g9015 ( 
.A(n_8349),
.Y(n_9015)
);

NOR2xp33_ASAP7_75t_L g9016 ( 
.A(n_8419),
.B(n_8266),
.Y(n_9016)
);

INVx1_ASAP7_75t_L g9017 ( 
.A(n_8690),
.Y(n_9017)
);

AOI22xp5_ASAP7_75t_L g9018 ( 
.A1(n_8540),
.A2(n_8272),
.B1(n_8273),
.B2(n_8270),
.Y(n_9018)
);

INVx1_ASAP7_75t_L g9019 ( 
.A(n_8726),
.Y(n_9019)
);

AND2x6_ASAP7_75t_SL g9020 ( 
.A(n_9001),
.B(n_8278),
.Y(n_9020)
);

BUFx3_ASAP7_75t_L g9021 ( 
.A(n_8596),
.Y(n_9021)
);

AND2x4_ASAP7_75t_L g9022 ( 
.A(n_8432),
.B(n_8280),
.Y(n_9022)
);

AND2x4_ASAP7_75t_L g9023 ( 
.A(n_8429),
.B(n_8281),
.Y(n_9023)
);

NAND2xp5_ASAP7_75t_L g9024 ( 
.A(n_8588),
.B(n_8108),
.Y(n_9024)
);

NAND2xp5_ASAP7_75t_L g9025 ( 
.A(n_8594),
.B(n_8109),
.Y(n_9025)
);

NAND2xp5_ASAP7_75t_L g9026 ( 
.A(n_8518),
.B(n_8110),
.Y(n_9026)
);

OR2x2_ASAP7_75t_L g9027 ( 
.A(n_8519),
.B(n_8283),
.Y(n_9027)
);

NAND2xp5_ASAP7_75t_SL g9028 ( 
.A(n_8501),
.B(n_8244),
.Y(n_9028)
);

O2A1O1Ixp5_ASAP7_75t_L g9029 ( 
.A1(n_8433),
.A2(n_7743),
.B(n_8249),
.C(n_8245),
.Y(n_9029)
);

AOI21xp5_ASAP7_75t_L g9030 ( 
.A1(n_8621),
.A2(n_8254),
.B(n_8305),
.Y(n_9030)
);

INVx1_ASAP7_75t_L g9031 ( 
.A(n_8730),
.Y(n_9031)
);

NOR2xp33_ASAP7_75t_L g9032 ( 
.A(n_8459),
.B(n_8288),
.Y(n_9032)
);

CKINVDCx5p33_ASAP7_75t_R g9033 ( 
.A(n_8431),
.Y(n_9033)
);

NAND2xp5_ASAP7_75t_L g9034 ( 
.A(n_8640),
.B(n_8113),
.Y(n_9034)
);

NAND2xp5_ASAP7_75t_L g9035 ( 
.A(n_8537),
.B(n_8116),
.Y(n_9035)
);

AND2x2_ASAP7_75t_L g9036 ( 
.A(n_8951),
.B(n_8289),
.Y(n_9036)
);

INVx1_ASAP7_75t_L g9037 ( 
.A(n_8748),
.Y(n_9037)
);

NAND2xp5_ASAP7_75t_SL g9038 ( 
.A(n_8422),
.B(n_8291),
.Y(n_9038)
);

AOI22xp5_ASAP7_75t_L g9039 ( 
.A1(n_8657),
.A2(n_8297),
.B1(n_8118),
.B2(n_8120),
.Y(n_9039)
);

AOI22xp5_ASAP7_75t_L g9040 ( 
.A1(n_8676),
.A2(n_8121),
.B1(n_8123),
.B2(n_8117),
.Y(n_9040)
);

NAND2xp5_ASAP7_75t_L g9041 ( 
.A(n_8525),
.B(n_8125),
.Y(n_9041)
);

NOR3xp33_ASAP7_75t_SL g9042 ( 
.A(n_8412),
.B(n_8763),
.C(n_8826),
.Y(n_9042)
);

NOR2xp33_ASAP7_75t_L g9043 ( 
.A(n_8421),
.B(n_8126),
.Y(n_9043)
);

AND2x4_ASAP7_75t_L g9044 ( 
.A(n_8814),
.B(n_8131),
.Y(n_9044)
);

NAND2xp5_ASAP7_75t_L g9045 ( 
.A(n_8489),
.B(n_8138),
.Y(n_9045)
);

NOR2xp33_ASAP7_75t_L g9046 ( 
.A(n_8427),
.B(n_8140),
.Y(n_9046)
);

NAND2xp5_ASAP7_75t_L g9047 ( 
.A(n_8499),
.B(n_8143),
.Y(n_9047)
);

NAND2xp5_ASAP7_75t_SL g9048 ( 
.A(n_8467),
.B(n_8749),
.Y(n_9048)
);

INVx2_ASAP7_75t_L g9049 ( 
.A(n_8528),
.Y(n_9049)
);

NAND2xp5_ASAP7_75t_L g9050 ( 
.A(n_8506),
.B(n_8144),
.Y(n_9050)
);

BUFx12f_ASAP7_75t_L g9051 ( 
.A(n_8598),
.Y(n_9051)
);

AND2x2_ASAP7_75t_L g9052 ( 
.A(n_8418),
.B(n_8149),
.Y(n_9052)
);

INVx2_ASAP7_75t_L g9053 ( 
.A(n_8530),
.Y(n_9053)
);

INVx2_ASAP7_75t_L g9054 ( 
.A(n_8532),
.Y(n_9054)
);

INVx2_ASAP7_75t_SL g9055 ( 
.A(n_8654),
.Y(n_9055)
);

AND2x4_ASAP7_75t_L g9056 ( 
.A(n_8622),
.B(n_8150),
.Y(n_9056)
);

CKINVDCx5p33_ASAP7_75t_R g9057 ( 
.A(n_8700),
.Y(n_9057)
);

AOI22xp5_ASAP7_75t_L g9058 ( 
.A1(n_8681),
.A2(n_8152),
.B1(n_8179),
.B2(n_8151),
.Y(n_9058)
);

INVx2_ASAP7_75t_L g9059 ( 
.A(n_8557),
.Y(n_9059)
);

OR2x4_ASAP7_75t_L g9060 ( 
.A(n_8477),
.B(n_8184),
.Y(n_9060)
);

NAND2xp5_ASAP7_75t_L g9061 ( 
.A(n_8526),
.B(n_8187),
.Y(n_9061)
);

INVx1_ASAP7_75t_L g9062 ( 
.A(n_8788),
.Y(n_9062)
);

NAND2xp5_ASAP7_75t_L g9063 ( 
.A(n_8517),
.B(n_8188),
.Y(n_9063)
);

INVx2_ASAP7_75t_L g9064 ( 
.A(n_8559),
.Y(n_9064)
);

OAI21xp33_ASAP7_75t_SL g9065 ( 
.A1(n_8701),
.A2(n_8192),
.B(n_8191),
.Y(n_9065)
);

BUFx6f_ASAP7_75t_L g9066 ( 
.A(n_8411),
.Y(n_9066)
);

BUFx8_ASAP7_75t_L g9067 ( 
.A(n_8693),
.Y(n_9067)
);

INVx1_ASAP7_75t_L g9068 ( 
.A(n_8813),
.Y(n_9068)
);

NAND3xp33_ASAP7_75t_SL g9069 ( 
.A(n_8437),
.B(n_8196),
.C(n_8194),
.Y(n_9069)
);

INVxp67_ASAP7_75t_L g9070 ( 
.A(n_8509),
.Y(n_9070)
);

INVx2_ASAP7_75t_L g9071 ( 
.A(n_8569),
.Y(n_9071)
);

INVx1_ASAP7_75t_SL g9072 ( 
.A(n_8575),
.Y(n_9072)
);

CKINVDCx5p33_ASAP7_75t_R g9073 ( 
.A(n_8700),
.Y(n_9073)
);

INVx1_ASAP7_75t_L g9074 ( 
.A(n_8834),
.Y(n_9074)
);

INVx2_ASAP7_75t_SL g9075 ( 
.A(n_8806),
.Y(n_9075)
);

NAND2xp5_ASAP7_75t_L g9076 ( 
.A(n_8476),
.B(n_8197),
.Y(n_9076)
);

INVx1_ASAP7_75t_L g9077 ( 
.A(n_8848),
.Y(n_9077)
);

NOR3xp33_ASAP7_75t_SL g9078 ( 
.A(n_8727),
.B(n_8199),
.C(n_8198),
.Y(n_9078)
);

CKINVDCx5p33_ASAP7_75t_R g9079 ( 
.A(n_8411),
.Y(n_9079)
);

NOR2xp33_ASAP7_75t_L g9080 ( 
.A(n_8430),
.B(n_8203),
.Y(n_9080)
);

AOI22xp33_ASAP7_75t_L g9081 ( 
.A1(n_8424),
.A2(n_8204),
.B1(n_8353),
.B2(n_8334),
.Y(n_9081)
);

NAND2xp5_ASAP7_75t_L g9082 ( 
.A(n_8514),
.B(n_8358),
.Y(n_9082)
);

INVx2_ASAP7_75t_L g9083 ( 
.A(n_8577),
.Y(n_9083)
);

INVx1_ASAP7_75t_L g9084 ( 
.A(n_8600),
.Y(n_9084)
);

INVx2_ASAP7_75t_L g9085 ( 
.A(n_8579),
.Y(n_9085)
);

NAND2xp5_ASAP7_75t_L g9086 ( 
.A(n_8446),
.B(n_140),
.Y(n_9086)
);

INVx1_ASAP7_75t_L g9087 ( 
.A(n_8414),
.Y(n_9087)
);

AND2x6_ASAP7_75t_SL g9088 ( 
.A(n_8551),
.B(n_140),
.Y(n_9088)
);

NAND2xp5_ASAP7_75t_L g9089 ( 
.A(n_8707),
.B(n_141),
.Y(n_9089)
);

NAND2xp5_ASAP7_75t_SL g9090 ( 
.A(n_8749),
.B(n_141),
.Y(n_9090)
);

NAND2xp5_ASAP7_75t_L g9091 ( 
.A(n_8512),
.B(n_141),
.Y(n_9091)
);

NAND2xp5_ASAP7_75t_SL g9092 ( 
.A(n_8749),
.B(n_142),
.Y(n_9092)
);

BUFx2_ASAP7_75t_L g9093 ( 
.A(n_8946),
.Y(n_9093)
);

INVx1_ASAP7_75t_L g9094 ( 
.A(n_8439),
.Y(n_9094)
);

BUFx2_ASAP7_75t_L g9095 ( 
.A(n_8521),
.Y(n_9095)
);

NAND2xp5_ASAP7_75t_L g9096 ( 
.A(n_8538),
.B(n_8547),
.Y(n_9096)
);

NAND2xp5_ASAP7_75t_L g9097 ( 
.A(n_8583),
.B(n_142),
.Y(n_9097)
);

INVx1_ASAP7_75t_L g9098 ( 
.A(n_8441),
.Y(n_9098)
);

AND2x6_ASAP7_75t_SL g9099 ( 
.A(n_8968),
.B(n_142),
.Y(n_9099)
);

NAND2xp5_ASAP7_75t_L g9100 ( 
.A(n_8591),
.B(n_143),
.Y(n_9100)
);

BUFx8_ASAP7_75t_L g9101 ( 
.A(n_8973),
.Y(n_9101)
);

OAI22xp5_ASAP7_75t_L g9102 ( 
.A1(n_8502),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_9102)
);

NOR2xp33_ASAP7_75t_L g9103 ( 
.A(n_8415),
.B(n_144),
.Y(n_9103)
);

NAND2xp5_ASAP7_75t_SL g9104 ( 
.A(n_8749),
.B(n_144),
.Y(n_9104)
);

NAND3xp33_ASAP7_75t_L g9105 ( 
.A(n_8638),
.B(n_145),
.C(n_146),
.Y(n_9105)
);

INVx2_ASAP7_75t_SL g9106 ( 
.A(n_8806),
.Y(n_9106)
);

NAND3xp33_ASAP7_75t_L g9107 ( 
.A(n_8484),
.B(n_8616),
.C(n_8491),
.Y(n_9107)
);

INVx1_ASAP7_75t_SL g9108 ( 
.A(n_8447),
.Y(n_9108)
);

NAND2xp5_ASAP7_75t_SL g9109 ( 
.A(n_8508),
.B(n_8451),
.Y(n_9109)
);

INVx2_ASAP7_75t_L g9110 ( 
.A(n_8584),
.Y(n_9110)
);

INVx2_ASAP7_75t_SL g9111 ( 
.A(n_8464),
.Y(n_9111)
);

INVxp67_ASAP7_75t_L g9112 ( 
.A(n_8487),
.Y(n_9112)
);

NAND2xp5_ASAP7_75t_L g9113 ( 
.A(n_8606),
.B(n_146),
.Y(n_9113)
);

BUFx6f_ASAP7_75t_SL g9114 ( 
.A(n_8903),
.Y(n_9114)
);

INVx2_ASAP7_75t_L g9115 ( 
.A(n_8592),
.Y(n_9115)
);

AOI22xp33_ASAP7_75t_L g9116 ( 
.A1(n_8426),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_9116)
);

INVx1_ASAP7_75t_L g9117 ( 
.A(n_8458),
.Y(n_9117)
);

INVx1_ASAP7_75t_L g9118 ( 
.A(n_8461),
.Y(n_9118)
);

INVx2_ASAP7_75t_L g9119 ( 
.A(n_8599),
.Y(n_9119)
);

BUFx3_ASAP7_75t_L g9120 ( 
.A(n_8950),
.Y(n_9120)
);

INVx2_ASAP7_75t_SL g9121 ( 
.A(n_8759),
.Y(n_9121)
);

AOI22xp33_ASAP7_75t_SL g9122 ( 
.A1(n_8767),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_9122)
);

NAND2xp5_ASAP7_75t_SL g9123 ( 
.A(n_8444),
.B(n_147),
.Y(n_9123)
);

INVx2_ASAP7_75t_L g9124 ( 
.A(n_8416),
.Y(n_9124)
);

NAND2xp5_ASAP7_75t_L g9125 ( 
.A(n_8513),
.B(n_148),
.Y(n_9125)
);

INVx1_ASAP7_75t_L g9126 ( 
.A(n_8462),
.Y(n_9126)
);

NAND2xp5_ASAP7_75t_L g9127 ( 
.A(n_8513),
.B(n_149),
.Y(n_9127)
);

NAND2xp5_ASAP7_75t_L g9128 ( 
.A(n_8513),
.B(n_150),
.Y(n_9128)
);

INVx3_ASAP7_75t_L g9129 ( 
.A(n_8759),
.Y(n_9129)
);

AOI22xp5_ASAP7_75t_L g9130 ( 
.A1(n_8685),
.A2(n_8667),
.B1(n_8648),
.B2(n_8553),
.Y(n_9130)
);

AND2x4_ASAP7_75t_L g9131 ( 
.A(n_8955),
.B(n_8542),
.Y(n_9131)
);

INVx3_ASAP7_75t_L g9132 ( 
.A(n_8434),
.Y(n_9132)
);

NAND2xp5_ASAP7_75t_L g9133 ( 
.A(n_8554),
.B(n_150),
.Y(n_9133)
);

NOR2xp33_ASAP7_75t_L g9134 ( 
.A(n_8440),
.B(n_150),
.Y(n_9134)
);

INVx2_ASAP7_75t_L g9135 ( 
.A(n_8417),
.Y(n_9135)
);

NAND2xp5_ASAP7_75t_SL g9136 ( 
.A(n_8607),
.B(n_8709),
.Y(n_9136)
);

INVx2_ASAP7_75t_SL g9137 ( 
.A(n_8885),
.Y(n_9137)
);

INVx3_ASAP7_75t_L g9138 ( 
.A(n_8881),
.Y(n_9138)
);

INVx1_ASAP7_75t_L g9139 ( 
.A(n_8466),
.Y(n_9139)
);

NAND2xp5_ASAP7_75t_L g9140 ( 
.A(n_8535),
.B(n_151),
.Y(n_9140)
);

OAI22xp5_ASAP7_75t_SL g9141 ( 
.A1(n_8661),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_9141)
);

AOI22xp33_ASAP7_75t_L g9142 ( 
.A1(n_8818),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_9142)
);

INVx5_ASAP7_75t_L g9143 ( 
.A(n_8604),
.Y(n_9143)
);

AOI22xp33_ASAP7_75t_L g9144 ( 
.A1(n_8869),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_9144)
);

NAND2xp5_ASAP7_75t_SL g9145 ( 
.A(n_8615),
.B(n_154),
.Y(n_9145)
);

INVx2_ASAP7_75t_L g9146 ( 
.A(n_8423),
.Y(n_9146)
);

INVx1_ASAP7_75t_L g9147 ( 
.A(n_8471),
.Y(n_9147)
);

INVx2_ASAP7_75t_L g9148 ( 
.A(n_8425),
.Y(n_9148)
);

HB1xp67_ASAP7_75t_L g9149 ( 
.A(n_8900),
.Y(n_9149)
);

INVx1_ASAP7_75t_L g9150 ( 
.A(n_8480),
.Y(n_9150)
);

NAND2xp5_ASAP7_75t_L g9151 ( 
.A(n_8527),
.B(n_155),
.Y(n_9151)
);

CKINVDCx20_ASAP7_75t_R g9152 ( 
.A(n_8651),
.Y(n_9152)
);

A2O1A1Ixp33_ASAP7_75t_L g9153 ( 
.A1(n_8545),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_9153)
);

AND2x6_ASAP7_75t_SL g9154 ( 
.A(n_8972),
.B(n_156),
.Y(n_9154)
);

INVx2_ASAP7_75t_L g9155 ( 
.A(n_8428),
.Y(n_9155)
);

INVxp67_ASAP7_75t_L g9156 ( 
.A(n_8445),
.Y(n_9156)
);

NAND2xp5_ASAP7_75t_L g9157 ( 
.A(n_8544),
.B(n_157),
.Y(n_9157)
);

NAND2xp5_ASAP7_75t_L g9158 ( 
.A(n_8980),
.B(n_158),
.Y(n_9158)
);

INVx3_ASAP7_75t_L g9159 ( 
.A(n_8881),
.Y(n_9159)
);

INVx4_ASAP7_75t_L g9160 ( 
.A(n_8955),
.Y(n_9160)
);

NAND2xp5_ASAP7_75t_SL g9161 ( 
.A(n_8624),
.B(n_158),
.Y(n_9161)
);

NAND2xp5_ASAP7_75t_SL g9162 ( 
.A(n_8628),
.B(n_158),
.Y(n_9162)
);

INVx1_ASAP7_75t_L g9163 ( 
.A(n_8485),
.Y(n_9163)
);

INVxp33_ASAP7_75t_SL g9164 ( 
.A(n_8548),
.Y(n_9164)
);

NOR2xp33_ASAP7_75t_L g9165 ( 
.A(n_8523),
.B(n_8495),
.Y(n_9165)
);

INVx1_ASAP7_75t_L g9166 ( 
.A(n_8486),
.Y(n_9166)
);

INVx1_ASAP7_75t_L g9167 ( 
.A(n_8493),
.Y(n_9167)
);

AOI22xp33_ASAP7_75t_L g9168 ( 
.A1(n_8703),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_9168)
);

AOI22xp5_ASAP7_75t_L g9169 ( 
.A1(n_8478),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_9169)
);

INVx2_ASAP7_75t_L g9170 ( 
.A(n_8435),
.Y(n_9170)
);

NAND2xp5_ASAP7_75t_L g9171 ( 
.A(n_8647),
.B(n_162),
.Y(n_9171)
);

NAND2xp5_ASAP7_75t_SL g9172 ( 
.A(n_8765),
.B(n_8799),
.Y(n_9172)
);

INVx2_ASAP7_75t_L g9173 ( 
.A(n_8438),
.Y(n_9173)
);

HB1xp67_ASAP7_75t_L g9174 ( 
.A(n_8921),
.Y(n_9174)
);

AOI21xp5_ASAP7_75t_L g9175 ( 
.A1(n_8539),
.A2(n_162),
.B(n_163),
.Y(n_9175)
);

INVx5_ASAP7_75t_L g9176 ( 
.A(n_8604),
.Y(n_9176)
);

NAND2xp5_ASAP7_75t_SL g9177 ( 
.A(n_8955),
.B(n_162),
.Y(n_9177)
);

OAI22xp5_ASAP7_75t_SL g9178 ( 
.A1(n_8620),
.A2(n_167),
.B1(n_164),
.B2(n_166),
.Y(n_9178)
);

NAND2xp5_ASAP7_75t_SL g9179 ( 
.A(n_8443),
.B(n_164),
.Y(n_9179)
);

NAND2xp5_ASAP7_75t_SL g9180 ( 
.A(n_8885),
.B(n_167),
.Y(n_9180)
);

INVx2_ASAP7_75t_L g9181 ( 
.A(n_8449),
.Y(n_9181)
);

NOR2xp33_ASAP7_75t_L g9182 ( 
.A(n_8420),
.B(n_168),
.Y(n_9182)
);

INVx2_ASAP7_75t_L g9183 ( 
.A(n_8452),
.Y(n_9183)
);

NOR3xp33_ASAP7_75t_SL g9184 ( 
.A(n_8675),
.B(n_168),
.C(n_169),
.Y(n_9184)
);

INVx1_ASAP7_75t_L g9185 ( 
.A(n_8498),
.Y(n_9185)
);

INVx1_ASAP7_75t_L g9186 ( 
.A(n_8511),
.Y(n_9186)
);

NAND2xp5_ASAP7_75t_L g9187 ( 
.A(n_8515),
.B(n_168),
.Y(n_9187)
);

INVx1_ASAP7_75t_L g9188 ( 
.A(n_8529),
.Y(n_9188)
);

INVx1_ASAP7_75t_L g9189 ( 
.A(n_8552),
.Y(n_9189)
);

HB1xp67_ASAP7_75t_L g9190 ( 
.A(n_8556),
.Y(n_9190)
);

INVx4_ASAP7_75t_L g9191 ( 
.A(n_8845),
.Y(n_9191)
);

INVx2_ASAP7_75t_L g9192 ( 
.A(n_8460),
.Y(n_9192)
);

NAND2xp5_ASAP7_75t_L g9193 ( 
.A(n_8566),
.B(n_169),
.Y(n_9193)
);

INVx1_ASAP7_75t_L g9194 ( 
.A(n_8567),
.Y(n_9194)
);

NAND2xp5_ASAP7_75t_L g9195 ( 
.A(n_8573),
.B(n_169),
.Y(n_9195)
);

NAND2xp5_ASAP7_75t_L g9196 ( 
.A(n_8574),
.B(n_170),
.Y(n_9196)
);

OR2x6_ASAP7_75t_L g9197 ( 
.A(n_8454),
.B(n_170),
.Y(n_9197)
);

AOI22xp33_ASAP7_75t_L g9198 ( 
.A1(n_8679),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_9198)
);

INVx2_ASAP7_75t_SL g9199 ( 
.A(n_8885),
.Y(n_9199)
);

AND2x4_ASAP7_75t_L g9200 ( 
.A(n_8453),
.B(n_8533),
.Y(n_9200)
);

INVx2_ASAP7_75t_L g9201 ( 
.A(n_8469),
.Y(n_9201)
);

NAND2xp5_ASAP7_75t_SL g9202 ( 
.A(n_8468),
.B(n_8549),
.Y(n_9202)
);

INVx1_ASAP7_75t_L g9203 ( 
.A(n_8581),
.Y(n_9203)
);

AOI22xp5_ASAP7_75t_L g9204 ( 
.A1(n_8842),
.A2(n_8909),
.B1(n_8660),
.B2(n_8666),
.Y(n_9204)
);

AOI22xp33_ASAP7_75t_SL g9205 ( 
.A1(n_8899),
.A2(n_174),
.B1(n_171),
.B2(n_172),
.Y(n_9205)
);

INVx2_ASAP7_75t_L g9206 ( 
.A(n_8470),
.Y(n_9206)
);

AND2x2_ASAP7_75t_L g9207 ( 
.A(n_8587),
.B(n_171),
.Y(n_9207)
);

NOR2xp33_ASAP7_75t_L g9208 ( 
.A(n_8560),
.B(n_172),
.Y(n_9208)
);

O2A1O1Ixp5_ASAP7_75t_L g9209 ( 
.A1(n_8614),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_9209)
);

AND2x4_ASAP7_75t_L g9210 ( 
.A(n_8413),
.B(n_174),
.Y(n_9210)
);

AND2x4_ASAP7_75t_L g9211 ( 
.A(n_8928),
.B(n_175),
.Y(n_9211)
);

INVx1_ASAP7_75t_L g9212 ( 
.A(n_8590),
.Y(n_9212)
);

AND2x6_ASAP7_75t_L g9213 ( 
.A(n_8866),
.B(n_175),
.Y(n_9213)
);

AOI22xp33_ASAP7_75t_L g9214 ( 
.A1(n_8854),
.A2(n_180),
.B1(n_177),
.B2(n_178),
.Y(n_9214)
);

AOI21xp5_ASAP7_75t_L g9215 ( 
.A1(n_8481),
.A2(n_177),
.B(n_178),
.Y(n_9215)
);

AND2x4_ASAP7_75t_L g9216 ( 
.A(n_8973),
.B(n_180),
.Y(n_9216)
);

NAND2xp5_ASAP7_75t_L g9217 ( 
.A(n_8597),
.B(n_180),
.Y(n_9217)
);

AND2x6_ASAP7_75t_L g9218 ( 
.A(n_8603),
.B(n_181),
.Y(n_9218)
);

AND2x4_ASAP7_75t_L g9219 ( 
.A(n_8639),
.B(n_181),
.Y(n_9219)
);

NAND2xp5_ASAP7_75t_L g9220 ( 
.A(n_8611),
.B(n_182),
.Y(n_9220)
);

NAND2xp5_ASAP7_75t_SL g9221 ( 
.A(n_8455),
.B(n_183),
.Y(n_9221)
);

NAND2xp5_ASAP7_75t_SL g9222 ( 
.A(n_8516),
.B(n_183),
.Y(n_9222)
);

NAND2xp5_ASAP7_75t_L g9223 ( 
.A(n_8612),
.B(n_183),
.Y(n_9223)
);

AOI22xp33_ASAP7_75t_L g9224 ( 
.A1(n_8561),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_9224)
);

OAI22xp33_ASAP7_75t_L g9225 ( 
.A1(n_8768),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_9225)
);

INVx1_ASAP7_75t_SL g9226 ( 
.A(n_8550),
.Y(n_9226)
);

NAND2xp5_ASAP7_75t_L g9227 ( 
.A(n_8617),
.B(n_8643),
.Y(n_9227)
);

INVx1_ASAP7_75t_L g9228 ( 
.A(n_8656),
.Y(n_9228)
);

NAND2xp5_ASAP7_75t_L g9229 ( 
.A(n_8665),
.B(n_8670),
.Y(n_9229)
);

AOI22xp33_ASAP7_75t_L g9230 ( 
.A1(n_8695),
.A2(n_187),
.B1(n_184),
.B2(n_185),
.Y(n_9230)
);

AND2x4_ASAP7_75t_L g9231 ( 
.A(n_8456),
.B(n_187),
.Y(n_9231)
);

INVx2_ASAP7_75t_L g9232 ( 
.A(n_8472),
.Y(n_9232)
);

INVx1_ASAP7_75t_L g9233 ( 
.A(n_8684),
.Y(n_9233)
);

NAND2xp5_ASAP7_75t_L g9234 ( 
.A(n_8706),
.B(n_188),
.Y(n_9234)
);

NAND2xp5_ASAP7_75t_SL g9235 ( 
.A(n_8536),
.B(n_188),
.Y(n_9235)
);

INVx1_ASAP7_75t_L g9236 ( 
.A(n_8715),
.Y(n_9236)
);

NOR2x2_ASAP7_75t_L g9237 ( 
.A(n_8580),
.B(n_188),
.Y(n_9237)
);

NAND2xp5_ASAP7_75t_SL g9238 ( 
.A(n_8629),
.B(n_189),
.Y(n_9238)
);

INVx3_ASAP7_75t_L g9239 ( 
.A(n_8448),
.Y(n_9239)
);

AOI22xp5_ASAP7_75t_L g9240 ( 
.A1(n_8901),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_9240)
);

NOR2x1_ASAP7_75t_R g9241 ( 
.A(n_8474),
.B(n_189),
.Y(n_9241)
);

INVx1_ASAP7_75t_L g9242 ( 
.A(n_8724),
.Y(n_9242)
);

INVx1_ASAP7_75t_L g9243 ( 
.A(n_8738),
.Y(n_9243)
);

BUFx2_ASAP7_75t_L g9244 ( 
.A(n_8855),
.Y(n_9244)
);

INVx2_ASAP7_75t_L g9245 ( 
.A(n_8482),
.Y(n_9245)
);

INVx1_ASAP7_75t_L g9246 ( 
.A(n_8739),
.Y(n_9246)
);

BUFx8_ASAP7_75t_L g9247 ( 
.A(n_8839),
.Y(n_9247)
);

NAND2xp5_ASAP7_75t_SL g9248 ( 
.A(n_8558),
.B(n_190),
.Y(n_9248)
);

AND2x2_ASAP7_75t_L g9249 ( 
.A(n_8613),
.B(n_190),
.Y(n_9249)
);

INVx1_ASAP7_75t_L g9250 ( 
.A(n_8740),
.Y(n_9250)
);

INVx2_ASAP7_75t_L g9251 ( 
.A(n_8483),
.Y(n_9251)
);

INVx2_ASAP7_75t_L g9252 ( 
.A(n_8488),
.Y(n_9252)
);

OR2x6_ASAP7_75t_L g9253 ( 
.A(n_8580),
.B(n_191),
.Y(n_9253)
);

AOI22xp33_ASAP7_75t_L g9254 ( 
.A1(n_8635),
.A2(n_195),
.B1(n_192),
.B2(n_194),
.Y(n_9254)
);

INVx4_ASAP7_75t_L g9255 ( 
.A(n_8646),
.Y(n_9255)
);

NAND2xp33_ASAP7_75t_SL g9256 ( 
.A(n_8571),
.B(n_192),
.Y(n_9256)
);

INVx2_ASAP7_75t_L g9257 ( 
.A(n_8494),
.Y(n_9257)
);

INVx1_ASAP7_75t_L g9258 ( 
.A(n_8741),
.Y(n_9258)
);

INVx2_ASAP7_75t_L g9259 ( 
.A(n_8908),
.Y(n_9259)
);

INVx1_ASAP7_75t_L g9260 ( 
.A(n_8743),
.Y(n_9260)
);

NAND2x1p5_ASAP7_75t_L g9261 ( 
.A(n_8677),
.B(n_192),
.Y(n_9261)
);

INVx1_ASAP7_75t_L g9262 ( 
.A(n_8760),
.Y(n_9262)
);

INVx5_ASAP7_75t_L g9263 ( 
.A(n_8604),
.Y(n_9263)
);

NAND2xp5_ASAP7_75t_L g9264 ( 
.A(n_8764),
.B(n_194),
.Y(n_9264)
);

INVx1_ASAP7_75t_L g9265 ( 
.A(n_8779),
.Y(n_9265)
);

INVx3_ASAP7_75t_L g9266 ( 
.A(n_8752),
.Y(n_9266)
);

AND2x2_ASAP7_75t_L g9267 ( 
.A(n_8731),
.B(n_194),
.Y(n_9267)
);

OAI21xp5_ASAP7_75t_L g9268 ( 
.A1(n_8649),
.A2(n_196),
.B(n_197),
.Y(n_9268)
);

INVx2_ASAP7_75t_L g9269 ( 
.A(n_8912),
.Y(n_9269)
);

NAND2xp5_ASAP7_75t_L g9270 ( 
.A(n_8789),
.B(n_196),
.Y(n_9270)
);

INVx1_ASAP7_75t_L g9271 ( 
.A(n_8792),
.Y(n_9271)
);

INVx2_ASAP7_75t_L g9272 ( 
.A(n_8653),
.Y(n_9272)
);

NOR2x2_ASAP7_75t_L g9273 ( 
.A(n_8959),
.B(n_196),
.Y(n_9273)
);

AND2x4_ASAP7_75t_L g9274 ( 
.A(n_8644),
.B(n_198),
.Y(n_9274)
);

INVx1_ASAP7_75t_L g9275 ( 
.A(n_8804),
.Y(n_9275)
);

INVx2_ASAP7_75t_SL g9276 ( 
.A(n_8671),
.Y(n_9276)
);

INVx2_ASAP7_75t_SL g9277 ( 
.A(n_8686),
.Y(n_9277)
);

INVxp67_ASAP7_75t_SL g9278 ( 
.A(n_8936),
.Y(n_9278)
);

INVx1_ASAP7_75t_L g9279 ( 
.A(n_8807),
.Y(n_9279)
);

NAND2xp5_ASAP7_75t_SL g9280 ( 
.A(n_8475),
.B(n_198),
.Y(n_9280)
);

INVx1_ASAP7_75t_L g9281 ( 
.A(n_8816),
.Y(n_9281)
);

NOR2xp33_ASAP7_75t_L g9282 ( 
.A(n_8572),
.B(n_198),
.Y(n_9282)
);

OAI22xp33_ASAP7_75t_L g9283 ( 
.A1(n_8595),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_9283)
);

BUFx4f_ASAP7_75t_L g9284 ( 
.A(n_8735),
.Y(n_9284)
);

INVx1_ASAP7_75t_SL g9285 ( 
.A(n_8744),
.Y(n_9285)
);

INVxp67_ASAP7_75t_L g9286 ( 
.A(n_8497),
.Y(n_9286)
);

BUFx12f_ASAP7_75t_L g9287 ( 
.A(n_8702),
.Y(n_9287)
);

INVx1_ASAP7_75t_L g9288 ( 
.A(n_8821),
.Y(n_9288)
);

NOR2xp33_ASAP7_75t_L g9289 ( 
.A(n_9008),
.B(n_8522),
.Y(n_9289)
);

INVx1_ASAP7_75t_L g9290 ( 
.A(n_8838),
.Y(n_9290)
);

AND2x6_ASAP7_75t_L g9291 ( 
.A(n_8858),
.B(n_199),
.Y(n_9291)
);

NAND2xp5_ASAP7_75t_L g9292 ( 
.A(n_8890),
.B(n_199),
.Y(n_9292)
);

NAND2xp5_ASAP7_75t_SL g9293 ( 
.A(n_8543),
.B(n_200),
.Y(n_9293)
);

INVx1_ASAP7_75t_SL g9294 ( 
.A(n_8750),
.Y(n_9294)
);

INVx2_ASAP7_75t_L g9295 ( 
.A(n_8655),
.Y(n_9295)
);

AOI22xp33_ASAP7_75t_L g9296 ( 
.A1(n_8710),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_9296)
);

INVx1_ASAP7_75t_L g9297 ( 
.A(n_8904),
.Y(n_9297)
);

NAND2xp5_ASAP7_75t_L g9298 ( 
.A(n_8963),
.B(n_201),
.Y(n_9298)
);

INVx1_ASAP7_75t_L g9299 ( 
.A(n_8906),
.Y(n_9299)
);

HB1xp67_ASAP7_75t_L g9300 ( 
.A(n_8918),
.Y(n_9300)
);

INVx1_ASAP7_75t_L g9301 ( 
.A(n_8929),
.Y(n_9301)
);

AOI21xp5_ASAP7_75t_L g9302 ( 
.A1(n_8541),
.A2(n_8524),
.B(n_8570),
.Y(n_9302)
);

INVx2_ASAP7_75t_L g9303 ( 
.A(n_8673),
.Y(n_9303)
);

NAND3xp33_ASAP7_75t_SL g9304 ( 
.A(n_8630),
.B(n_8637),
.C(n_8631),
.Y(n_9304)
);

INVx1_ASAP7_75t_L g9305 ( 
.A(n_8410),
.Y(n_9305)
);

NAND2xp5_ASAP7_75t_L g9306 ( 
.A(n_8496),
.B(n_202),
.Y(n_9306)
);

NAND2xp5_ASAP7_75t_L g9307 ( 
.A(n_8503),
.B(n_202),
.Y(n_9307)
);

NAND2xp5_ASAP7_75t_L g9308 ( 
.A(n_8505),
.B(n_203),
.Y(n_9308)
);

INVx3_ASAP7_75t_L g9309 ( 
.A(n_8546),
.Y(n_9309)
);

AOI22xp33_ASAP7_75t_L g9310 ( 
.A1(n_9007),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_9310)
);

INVx1_ASAP7_75t_L g9311 ( 
.A(n_8943),
.Y(n_9311)
);

NAND2xp5_ASAP7_75t_L g9312 ( 
.A(n_8642),
.B(n_204),
.Y(n_9312)
);

AND2x2_ASAP7_75t_SL g9313 ( 
.A(n_8877),
.B(n_204),
.Y(n_9313)
);

INVx2_ASAP7_75t_L g9314 ( 
.A(n_8680),
.Y(n_9314)
);

INVx1_ASAP7_75t_L g9315 ( 
.A(n_8945),
.Y(n_9315)
);

INVx1_ASAP7_75t_L g9316 ( 
.A(n_8948),
.Y(n_9316)
);

INVx1_ASAP7_75t_L g9317 ( 
.A(n_8965),
.Y(n_9317)
);

INVx1_ASAP7_75t_L g9318 ( 
.A(n_8982),
.Y(n_9318)
);

NAND2xp5_ASAP7_75t_SL g9319 ( 
.A(n_8565),
.B(n_205),
.Y(n_9319)
);

BUFx6f_ASAP7_75t_L g9320 ( 
.A(n_8754),
.Y(n_9320)
);

AOI22xp33_ASAP7_75t_L g9321 ( 
.A1(n_8634),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_8998),
.Y(n_9322)
);

NAND2xp33_ASAP7_75t_SL g9323 ( 
.A(n_8601),
.B(n_206),
.Y(n_9323)
);

AOI22xp5_ASAP7_75t_L g9324 ( 
.A1(n_8436),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_9324)
);

AOI22xp5_ASAP7_75t_L g9325 ( 
.A1(n_8625),
.A2(n_210),
.B1(n_207),
.B2(n_209),
.Y(n_9325)
);

INVx2_ASAP7_75t_SL g9326 ( 
.A(n_8859),
.Y(n_9326)
);

INVx1_ASAP7_75t_L g9327 ( 
.A(n_9012),
.Y(n_9327)
);

AND2x4_ASAP7_75t_SL g9328 ( 
.A(n_9015),
.B(n_8959),
.Y(n_9328)
);

INVx1_ASAP7_75t_L g9329 ( 
.A(n_8682),
.Y(n_9329)
);

AOI22xp5_ASAP7_75t_L g9330 ( 
.A1(n_8531),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_9330)
);

AND3x1_ASAP7_75t_SL g9331 ( 
.A(n_8705),
.B(n_211),
.C(n_212),
.Y(n_9331)
);

AOI22xp33_ASAP7_75t_L g9332 ( 
.A1(n_8633),
.A2(n_214),
.B1(n_211),
.B2(n_213),
.Y(n_9332)
);

OAI22xp5_ASAP7_75t_L g9333 ( 
.A1(n_8555),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_9333)
);

INVx1_ASAP7_75t_L g9334 ( 
.A(n_8689),
.Y(n_9334)
);

AND2x4_ASAP7_75t_L g9335 ( 
.A(n_8775),
.B(n_216),
.Y(n_9335)
);

NOR2xp33_ASAP7_75t_L g9336 ( 
.A(n_8879),
.B(n_216),
.Y(n_9336)
);

INVx1_ASAP7_75t_L g9337 ( 
.A(n_8721),
.Y(n_9337)
);

INVx5_ASAP7_75t_L g9338 ( 
.A(n_8442),
.Y(n_9338)
);

BUFx2_ASAP7_75t_L g9339 ( 
.A(n_8790),
.Y(n_9339)
);

INVx2_ASAP7_75t_L g9340 ( 
.A(n_8723),
.Y(n_9340)
);

NAND2xp5_ASAP7_75t_L g9341 ( 
.A(n_8641),
.B(n_217),
.Y(n_9341)
);

NOR2x1_ASAP7_75t_L g9342 ( 
.A(n_8883),
.B(n_217),
.Y(n_9342)
);

CKINVDCx5p33_ASAP7_75t_R g9343 ( 
.A(n_8996),
.Y(n_9343)
);

INVx1_ASAP7_75t_L g9344 ( 
.A(n_8732),
.Y(n_9344)
);

AOI22xp5_ASAP7_75t_L g9345 ( 
.A1(n_9002),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_9345)
);

INVx2_ASAP7_75t_L g9346 ( 
.A(n_8942),
.Y(n_9346)
);

NAND2xp5_ASAP7_75t_L g9347 ( 
.A(n_8836),
.B(n_218),
.Y(n_9347)
);

NOR2xp33_ASAP7_75t_L g9348 ( 
.A(n_8564),
.B(n_218),
.Y(n_9348)
);

INVx1_ASAP7_75t_L g9349 ( 
.A(n_8944),
.Y(n_9349)
);

AND2x4_ASAP7_75t_SL g9350 ( 
.A(n_8911),
.B(n_219),
.Y(n_9350)
);

NAND2x1p5_ASAP7_75t_L g9351 ( 
.A(n_8810),
.B(n_219),
.Y(n_9351)
);

OAI22xp5_ASAP7_75t_L g9352 ( 
.A1(n_8781),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_9352)
);

AOI22xp5_ASAP7_75t_L g9353 ( 
.A1(n_8713),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_9353)
);

INVx1_ASAP7_75t_L g9354 ( 
.A(n_8953),
.Y(n_9354)
);

AND2x4_ASAP7_75t_L g9355 ( 
.A(n_8683),
.B(n_221),
.Y(n_9355)
);

HB1xp67_ASAP7_75t_L g9356 ( 
.A(n_9000),
.Y(n_9356)
);

INVx2_ASAP7_75t_L g9357 ( 
.A(n_8962),
.Y(n_9357)
);

AND2x2_ASAP7_75t_L g9358 ( 
.A(n_8737),
.B(n_222),
.Y(n_9358)
);

NOR2xp33_ASAP7_75t_R g9359 ( 
.A(n_8896),
.B(n_223),
.Y(n_9359)
);

NAND2xp5_ASAP7_75t_L g9360 ( 
.A(n_8843),
.B(n_223),
.Y(n_9360)
);

INVx5_ASAP7_75t_L g9361 ( 
.A(n_8888),
.Y(n_9361)
);

A2O1A1Ixp33_ASAP7_75t_L g9362 ( 
.A1(n_8534),
.A2(n_226),
.B(n_224),
.C(n_225),
.Y(n_9362)
);

INVx1_ASAP7_75t_L g9363 ( 
.A(n_8967),
.Y(n_9363)
);

AND2x6_ASAP7_75t_L g9364 ( 
.A(n_8979),
.B(n_224),
.Y(n_9364)
);

INVx1_ASAP7_75t_L g9365 ( 
.A(n_8986),
.Y(n_9365)
);

NAND2xp5_ASAP7_75t_L g9366 ( 
.A(n_8582),
.B(n_224),
.Y(n_9366)
);

INVx4_ASAP7_75t_L g9367 ( 
.A(n_8920),
.Y(n_9367)
);

NOR3xp33_ASAP7_75t_SL g9368 ( 
.A(n_8711),
.B(n_225),
.C(n_226),
.Y(n_9368)
);

BUFx2_ASAP7_75t_L g9369 ( 
.A(n_8824),
.Y(n_9369)
);

INVx3_ASAP7_75t_L g9370 ( 
.A(n_8993),
.Y(n_9370)
);

NAND2xp5_ASAP7_75t_SL g9371 ( 
.A(n_8578),
.B(n_227),
.Y(n_9371)
);

INVx2_ASAP7_75t_SL g9372 ( 
.A(n_8457),
.Y(n_9372)
);

AOI22xp33_ASAP7_75t_L g9373 ( 
.A1(n_8672),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_9373)
);

NOR2xp33_ASAP7_75t_L g9374 ( 
.A(n_8960),
.B(n_228),
.Y(n_9374)
);

OAI22xp5_ASAP7_75t_L g9375 ( 
.A1(n_8793),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_9375)
);

BUFx2_ASAP7_75t_L g9376 ( 
.A(n_8829),
.Y(n_9376)
);

INVx2_ASAP7_75t_L g9377 ( 
.A(n_8999),
.Y(n_9377)
);

NAND2xp5_ASAP7_75t_L g9378 ( 
.A(n_8463),
.B(n_229),
.Y(n_9378)
);

OAI22xp5_ASAP7_75t_L g9379 ( 
.A1(n_8610),
.A2(n_8872),
.B1(n_8941),
.B2(n_8822),
.Y(n_9379)
);

BUFx3_ASAP7_75t_L g9380 ( 
.A(n_8473),
.Y(n_9380)
);

AOI22xp33_ASAP7_75t_L g9381 ( 
.A1(n_8956),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_9381)
);

NAND2xp5_ASAP7_75t_SL g9382 ( 
.A(n_8568),
.B(n_231),
.Y(n_9382)
);

OAI22xp5_ASAP7_75t_L g9383 ( 
.A1(n_8782),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_9383)
);

OR2x2_ASAP7_75t_L g9384 ( 
.A(n_8970),
.B(n_232),
.Y(n_9384)
);

INVx2_ASAP7_75t_SL g9385 ( 
.A(n_8479),
.Y(n_9385)
);

AND2x2_ASAP7_75t_L g9386 ( 
.A(n_8756),
.B(n_234),
.Y(n_9386)
);

OAI21xp33_ASAP7_75t_L g9387 ( 
.A1(n_8771),
.A2(n_234),
.B(n_235),
.Y(n_9387)
);

INVx3_ASAP7_75t_L g9388 ( 
.A(n_9009),
.Y(n_9388)
);

BUFx3_ASAP7_75t_L g9389 ( 
.A(n_8490),
.Y(n_9389)
);

INVx2_ASAP7_75t_L g9390 ( 
.A(n_8500),
.Y(n_9390)
);

NOR3xp33_ASAP7_75t_L g9391 ( 
.A(n_8757),
.B(n_234),
.C(n_235),
.Y(n_9391)
);

AOI22xp5_ASAP7_75t_L g9392 ( 
.A1(n_8770),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_9392)
);

INVx3_ASAP7_75t_L g9393 ( 
.A(n_9010),
.Y(n_9393)
);

INVx1_ASAP7_75t_L g9394 ( 
.A(n_8930),
.Y(n_9394)
);

NOR2xp33_ASAP7_75t_SL g9395 ( 
.A(n_8520),
.B(n_236),
.Y(n_9395)
);

AOI22xp33_ASAP7_75t_L g9396 ( 
.A1(n_8957),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_9396)
);

INVx2_ASAP7_75t_L g9397 ( 
.A(n_8504),
.Y(n_9397)
);

INVx1_ASAP7_75t_L g9398 ( 
.A(n_8933),
.Y(n_9398)
);

NAND2xp5_ASAP7_75t_L g9399 ( 
.A(n_8507),
.B(n_237),
.Y(n_9399)
);

HB1xp67_ASAP7_75t_L g9400 ( 
.A(n_8882),
.Y(n_9400)
);

NAND2xp5_ASAP7_75t_SL g9401 ( 
.A(n_8576),
.B(n_238),
.Y(n_9401)
);

INVx2_ASAP7_75t_L g9402 ( 
.A(n_8510),
.Y(n_9402)
);

INVx5_ASAP7_75t_L g9403 ( 
.A(n_8823),
.Y(n_9403)
);

AND2x6_ASAP7_75t_SL g9404 ( 
.A(n_8977),
.B(n_8987),
.Y(n_9404)
);

INVx2_ASAP7_75t_SL g9405 ( 
.A(n_8777),
.Y(n_9405)
);

BUFx3_ASAP7_75t_L g9406 ( 
.A(n_8867),
.Y(n_9406)
);

INVx3_ASAP7_75t_L g9407 ( 
.A(n_8746),
.Y(n_9407)
);

INVx2_ASAP7_75t_L g9408 ( 
.A(n_8762),
.Y(n_9408)
);

CKINVDCx5p33_ASAP7_75t_R g9409 ( 
.A(n_8915),
.Y(n_9409)
);

BUFx6f_ASAP7_75t_L g9410 ( 
.A(n_8492),
.Y(n_9410)
);

INVx2_ASAP7_75t_L g9411 ( 
.A(n_8812),
.Y(n_9411)
);

INVx2_ASAP7_75t_L g9412 ( 
.A(n_8830),
.Y(n_9412)
);

INVx1_ASAP7_75t_L g9413 ( 
.A(n_8847),
.Y(n_9413)
);

AOI21xp5_ASAP7_75t_L g9414 ( 
.A1(n_8669),
.A2(n_238),
.B(n_239),
.Y(n_9414)
);

NAND3xp33_ASAP7_75t_SL g9415 ( 
.A(n_8907),
.B(n_239),
.C(n_240),
.Y(n_9415)
);

NAND2xp5_ASAP7_75t_L g9416 ( 
.A(n_8608),
.B(n_239),
.Y(n_9416)
);

AND2x2_ASAP7_75t_L g9417 ( 
.A(n_8798),
.B(n_241),
.Y(n_9417)
);

INVx1_ASAP7_75t_L g9418 ( 
.A(n_8853),
.Y(n_9418)
);

INVx2_ASAP7_75t_L g9419 ( 
.A(n_8856),
.Y(n_9419)
);

INVx3_ASAP7_75t_L g9420 ( 
.A(n_8857),
.Y(n_9420)
);

BUFx3_ASAP7_75t_L g9421 ( 
.A(n_8697),
.Y(n_9421)
);

INVx1_ASAP7_75t_L g9422 ( 
.A(n_8863),
.Y(n_9422)
);

NAND2xp33_ASAP7_75t_L g9423 ( 
.A(n_8786),
.B(n_241),
.Y(n_9423)
);

O2A1O1Ixp33_ASAP7_75t_L g9424 ( 
.A1(n_8605),
.A2(n_243),
.B(n_241),
.C(n_242),
.Y(n_9424)
);

INVx2_ASAP7_75t_L g9425 ( 
.A(n_8865),
.Y(n_9425)
);

AOI22xp33_ASAP7_75t_L g9426 ( 
.A1(n_8827),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_9426)
);

INVx1_ASAP7_75t_L g9427 ( 
.A(n_8868),
.Y(n_9427)
);

BUFx3_ASAP7_75t_L g9428 ( 
.A(n_8801),
.Y(n_9428)
);

INVx2_ASAP7_75t_L g9429 ( 
.A(n_8870),
.Y(n_9429)
);

NOR2xp33_ASAP7_75t_L g9430 ( 
.A(n_8961),
.B(n_242),
.Y(n_9430)
);

NOR3xp33_ASAP7_75t_L g9431 ( 
.A(n_8733),
.B(n_244),
.C(n_245),
.Y(n_9431)
);

NOR2xp33_ASAP7_75t_R g9432 ( 
.A(n_8585),
.B(n_244),
.Y(n_9432)
);

HB1xp67_ASAP7_75t_L g9433 ( 
.A(n_8894),
.Y(n_9433)
);

OAI22xp5_ASAP7_75t_SL g9434 ( 
.A1(n_8846),
.A2(n_8990),
.B1(n_8992),
.B2(n_8783),
.Y(n_9434)
);

INVx2_ASAP7_75t_L g9435 ( 
.A(n_8887),
.Y(n_9435)
);

INVxp67_ASAP7_75t_L g9436 ( 
.A(n_8840),
.Y(n_9436)
);

INVx2_ASAP7_75t_L g9437 ( 
.A(n_8891),
.Y(n_9437)
);

INVx2_ASAP7_75t_L g9438 ( 
.A(n_8902),
.Y(n_9438)
);

NAND2x1p5_ASAP7_75t_L g9439 ( 
.A(n_8450),
.B(n_245),
.Y(n_9439)
);

CKINVDCx5p33_ASAP7_75t_R g9440 ( 
.A(n_8586),
.Y(n_9440)
);

A2O1A1Ixp33_ASAP7_75t_L g9441 ( 
.A1(n_8668),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_9441)
);

INVx1_ASAP7_75t_L g9442 ( 
.A(n_8934),
.Y(n_9442)
);

AND2x4_ASAP7_75t_L g9443 ( 
.A(n_8589),
.B(n_246),
.Y(n_9443)
);

INVx5_ASAP7_75t_L g9444 ( 
.A(n_8811),
.Y(n_9444)
);

NOR3xp33_ASAP7_75t_SL g9445 ( 
.A(n_8632),
.B(n_247),
.C(n_248),
.Y(n_9445)
);

NAND2xp5_ASAP7_75t_L g9446 ( 
.A(n_8897),
.B(n_247),
.Y(n_9446)
);

INVxp67_ASAP7_75t_L g9447 ( 
.A(n_8593),
.Y(n_9447)
);

INVx1_ASAP7_75t_L g9448 ( 
.A(n_9006),
.Y(n_9448)
);

BUFx3_ASAP7_75t_L g9449 ( 
.A(n_9003),
.Y(n_9449)
);

AOI22xp5_ASAP7_75t_L g9450 ( 
.A1(n_8785),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_9450)
);

INVx1_ASAP7_75t_L g9451 ( 
.A(n_8926),
.Y(n_9451)
);

INVx1_ASAP7_75t_L g9452 ( 
.A(n_8954),
.Y(n_9452)
);

INVx1_ASAP7_75t_L g9453 ( 
.A(n_8958),
.Y(n_9453)
);

AOI22xp5_ASAP7_75t_L g9454 ( 
.A1(n_8819),
.A2(n_251),
.B1(n_248),
.B2(n_249),
.Y(n_9454)
);

AOI21xp5_ASAP7_75t_L g9455 ( 
.A1(n_8678),
.A2(n_252),
.B(n_253),
.Y(n_9455)
);

INVx1_ASAP7_75t_L g9456 ( 
.A(n_8964),
.Y(n_9456)
);

NAND2xp5_ASAP7_75t_SL g9457 ( 
.A(n_8831),
.B(n_252),
.Y(n_9457)
);

INVx1_ASAP7_75t_L g9458 ( 
.A(n_8966),
.Y(n_9458)
);

BUFx4f_ASAP7_75t_L g9459 ( 
.A(n_8989),
.Y(n_9459)
);

INVx1_ASAP7_75t_L g9460 ( 
.A(n_8969),
.Y(n_9460)
);

BUFx6f_ASAP7_75t_L g9461 ( 
.A(n_8465),
.Y(n_9461)
);

NAND2xp5_ASAP7_75t_SL g9462 ( 
.A(n_8833),
.B(n_252),
.Y(n_9462)
);

AND2x2_ASAP7_75t_L g9463 ( 
.A(n_8849),
.B(n_253),
.Y(n_9463)
);

NAND2xp5_ASAP7_75t_L g9464 ( 
.A(n_8884),
.B(n_253),
.Y(n_9464)
);

BUFx6f_ASAP7_75t_L g9465 ( 
.A(n_8742),
.Y(n_9465)
);

NOR2xp33_ASAP7_75t_L g9466 ( 
.A(n_8871),
.B(n_254),
.Y(n_9466)
);

INVx2_ASAP7_75t_L g9467 ( 
.A(n_8947),
.Y(n_9467)
);

INVx3_ASAP7_75t_L g9468 ( 
.A(n_8618),
.Y(n_9468)
);

BUFx4f_ASAP7_75t_L g9469 ( 
.A(n_8714),
.Y(n_9469)
);

INVxp67_ASAP7_75t_SL g9470 ( 
.A(n_8850),
.Y(n_9470)
);

NOR2x2_ASAP7_75t_L g9471 ( 
.A(n_8841),
.B(n_254),
.Y(n_9471)
);

INVx1_ASAP7_75t_L g9472 ( 
.A(n_8975),
.Y(n_9472)
);

BUFx3_ASAP7_75t_L g9473 ( 
.A(n_8716),
.Y(n_9473)
);

INVx4_ASAP7_75t_L g9474 ( 
.A(n_8917),
.Y(n_9474)
);

AND2x4_ASAP7_75t_L g9475 ( 
.A(n_8602),
.B(n_255),
.Y(n_9475)
);

OR2x6_ASAP7_75t_L g9476 ( 
.A(n_8828),
.B(n_255),
.Y(n_9476)
);

INVx3_ASAP7_75t_L g9477 ( 
.A(n_8949),
.Y(n_9477)
);

NAND2xp5_ASAP7_75t_L g9478 ( 
.A(n_8895),
.B(n_256),
.Y(n_9478)
);

NAND2xp5_ASAP7_75t_L g9479 ( 
.A(n_8837),
.B(n_8645),
.Y(n_9479)
);

NOR2x1_ASAP7_75t_L g9480 ( 
.A(n_8919),
.B(n_8658),
.Y(n_9480)
);

HB1xp67_ASAP7_75t_L g9481 ( 
.A(n_8976),
.Y(n_9481)
);

INVx2_ASAP7_75t_L g9482 ( 
.A(n_8978),
.Y(n_9482)
);

AOI22xp33_ASAP7_75t_SL g9483 ( 
.A1(n_8910),
.A2(n_8815),
.B1(n_8984),
.B2(n_8780),
.Y(n_9483)
);

INVx1_ASAP7_75t_L g9484 ( 
.A(n_8983),
.Y(n_9484)
);

NAND2xp5_ASAP7_75t_L g9485 ( 
.A(n_8652),
.B(n_256),
.Y(n_9485)
);

INVx1_ASAP7_75t_L g9486 ( 
.A(n_8994),
.Y(n_9486)
);

AOI22xp33_ASAP7_75t_L g9487 ( 
.A1(n_9005),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_9487)
);

AOI21xp5_ASAP7_75t_L g9488 ( 
.A1(n_8687),
.A2(n_257),
.B(n_258),
.Y(n_9488)
);

INVx1_ASAP7_75t_L g9489 ( 
.A(n_8997),
.Y(n_9489)
);

NAND2xp5_ASAP7_75t_L g9490 ( 
.A(n_8659),
.B(n_258),
.Y(n_9490)
);

BUFx2_ASAP7_75t_L g9491 ( 
.A(n_9011),
.Y(n_9491)
);

NAND3xp33_ASAP7_75t_SL g9492 ( 
.A(n_8844),
.B(n_259),
.C(n_260),
.Y(n_9492)
);

NOR2x1p5_ASAP7_75t_L g9493 ( 
.A(n_8662),
.B(n_260),
.Y(n_9493)
);

INVx2_ASAP7_75t_L g9494 ( 
.A(n_9013),
.Y(n_9494)
);

NAND2xp5_ASAP7_75t_L g9495 ( 
.A(n_8663),
.B(n_260),
.Y(n_9495)
);

INVx2_ASAP7_75t_SL g9496 ( 
.A(n_8922),
.Y(n_9496)
);

INVxp67_ASAP7_75t_L g9497 ( 
.A(n_8609),
.Y(n_9497)
);

NAND2xp33_ASAP7_75t_L g9498 ( 
.A(n_8751),
.B(n_261),
.Y(n_9498)
);

BUFx3_ASAP7_75t_L g9499 ( 
.A(n_8722),
.Y(n_9499)
);

NAND2xp5_ASAP7_75t_SL g9500 ( 
.A(n_8937),
.B(n_261),
.Y(n_9500)
);

INVx2_ASAP7_75t_L g9501 ( 
.A(n_8914),
.Y(n_9501)
);

NAND2xp5_ASAP7_75t_L g9502 ( 
.A(n_8664),
.B(n_262),
.Y(n_9502)
);

A2O1A1Ixp33_ASAP7_75t_L g9503 ( 
.A1(n_8650),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_9503)
);

INVx1_ASAP7_75t_L g9504 ( 
.A(n_8916),
.Y(n_9504)
);

NAND2xp33_ASAP7_75t_L g9505 ( 
.A(n_8974),
.B(n_263),
.Y(n_9505)
);

BUFx3_ASAP7_75t_L g9506 ( 
.A(n_8794),
.Y(n_9506)
);

AND2x6_ASAP7_75t_SL g9507 ( 
.A(n_8626),
.B(n_8636),
.Y(n_9507)
);

NAND2xp5_ASAP7_75t_L g9508 ( 
.A(n_8674),
.B(n_263),
.Y(n_9508)
);

NOR3xp33_ASAP7_75t_L g9509 ( 
.A(n_8852),
.B(n_8835),
.C(n_8825),
.Y(n_9509)
);

OAI22xp5_ASAP7_75t_SL g9510 ( 
.A1(n_8886),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_9510)
);

NAND2xp5_ASAP7_75t_SL g9511 ( 
.A(n_8691),
.B(n_265),
.Y(n_9511)
);

NOR2xp33_ASAP7_75t_R g9512 ( 
.A(n_8688),
.B(n_266),
.Y(n_9512)
);

INVx2_ASAP7_75t_L g9513 ( 
.A(n_8923),
.Y(n_9513)
);

INVx1_ASAP7_75t_L g9514 ( 
.A(n_8924),
.Y(n_9514)
);

NAND2xp5_ASAP7_75t_L g9515 ( 
.A(n_8692),
.B(n_266),
.Y(n_9515)
);

NAND2xp5_ASAP7_75t_L g9516 ( 
.A(n_8698),
.B(n_267),
.Y(n_9516)
);

NAND2xp5_ASAP7_75t_SL g9517 ( 
.A(n_8694),
.B(n_268),
.Y(n_9517)
);

AND2x2_ASAP7_75t_L g9518 ( 
.A(n_8860),
.B(n_268),
.Y(n_9518)
);

INVx2_ASAP7_75t_L g9519 ( 
.A(n_8925),
.Y(n_9519)
);

INVx1_ASAP7_75t_L g9520 ( 
.A(n_8931),
.Y(n_9520)
);

BUFx2_ASAP7_75t_L g9521 ( 
.A(n_8932),
.Y(n_9521)
);

NAND2xp5_ASAP7_75t_L g9522 ( 
.A(n_8699),
.B(n_268),
.Y(n_9522)
);

NAND2xp5_ASAP7_75t_SL g9523 ( 
.A(n_8696),
.B(n_269),
.Y(n_9523)
);

INVx1_ASAP7_75t_L g9524 ( 
.A(n_8704),
.Y(n_9524)
);

INVx2_ASAP7_75t_SL g9525 ( 
.A(n_8991),
.Y(n_9525)
);

INVx1_ASAP7_75t_L g9526 ( 
.A(n_8717),
.Y(n_9526)
);

NAND2xp5_ASAP7_75t_L g9527 ( 
.A(n_8725),
.B(n_269),
.Y(n_9527)
);

INVx3_ASAP7_75t_L g9528 ( 
.A(n_8728),
.Y(n_9528)
);

NOR2xp33_ASAP7_75t_L g9529 ( 
.A(n_8755),
.B(n_269),
.Y(n_9529)
);

INVx2_ASAP7_75t_L g9530 ( 
.A(n_8734),
.Y(n_9530)
);

CKINVDCx5p33_ASAP7_75t_R g9531 ( 
.A(n_8758),
.Y(n_9531)
);

AND2x4_ASAP7_75t_L g9532 ( 
.A(n_8619),
.B(n_270),
.Y(n_9532)
);

INVx2_ASAP7_75t_L g9533 ( 
.A(n_8736),
.Y(n_9533)
);

NAND2xp5_ASAP7_75t_L g9534 ( 
.A(n_8745),
.B(n_8753),
.Y(n_9534)
);

AND2x4_ASAP7_75t_L g9535 ( 
.A(n_8562),
.B(n_270),
.Y(n_9535)
);

INVx1_ASAP7_75t_L g9536 ( 
.A(n_8761),
.Y(n_9536)
);

AOI22xp5_ASAP7_75t_L g9537 ( 
.A1(n_8820),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_9537)
);

BUFx3_ASAP7_75t_L g9538 ( 
.A(n_8766),
.Y(n_9538)
);

AND2x4_ASAP7_75t_L g9539 ( 
.A(n_8563),
.B(n_271),
.Y(n_9539)
);

INVx1_ASAP7_75t_L g9540 ( 
.A(n_8769),
.Y(n_9540)
);

INVx2_ASAP7_75t_L g9541 ( 
.A(n_8772),
.Y(n_9541)
);

INVx1_ASAP7_75t_L g9542 ( 
.A(n_8773),
.Y(n_9542)
);

INVx2_ASAP7_75t_L g9543 ( 
.A(n_8778),
.Y(n_9543)
);

AOI22xp5_ASAP7_75t_L g9544 ( 
.A1(n_8971),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_9544)
);

NAND2xp5_ASAP7_75t_L g9545 ( 
.A(n_8791),
.B(n_272),
.Y(n_9545)
);

NAND2xp5_ASAP7_75t_SL g9546 ( 
.A(n_8708),
.B(n_273),
.Y(n_9546)
);

AND2x2_ASAP7_75t_L g9547 ( 
.A(n_8800),
.B(n_273),
.Y(n_9547)
);

A2O1A1Ixp33_ASAP7_75t_SL g9548 ( 
.A1(n_8787),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_9548)
);

NAND2x1p5_ASAP7_75t_L g9549 ( 
.A(n_8712),
.B(n_274),
.Y(n_9549)
);

INVx2_ASAP7_75t_SL g9550 ( 
.A(n_8796),
.Y(n_9550)
);

NAND2xp5_ASAP7_75t_L g9551 ( 
.A(n_8797),
.B(n_275),
.Y(n_9551)
);

AND2x4_ASAP7_75t_L g9552 ( 
.A(n_9004),
.B(n_275),
.Y(n_9552)
);

INVx1_ASAP7_75t_L g9553 ( 
.A(n_8802),
.Y(n_9553)
);

NAND2xp5_ASAP7_75t_L g9554 ( 
.A(n_8803),
.B(n_276),
.Y(n_9554)
);

OAI22xp5_ASAP7_75t_L g9555 ( 
.A1(n_8747),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_9555)
);

INVx1_ASAP7_75t_L g9556 ( 
.A(n_8805),
.Y(n_9556)
);

INVx2_ASAP7_75t_L g9557 ( 
.A(n_8808),
.Y(n_9557)
);

INVx1_ASAP7_75t_L g9558 ( 
.A(n_8809),
.Y(n_9558)
);

AND2x4_ASAP7_75t_L g9559 ( 
.A(n_9014),
.B(n_277),
.Y(n_9559)
);

AOI22xp33_ASAP7_75t_L g9560 ( 
.A1(n_8935),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_9560)
);

AND2x4_ASAP7_75t_L g9561 ( 
.A(n_8938),
.B(n_278),
.Y(n_9561)
);

INVx1_ASAP7_75t_L g9562 ( 
.A(n_8817),
.Y(n_9562)
);

NAND2xp33_ASAP7_75t_L g9563 ( 
.A(n_8832),
.B(n_279),
.Y(n_9563)
);

NAND2xp5_ASAP7_75t_SL g9564 ( 
.A(n_8718),
.B(n_280),
.Y(n_9564)
);

NAND2xp5_ASAP7_75t_L g9565 ( 
.A(n_8861),
.B(n_280),
.Y(n_9565)
);

INVx1_ASAP7_75t_L g9566 ( 
.A(n_8864),
.Y(n_9566)
);

INVx1_ASAP7_75t_L g9567 ( 
.A(n_8873),
.Y(n_9567)
);

INVx1_ASAP7_75t_L g9568 ( 
.A(n_8874),
.Y(n_9568)
);

AOI22xp33_ASAP7_75t_L g9569 ( 
.A1(n_8985),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_9569)
);

OR2x6_ASAP7_75t_L g9570 ( 
.A(n_8851),
.B(n_281),
.Y(n_9570)
);

BUFx2_ASAP7_75t_L g9571 ( 
.A(n_8875),
.Y(n_9571)
);

NOR2xp33_ASAP7_75t_L g9572 ( 
.A(n_8774),
.B(n_281),
.Y(n_9572)
);

NAND2x1p5_ASAP7_75t_L g9573 ( 
.A(n_8719),
.B(n_283),
.Y(n_9573)
);

NAND2xp5_ASAP7_75t_L g9574 ( 
.A(n_8876),
.B(n_284),
.Y(n_9574)
);

AOI21xp5_ASAP7_75t_L g9575 ( 
.A1(n_8720),
.A2(n_285),
.B(n_286),
.Y(n_9575)
);

NOR2xp33_ASAP7_75t_L g9576 ( 
.A(n_8776),
.B(n_285),
.Y(n_9576)
);

AOI22xp5_ASAP7_75t_L g9577 ( 
.A1(n_8892),
.A2(n_288),
.B1(n_285),
.B2(n_287),
.Y(n_9577)
);

INVx3_ASAP7_75t_L g9578 ( 
.A(n_8878),
.Y(n_9578)
);

AND2x2_ASAP7_75t_L g9579 ( 
.A(n_8880),
.B(n_8893),
.Y(n_9579)
);

NAND2xp33_ASAP7_75t_L g9580 ( 
.A(n_8898),
.B(n_287),
.Y(n_9580)
);

INVx2_ASAP7_75t_SL g9581 ( 
.A(n_8905),
.Y(n_9581)
);

AOI22xp5_ASAP7_75t_L g9582 ( 
.A1(n_8623),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_9582)
);

NOR3xp33_ASAP7_75t_SL g9583 ( 
.A(n_8784),
.B(n_288),
.C(n_289),
.Y(n_9583)
);

BUFx6f_ASAP7_75t_L g9584 ( 
.A(n_8627),
.Y(n_9584)
);

NAND2xp5_ASAP7_75t_SL g9585 ( 
.A(n_8862),
.B(n_290),
.Y(n_9585)
);

INVx2_ASAP7_75t_SL g9586 ( 
.A(n_8795),
.Y(n_9586)
);

INVx1_ASAP7_75t_L g9587 ( 
.A(n_8939),
.Y(n_9587)
);

INVx1_ASAP7_75t_L g9588 ( 
.A(n_8940),
.Y(n_9588)
);

BUFx2_ASAP7_75t_L g9589 ( 
.A(n_8952),
.Y(n_9589)
);

O2A1O1Ixp33_ASAP7_75t_L g9590 ( 
.A1(n_8913),
.A2(n_8729),
.B(n_8889),
.C(n_8981),
.Y(n_9590)
);

INVx1_ASAP7_75t_L g9591 ( 
.A(n_8927),
.Y(n_9591)
);

AND3x1_ASAP7_75t_L g9592 ( 
.A(n_8988),
.B(n_290),
.C(n_291),
.Y(n_9592)
);

NAND2xp5_ASAP7_75t_SL g9593 ( 
.A(n_8995),
.B(n_291),
.Y(n_9593)
);

BUFx6f_ASAP7_75t_L g9594 ( 
.A(n_8654),
.Y(n_9594)
);

NAND2xp5_ASAP7_75t_L g9595 ( 
.A(n_8588),
.B(n_291),
.Y(n_9595)
);

INVx1_ASAP7_75t_L g9596 ( 
.A(n_8690),
.Y(n_9596)
);

INVx1_ASAP7_75t_L g9597 ( 
.A(n_8690),
.Y(n_9597)
);

INVx2_ASAP7_75t_SL g9598 ( 
.A(n_8654),
.Y(n_9598)
);

NAND2xp5_ASAP7_75t_SL g9599 ( 
.A(n_8419),
.B(n_292),
.Y(n_9599)
);

BUFx4f_ASAP7_75t_SL g9600 ( 
.A(n_8431),
.Y(n_9600)
);

INVx2_ASAP7_75t_L g9601 ( 
.A(n_8528),
.Y(n_9601)
);

INVx2_ASAP7_75t_L g9602 ( 
.A(n_8528),
.Y(n_9602)
);

NOR2xp33_ASAP7_75t_L g9603 ( 
.A(n_8419),
.B(n_292),
.Y(n_9603)
);

XOR2xp5_ASAP7_75t_L g9604 ( 
.A(n_9033),
.B(n_292),
.Y(n_9604)
);

NAND2xp5_ASAP7_75t_L g9605 ( 
.A(n_9095),
.B(n_9017),
.Y(n_9605)
);

NOR2xp33_ASAP7_75t_L g9606 ( 
.A(n_9164),
.B(n_293),
.Y(n_9606)
);

NAND2xp33_ASAP7_75t_L g9607 ( 
.A(n_9213),
.B(n_293),
.Y(n_9607)
);

NAND2xp5_ASAP7_75t_L g9608 ( 
.A(n_9019),
.B(n_293),
.Y(n_9608)
);

A2O1A1Ixp33_ASAP7_75t_L g9609 ( 
.A1(n_9107),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_9609)
);

INVx1_ASAP7_75t_SL g9610 ( 
.A(n_9226),
.Y(n_9610)
);

NAND2xp5_ASAP7_75t_L g9611 ( 
.A(n_9031),
.B(n_294),
.Y(n_9611)
);

CKINVDCx10_ASAP7_75t_R g9612 ( 
.A(n_9114),
.Y(n_9612)
);

AOI21x1_ASAP7_75t_L g9613 ( 
.A1(n_9028),
.A2(n_294),
.B(n_295),
.Y(n_9613)
);

OAI22xp5_ASAP7_75t_SL g9614 ( 
.A1(n_9253),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_9614)
);

BUFx8_ASAP7_75t_L g9615 ( 
.A(n_9120),
.Y(n_9615)
);

INVx2_ASAP7_75t_L g9616 ( 
.A(n_9049),
.Y(n_9616)
);

OAI22xp5_ASAP7_75t_L g9617 ( 
.A1(n_9483),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_9617)
);

NOR3xp33_ASAP7_75t_L g9618 ( 
.A(n_9293),
.B(n_297),
.C(n_298),
.Y(n_9618)
);

INVx1_ASAP7_75t_L g9619 ( 
.A(n_9190),
.Y(n_9619)
);

AOI21x1_ASAP7_75t_L g9620 ( 
.A1(n_9172),
.A2(n_9202),
.B(n_9048),
.Y(n_9620)
);

BUFx4f_ASAP7_75t_L g9621 ( 
.A(n_9594),
.Y(n_9621)
);

BUFx6f_ASAP7_75t_L g9622 ( 
.A(n_9594),
.Y(n_9622)
);

NAND2xp5_ASAP7_75t_L g9623 ( 
.A(n_9037),
.B(n_298),
.Y(n_9623)
);

NAND3xp33_ASAP7_75t_L g9624 ( 
.A(n_9065),
.B(n_299),
.C(n_300),
.Y(n_9624)
);

OR2x2_ASAP7_75t_L g9625 ( 
.A(n_9149),
.B(n_299),
.Y(n_9625)
);

INVx2_ASAP7_75t_L g9626 ( 
.A(n_9601),
.Y(n_9626)
);

NAND2xp5_ASAP7_75t_L g9627 ( 
.A(n_9062),
.B(n_300),
.Y(n_9627)
);

NAND2xp5_ASAP7_75t_L g9628 ( 
.A(n_9068),
.B(n_9596),
.Y(n_9628)
);

OAI22xp5_ASAP7_75t_L g9629 ( 
.A1(n_9130),
.A2(n_9089),
.B1(n_9454),
.B2(n_9450),
.Y(n_9629)
);

INVx1_ASAP7_75t_L g9630 ( 
.A(n_9300),
.Y(n_9630)
);

AOI21xp5_ASAP7_75t_L g9631 ( 
.A1(n_9030),
.A2(n_300),
.B(n_301),
.Y(n_9631)
);

O2A1O1Ixp33_ASAP7_75t_L g9632 ( 
.A1(n_9423),
.A2(n_303),
.B(n_301),
.C(n_302),
.Y(n_9632)
);

AOI22xp33_ASAP7_75t_L g9633 ( 
.A1(n_9141),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_9633)
);

BUFx3_ASAP7_75t_L g9634 ( 
.A(n_9066),
.Y(n_9634)
);

NAND2xp5_ASAP7_75t_L g9635 ( 
.A(n_9597),
.B(n_302),
.Y(n_9635)
);

AOI21xp5_ASAP7_75t_L g9636 ( 
.A1(n_9136),
.A2(n_304),
.B(n_305),
.Y(n_9636)
);

BUFx3_ASAP7_75t_L g9637 ( 
.A(n_9066),
.Y(n_9637)
);

NAND2xp5_ASAP7_75t_L g9638 ( 
.A(n_9108),
.B(n_304),
.Y(n_9638)
);

INVx2_ASAP7_75t_L g9639 ( 
.A(n_9602),
.Y(n_9639)
);

AOI21x1_ASAP7_75t_L g9640 ( 
.A1(n_9125),
.A2(n_305),
.B(n_306),
.Y(n_9640)
);

OAI21xp5_ASAP7_75t_L g9641 ( 
.A1(n_9175),
.A2(n_305),
.B(n_306),
.Y(n_9641)
);

NAND2xp5_ASAP7_75t_SL g9642 ( 
.A(n_9143),
.B(n_307),
.Y(n_9642)
);

NAND2xp5_ASAP7_75t_SL g9643 ( 
.A(n_9143),
.B(n_307),
.Y(n_9643)
);

AOI21xp5_ASAP7_75t_L g9644 ( 
.A1(n_9278),
.A2(n_307),
.B(n_308),
.Y(n_9644)
);

NAND2xp5_ASAP7_75t_L g9645 ( 
.A(n_9016),
.B(n_9380),
.Y(n_9645)
);

BUFx6f_ASAP7_75t_L g9646 ( 
.A(n_9284),
.Y(n_9646)
);

NAND2xp33_ASAP7_75t_L g9647 ( 
.A(n_9213),
.B(n_308),
.Y(n_9647)
);

INVx1_ASAP7_75t_L g9648 ( 
.A(n_9087),
.Y(n_9648)
);

NAND2xp5_ASAP7_75t_L g9649 ( 
.A(n_9389),
.B(n_308),
.Y(n_9649)
);

AOI21xp5_ASAP7_75t_L g9650 ( 
.A1(n_9302),
.A2(n_309),
.B(n_310),
.Y(n_9650)
);

OAI22xp5_ASAP7_75t_L g9651 ( 
.A1(n_9603),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_9651)
);

AOI21xp5_ASAP7_75t_L g9652 ( 
.A1(n_9590),
.A2(n_309),
.B(n_310),
.Y(n_9652)
);

AOI21xp5_ASAP7_75t_L g9653 ( 
.A1(n_9387),
.A2(n_312),
.B(n_313),
.Y(n_9653)
);

AOI21x1_ASAP7_75t_L g9654 ( 
.A1(n_9127),
.A2(n_312),
.B(n_313),
.Y(n_9654)
);

NAND2xp5_ASAP7_75t_L g9655 ( 
.A(n_9070),
.B(n_312),
.Y(n_9655)
);

NAND2xp5_ASAP7_75t_L g9656 ( 
.A(n_9093),
.B(n_313),
.Y(n_9656)
);

BUFx3_ASAP7_75t_L g9657 ( 
.A(n_9101),
.Y(n_9657)
);

INVx2_ASAP7_75t_L g9658 ( 
.A(n_9053),
.Y(n_9658)
);

NAND2xp5_ASAP7_75t_L g9659 ( 
.A(n_9174),
.B(n_314),
.Y(n_9659)
);

NAND2xp5_ASAP7_75t_L g9660 ( 
.A(n_9356),
.B(n_314),
.Y(n_9660)
);

AOI21xp5_ASAP7_75t_L g9661 ( 
.A1(n_9215),
.A2(n_315),
.B(n_316),
.Y(n_9661)
);

NAND2xp5_ASAP7_75t_L g9662 ( 
.A(n_9024),
.B(n_9025),
.Y(n_9662)
);

AOI21xp5_ASAP7_75t_L g9663 ( 
.A1(n_9153),
.A2(n_315),
.B(n_316),
.Y(n_9663)
);

NAND2xp5_ASAP7_75t_L g9664 ( 
.A(n_9372),
.B(n_316),
.Y(n_9664)
);

AOI22xp5_ASAP7_75t_L g9665 ( 
.A1(n_9213),
.A2(n_320),
.B1(n_317),
.B2(n_318),
.Y(n_9665)
);

AND2x2_ASAP7_75t_L g9666 ( 
.A(n_9468),
.B(n_317),
.Y(n_9666)
);

NAND2xp5_ASAP7_75t_L g9667 ( 
.A(n_9385),
.B(n_320),
.Y(n_9667)
);

OAI22xp5_ASAP7_75t_L g9668 ( 
.A1(n_9204),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_9668)
);

AOI21xp5_ASAP7_75t_L g9669 ( 
.A1(n_9123),
.A2(n_321),
.B(n_322),
.Y(n_9669)
);

NAND2xp5_ASAP7_75t_L g9670 ( 
.A(n_9400),
.B(n_322),
.Y(n_9670)
);

HB1xp67_ASAP7_75t_L g9671 ( 
.A(n_9433),
.Y(n_9671)
);

AOI21xp5_ASAP7_75t_L g9672 ( 
.A1(n_9029),
.A2(n_323),
.B(n_324),
.Y(n_9672)
);

AO32x1_ASAP7_75t_L g9673 ( 
.A1(n_9550),
.A2(n_325),
.A3(n_323),
.B1(n_324),
.B2(n_326),
.Y(n_9673)
);

NAND2xp5_ASAP7_75t_L g9674 ( 
.A(n_9571),
.B(n_325),
.Y(n_9674)
);

OAI22xp5_ASAP7_75t_SL g9675 ( 
.A1(n_9253),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_9675)
);

AND2x4_ASAP7_75t_L g9676 ( 
.A(n_9176),
.B(n_9263),
.Y(n_9676)
);

INVx1_ASAP7_75t_L g9677 ( 
.A(n_9094),
.Y(n_9677)
);

INVx1_ASAP7_75t_L g9678 ( 
.A(n_9098),
.Y(n_9678)
);

NAND2xp5_ASAP7_75t_L g9679 ( 
.A(n_9369),
.B(n_326),
.Y(n_9679)
);

AOI22xp5_ASAP7_75t_L g9680 ( 
.A1(n_9178),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_9680)
);

OAI22xp5_ASAP7_75t_L g9681 ( 
.A1(n_9184),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_9681)
);

NAND2xp5_ASAP7_75t_L g9682 ( 
.A(n_9376),
.B(n_9156),
.Y(n_9682)
);

AND2x2_ASAP7_75t_L g9683 ( 
.A(n_9036),
.B(n_330),
.Y(n_9683)
);

BUFx8_ASAP7_75t_L g9684 ( 
.A(n_9051),
.Y(n_9684)
);

INVx2_ASAP7_75t_L g9685 ( 
.A(n_9054),
.Y(n_9685)
);

AOI22xp33_ASAP7_75t_L g9686 ( 
.A1(n_9434),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_9686)
);

NOR3xp33_ASAP7_75t_L g9687 ( 
.A(n_9304),
.B(n_331),
.C(n_332),
.Y(n_9687)
);

AOI21xp5_ASAP7_75t_L g9688 ( 
.A1(n_9498),
.A2(n_331),
.B(n_334),
.Y(n_9688)
);

OAI21xp5_ASAP7_75t_L g9689 ( 
.A1(n_9362),
.A2(n_334),
.B(n_335),
.Y(n_9689)
);

AOI21xp5_ASAP7_75t_L g9690 ( 
.A1(n_9505),
.A2(n_334),
.B(n_335),
.Y(n_9690)
);

AOI21xp5_ASAP7_75t_L g9691 ( 
.A1(n_9128),
.A2(n_335),
.B(n_336),
.Y(n_9691)
);

AOI22xp5_ASAP7_75t_L g9692 ( 
.A1(n_9208),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_9692)
);

OAI22xp5_ASAP7_75t_L g9693 ( 
.A1(n_9368),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_9693)
);

NAND2xp5_ASAP7_75t_L g9694 ( 
.A(n_9481),
.B(n_337),
.Y(n_9694)
);

NAND2xp33_ASAP7_75t_L g9695 ( 
.A(n_9445),
.B(n_338),
.Y(n_9695)
);

AND2x2_ASAP7_75t_L g9696 ( 
.A(n_9444),
.B(n_339),
.Y(n_9696)
);

AND2x2_ASAP7_75t_L g9697 ( 
.A(n_9444),
.B(n_339),
.Y(n_9697)
);

NOR2xp33_ASAP7_75t_L g9698 ( 
.A(n_9165),
.B(n_339),
.Y(n_9698)
);

NAND2xp5_ASAP7_75t_SL g9699 ( 
.A(n_9176),
.B(n_340),
.Y(n_9699)
);

OAI22xp5_ASAP7_75t_L g9700 ( 
.A1(n_9168),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_9700)
);

AOI21x1_ASAP7_75t_L g9701 ( 
.A1(n_9109),
.A2(n_340),
.B(n_341),
.Y(n_9701)
);

AOI21xp5_ASAP7_75t_L g9702 ( 
.A1(n_9534),
.A2(n_9570),
.B(n_9222),
.Y(n_9702)
);

NAND2xp5_ASAP7_75t_L g9703 ( 
.A(n_9491),
.B(n_341),
.Y(n_9703)
);

NAND2xp5_ASAP7_75t_L g9704 ( 
.A(n_9521),
.B(n_342),
.Y(n_9704)
);

BUFx6f_ASAP7_75t_L g9705 ( 
.A(n_9320),
.Y(n_9705)
);

NAND2xp5_ASAP7_75t_L g9706 ( 
.A(n_9579),
.B(n_343),
.Y(n_9706)
);

NAND2xp5_ASAP7_75t_SL g9707 ( 
.A(n_9263),
.B(n_9040),
.Y(n_9707)
);

OR2x6_ASAP7_75t_L g9708 ( 
.A(n_9131),
.B(n_9160),
.Y(n_9708)
);

NAND2xp5_ASAP7_75t_L g9709 ( 
.A(n_9027),
.B(n_343),
.Y(n_9709)
);

NAND2xp5_ASAP7_75t_SL g9710 ( 
.A(n_9058),
.B(n_343),
.Y(n_9710)
);

AOI21xp5_ASAP7_75t_L g9711 ( 
.A1(n_9570),
.A2(n_344),
.B(n_345),
.Y(n_9711)
);

NAND2xp5_ASAP7_75t_L g9712 ( 
.A(n_9034),
.B(n_344),
.Y(n_9712)
);

BUFx3_ASAP7_75t_L g9713 ( 
.A(n_9079),
.Y(n_9713)
);

INVx2_ASAP7_75t_L g9714 ( 
.A(n_9059),
.Y(n_9714)
);

NOR2xp33_ASAP7_75t_L g9715 ( 
.A(n_9286),
.B(n_345),
.Y(n_9715)
);

INVxp67_ASAP7_75t_L g9716 ( 
.A(n_9046),
.Y(n_9716)
);

INVx2_ASAP7_75t_L g9717 ( 
.A(n_9064),
.Y(n_9717)
);

AOI21xp5_ASAP7_75t_L g9718 ( 
.A1(n_9074),
.A2(n_346),
.B(n_347),
.Y(n_9718)
);

O2A1O1Ixp33_ASAP7_75t_L g9719 ( 
.A1(n_9457),
.A2(n_348),
.B(n_346),
.C(n_347),
.Y(n_9719)
);

NOR2xp33_ASAP7_75t_L g9720 ( 
.A(n_9112),
.B(n_348),
.Y(n_9720)
);

INVx1_ASAP7_75t_L g9721 ( 
.A(n_9117),
.Y(n_9721)
);

BUFx8_ASAP7_75t_L g9722 ( 
.A(n_9287),
.Y(n_9722)
);

AND2x2_ASAP7_75t_L g9723 ( 
.A(n_9538),
.B(n_348),
.Y(n_9723)
);

AOI21xp5_ASAP7_75t_L g9724 ( 
.A1(n_9077),
.A2(n_349),
.B(n_351),
.Y(n_9724)
);

AOI21xp5_ASAP7_75t_L g9725 ( 
.A1(n_9268),
.A2(n_349),
.B(n_351),
.Y(n_9725)
);

INVx2_ASAP7_75t_L g9726 ( 
.A(n_9071),
.Y(n_9726)
);

AOI21xp5_ASAP7_75t_L g9727 ( 
.A1(n_9038),
.A2(n_9069),
.B(n_9563),
.Y(n_9727)
);

INVx4_ASAP7_75t_L g9728 ( 
.A(n_9600),
.Y(n_9728)
);

AOI21xp5_ASAP7_75t_L g9729 ( 
.A1(n_9580),
.A2(n_349),
.B(n_351),
.Y(n_9729)
);

BUFx6f_ASAP7_75t_L g9730 ( 
.A(n_9320),
.Y(n_9730)
);

OAI21xp33_ASAP7_75t_L g9731 ( 
.A1(n_9345),
.A2(n_352),
.B(n_353),
.Y(n_9731)
);

CKINVDCx16_ASAP7_75t_R g9732 ( 
.A(n_9152),
.Y(n_9732)
);

OAI21xp5_ASAP7_75t_L g9733 ( 
.A1(n_9105),
.A2(n_352),
.B(n_353),
.Y(n_9733)
);

INVx2_ASAP7_75t_L g9734 ( 
.A(n_9083),
.Y(n_9734)
);

INVx1_ASAP7_75t_L g9735 ( 
.A(n_9118),
.Y(n_9735)
);

AOI21xp5_ASAP7_75t_L g9736 ( 
.A1(n_9479),
.A2(n_352),
.B(n_353),
.Y(n_9736)
);

AOI21x1_ASAP7_75t_L g9737 ( 
.A1(n_9235),
.A2(n_354),
.B(n_355),
.Y(n_9737)
);

NAND2xp5_ASAP7_75t_SL g9738 ( 
.A(n_9528),
.B(n_354),
.Y(n_9738)
);

NAND2xp5_ASAP7_75t_L g9739 ( 
.A(n_9530),
.B(n_354),
.Y(n_9739)
);

AOI21xp5_ASAP7_75t_L g9740 ( 
.A1(n_9090),
.A2(n_355),
.B(n_356),
.Y(n_9740)
);

INVx2_ASAP7_75t_L g9741 ( 
.A(n_9085),
.Y(n_9741)
);

INVx2_ASAP7_75t_L g9742 ( 
.A(n_9110),
.Y(n_9742)
);

AOI21xp5_ASAP7_75t_L g9743 ( 
.A1(n_9092),
.A2(n_355),
.B(n_356),
.Y(n_9743)
);

NAND2xp5_ASAP7_75t_SL g9744 ( 
.A(n_9578),
.B(n_356),
.Y(n_9744)
);

OAI22xp5_ASAP7_75t_L g9745 ( 
.A1(n_9198),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_9745)
);

INVx1_ASAP7_75t_L g9746 ( 
.A(n_9126),
.Y(n_9746)
);

INVx3_ASAP7_75t_L g9747 ( 
.A(n_9255),
.Y(n_9747)
);

NAND3xp33_ASAP7_75t_L g9748 ( 
.A(n_9431),
.B(n_357),
.C(n_358),
.Y(n_9748)
);

OAI22xp5_ASAP7_75t_L g9749 ( 
.A1(n_9330),
.A2(n_360),
.B1(n_357),
.B2(n_359),
.Y(n_9749)
);

NAND2xp5_ASAP7_75t_SL g9750 ( 
.A(n_9477),
.B(n_359),
.Y(n_9750)
);

OAI22xp5_ASAP7_75t_L g9751 ( 
.A1(n_9169),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_9751)
);

HB1xp67_ASAP7_75t_L g9752 ( 
.A(n_9448),
.Y(n_9752)
);

AOI22xp5_ASAP7_75t_L g9753 ( 
.A1(n_9134),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_9753)
);

INVx1_ASAP7_75t_L g9754 ( 
.A(n_9139),
.Y(n_9754)
);

OAI22xp5_ASAP7_75t_L g9755 ( 
.A1(n_9464),
.A2(n_364),
.B1(n_361),
.B2(n_363),
.Y(n_9755)
);

AOI21xp5_ASAP7_75t_L g9756 ( 
.A1(n_9104),
.A2(n_363),
.B(n_364),
.Y(n_9756)
);

AOI21xp5_ASAP7_75t_L g9757 ( 
.A1(n_9045),
.A2(n_365),
.B(n_366),
.Y(n_9757)
);

NAND2xp5_ASAP7_75t_L g9758 ( 
.A(n_9533),
.B(n_366),
.Y(n_9758)
);

NAND2xp5_ASAP7_75t_SL g9759 ( 
.A(n_9080),
.B(n_366),
.Y(n_9759)
);

NAND2xp5_ASAP7_75t_SL g9760 ( 
.A(n_9584),
.B(n_367),
.Y(n_9760)
);

INVx1_ASAP7_75t_L g9761 ( 
.A(n_9147),
.Y(n_9761)
);

NAND2xp5_ASAP7_75t_L g9762 ( 
.A(n_9541),
.B(n_367),
.Y(n_9762)
);

O2A1O1Ixp33_ASAP7_75t_L g9763 ( 
.A1(n_9462),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_9763)
);

AOI21xp5_ASAP7_75t_L g9764 ( 
.A1(n_9047),
.A2(n_368),
.B(n_369),
.Y(n_9764)
);

BUFx6f_ASAP7_75t_L g9765 ( 
.A(n_9055),
.Y(n_9765)
);

AOI21xp5_ASAP7_75t_L g9766 ( 
.A1(n_9050),
.A2(n_368),
.B(n_370),
.Y(n_9766)
);

NAND2xp5_ASAP7_75t_L g9767 ( 
.A(n_9543),
.B(n_370),
.Y(n_9767)
);

NAND2xp5_ASAP7_75t_L g9768 ( 
.A(n_9557),
.B(n_370),
.Y(n_9768)
);

AOI21xp5_ASAP7_75t_L g9769 ( 
.A1(n_9379),
.A2(n_9469),
.B(n_9548),
.Y(n_9769)
);

NAND2xp5_ASAP7_75t_L g9770 ( 
.A(n_9076),
.B(n_371),
.Y(n_9770)
);

NAND3xp33_ASAP7_75t_L g9771 ( 
.A(n_9116),
.B(n_371),
.C(n_372),
.Y(n_9771)
);

OAI21xp5_ASAP7_75t_L g9772 ( 
.A1(n_9441),
.A2(n_371),
.B(n_372),
.Y(n_9772)
);

AOI21xp5_ASAP7_75t_L g9773 ( 
.A1(n_9424),
.A2(n_9470),
.B(n_9248),
.Y(n_9773)
);

INVx1_ASAP7_75t_L g9774 ( 
.A(n_9150),
.Y(n_9774)
);

BUFx8_ASAP7_75t_L g9775 ( 
.A(n_9339),
.Y(n_9775)
);

NAND2xp5_ASAP7_75t_L g9776 ( 
.A(n_9524),
.B(n_373),
.Y(n_9776)
);

NAND2xp5_ASAP7_75t_L g9777 ( 
.A(n_9526),
.B(n_373),
.Y(n_9777)
);

OAI22xp5_ASAP7_75t_L g9778 ( 
.A1(n_9478),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_9778)
);

OAI22xp5_ASAP7_75t_L g9779 ( 
.A1(n_9392),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_9779)
);

BUFx6f_ASAP7_75t_L g9780 ( 
.A(n_9598),
.Y(n_9780)
);

INVx4_ASAP7_75t_L g9781 ( 
.A(n_9057),
.Y(n_9781)
);

OAI21xp5_ASAP7_75t_L g9782 ( 
.A1(n_9503),
.A2(n_374),
.B(n_377),
.Y(n_9782)
);

AO22x1_ASAP7_75t_L g9783 ( 
.A1(n_9364),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_9783)
);

NAND2xp5_ASAP7_75t_L g9784 ( 
.A(n_9536),
.B(n_378),
.Y(n_9784)
);

INVx2_ASAP7_75t_L g9785 ( 
.A(n_9115),
.Y(n_9785)
);

A2O1A1Ixp33_ASAP7_75t_L g9786 ( 
.A1(n_9391),
.A2(n_381),
.B(n_379),
.C(n_380),
.Y(n_9786)
);

CKINVDCx10_ASAP7_75t_R g9787 ( 
.A(n_9197),
.Y(n_9787)
);

NAND2xp5_ASAP7_75t_L g9788 ( 
.A(n_9540),
.B(n_9542),
.Y(n_9788)
);

NAND2xp5_ASAP7_75t_SL g9789 ( 
.A(n_9584),
.B(n_379),
.Y(n_9789)
);

AND2x6_ASAP7_75t_SL g9790 ( 
.A(n_9289),
.B(n_9336),
.Y(n_9790)
);

NOR2x1_ASAP7_75t_L g9791 ( 
.A(n_9393),
.B(n_380),
.Y(n_9791)
);

O2A1O1Ixp33_ASAP7_75t_L g9792 ( 
.A1(n_9157),
.A2(n_382),
.B(n_380),
.C(n_381),
.Y(n_9792)
);

INVx3_ASAP7_75t_L g9793 ( 
.A(n_9044),
.Y(n_9793)
);

NOR2xp33_ASAP7_75t_L g9794 ( 
.A(n_9241),
.B(n_382),
.Y(n_9794)
);

A2O1A1Ixp33_ASAP7_75t_L g9795 ( 
.A1(n_9323),
.A2(n_384),
.B(n_382),
.C(n_383),
.Y(n_9795)
);

AND2x6_ASAP7_75t_L g9796 ( 
.A(n_9052),
.B(n_9552),
.Y(n_9796)
);

AO32x1_ASAP7_75t_L g9797 ( 
.A1(n_9581),
.A2(n_385),
.A3(n_383),
.B1(n_384),
.B2(n_386),
.Y(n_9797)
);

OR2x6_ASAP7_75t_L g9798 ( 
.A(n_9111),
.B(n_383),
.Y(n_9798)
);

AOI21xp5_ASAP7_75t_L g9799 ( 
.A1(n_9511),
.A2(n_385),
.B(n_386),
.Y(n_9799)
);

AOI21xp5_ASAP7_75t_L g9800 ( 
.A1(n_9517),
.A2(n_386),
.B(n_387),
.Y(n_9800)
);

OAI22xp5_ASAP7_75t_SL g9801 ( 
.A1(n_9122),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_9801)
);

A2O1A1Ixp33_ASAP7_75t_L g9802 ( 
.A1(n_9078),
.A2(n_389),
.B(n_387),
.C(n_388),
.Y(n_9802)
);

NAND2xp5_ASAP7_75t_SL g9803 ( 
.A(n_9410),
.B(n_389),
.Y(n_9803)
);

NAND2xp5_ASAP7_75t_L g9804 ( 
.A(n_9553),
.B(n_390),
.Y(n_9804)
);

NAND2xp5_ASAP7_75t_L g9805 ( 
.A(n_9556),
.B(n_391),
.Y(n_9805)
);

AND2x2_ASAP7_75t_L g9806 ( 
.A(n_9244),
.B(n_391),
.Y(n_9806)
);

O2A1O1Ixp33_ASAP7_75t_L g9807 ( 
.A1(n_9599),
.A2(n_394),
.B(n_392),
.C(n_393),
.Y(n_9807)
);

BUFx6f_ASAP7_75t_L g9808 ( 
.A(n_9021),
.Y(n_9808)
);

OR2x2_ASAP7_75t_L g9809 ( 
.A(n_9227),
.B(n_392),
.Y(n_9809)
);

INVx1_ASAP7_75t_L g9810 ( 
.A(n_9163),
.Y(n_9810)
);

AOI21xp5_ASAP7_75t_L g9811 ( 
.A1(n_9523),
.A2(n_392),
.B(n_393),
.Y(n_9811)
);

AOI21xp5_ASAP7_75t_L g9812 ( 
.A1(n_9546),
.A2(n_393),
.B(n_394),
.Y(n_9812)
);

NAND2xp5_ASAP7_75t_L g9813 ( 
.A(n_9558),
.B(n_9562),
.Y(n_9813)
);

INVx11_ASAP7_75t_L g9814 ( 
.A(n_9067),
.Y(n_9814)
);

NAND2xp5_ASAP7_75t_L g9815 ( 
.A(n_9566),
.B(n_394),
.Y(n_9815)
);

A2O1A1Ixp33_ASAP7_75t_L g9816 ( 
.A1(n_9529),
.A2(n_397),
.B(n_395),
.C(n_396),
.Y(n_9816)
);

NAND2xp5_ASAP7_75t_L g9817 ( 
.A(n_9567),
.B(n_395),
.Y(n_9817)
);

NAND2xp5_ASAP7_75t_L g9818 ( 
.A(n_9568),
.B(n_396),
.Y(n_9818)
);

NAND2xp5_ASAP7_75t_L g9819 ( 
.A(n_9451),
.B(n_396),
.Y(n_9819)
);

AOI21xp5_ASAP7_75t_L g9820 ( 
.A1(n_9564),
.A2(n_397),
.B(n_398),
.Y(n_9820)
);

O2A1O1Ixp33_ASAP7_75t_SL g9821 ( 
.A1(n_9283),
.A2(n_399),
.B(n_397),
.C(n_398),
.Y(n_9821)
);

AOI21xp5_ASAP7_75t_L g9822 ( 
.A1(n_9229),
.A2(n_398),
.B(n_399),
.Y(n_9822)
);

NOR2xp33_ASAP7_75t_L g9823 ( 
.A(n_9367),
.B(n_399),
.Y(n_9823)
);

OAI22xp5_ASAP7_75t_L g9824 ( 
.A1(n_9240),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_9824)
);

A2O1A1Ixp33_ASAP7_75t_L g9825 ( 
.A1(n_9342),
.A2(n_9353),
.B(n_9583),
.C(n_9282),
.Y(n_9825)
);

NOR2xp33_ASAP7_75t_L g9826 ( 
.A(n_9191),
.B(n_400),
.Y(n_9826)
);

INVx1_ASAP7_75t_L g9827 ( 
.A(n_9166),
.Y(n_9827)
);

NOR2xp33_ASAP7_75t_L g9828 ( 
.A(n_9409),
.B(n_400),
.Y(n_9828)
);

AND2x2_ASAP7_75t_L g9829 ( 
.A(n_9267),
.B(n_401),
.Y(n_9829)
);

AOI21xp5_ASAP7_75t_L g9830 ( 
.A1(n_9492),
.A2(n_402),
.B(n_403),
.Y(n_9830)
);

AOI21xp5_ASAP7_75t_L g9831 ( 
.A1(n_9587),
.A2(n_402),
.B(n_403),
.Y(n_9831)
);

NAND2xp5_ASAP7_75t_L g9832 ( 
.A(n_9096),
.B(n_403),
.Y(n_9832)
);

NOR2xp33_ASAP7_75t_L g9833 ( 
.A(n_9405),
.B(n_9072),
.Y(n_9833)
);

NOR2xp33_ASAP7_75t_L g9834 ( 
.A(n_9343),
.B(n_404),
.Y(n_9834)
);

NAND2xp5_ASAP7_75t_L g9835 ( 
.A(n_9452),
.B(n_404),
.Y(n_9835)
);

NAND2xp5_ASAP7_75t_L g9836 ( 
.A(n_9453),
.B(n_404),
.Y(n_9836)
);

NAND2xp5_ASAP7_75t_L g9837 ( 
.A(n_9456),
.B(n_405),
.Y(n_9837)
);

INVx2_ASAP7_75t_L g9838 ( 
.A(n_9119),
.Y(n_9838)
);

INVxp67_ASAP7_75t_L g9839 ( 
.A(n_9032),
.Y(n_9839)
);

AOI21xp5_ASAP7_75t_L g9840 ( 
.A1(n_9588),
.A2(n_405),
.B(n_406),
.Y(n_9840)
);

INVx3_ASAP7_75t_L g9841 ( 
.A(n_9129),
.Y(n_9841)
);

AOI22xp5_ASAP7_75t_L g9842 ( 
.A1(n_9348),
.A2(n_9510),
.B1(n_9592),
.B2(n_9256),
.Y(n_9842)
);

AOI22x1_ASAP7_75t_L g9843 ( 
.A1(n_9474),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_9843)
);

AOI21xp5_ASAP7_75t_L g9844 ( 
.A1(n_9102),
.A2(n_406),
.B(n_407),
.Y(n_9844)
);

NAND2xp5_ASAP7_75t_L g9845 ( 
.A(n_9458),
.B(n_408),
.Y(n_9845)
);

NOR2x1_ASAP7_75t_L g9846 ( 
.A(n_9480),
.B(n_408),
.Y(n_9846)
);

INVx2_ASAP7_75t_L g9847 ( 
.A(n_9272),
.Y(n_9847)
);

INVx1_ASAP7_75t_L g9848 ( 
.A(n_9167),
.Y(n_9848)
);

AOI22xp5_ASAP7_75t_L g9849 ( 
.A1(n_9395),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_9849)
);

AOI21xp5_ASAP7_75t_L g9850 ( 
.A1(n_9460),
.A2(n_409),
.B(n_410),
.Y(n_9850)
);

AOI21xp5_ASAP7_75t_L g9851 ( 
.A1(n_9472),
.A2(n_409),
.B(n_410),
.Y(n_9851)
);

NOR2xp33_ASAP7_75t_L g9852 ( 
.A(n_9138),
.B(n_412),
.Y(n_9852)
);

AOI21xp5_ASAP7_75t_L g9853 ( 
.A1(n_9484),
.A2(n_412),
.B(n_413),
.Y(n_9853)
);

HB1xp67_ASAP7_75t_L g9854 ( 
.A(n_9185),
.Y(n_9854)
);

OAI21xp5_ASAP7_75t_L g9855 ( 
.A1(n_9209),
.A2(n_413),
.B(n_414),
.Y(n_9855)
);

NAND2xp5_ASAP7_75t_L g9856 ( 
.A(n_9486),
.B(n_9489),
.Y(n_9856)
);

AOI21xp5_ASAP7_75t_L g9857 ( 
.A1(n_9504),
.A2(n_413),
.B(n_414),
.Y(n_9857)
);

NAND2xp5_ASAP7_75t_SL g9858 ( 
.A(n_9410),
.B(n_9137),
.Y(n_9858)
);

NAND2xp5_ASAP7_75t_L g9859 ( 
.A(n_9514),
.B(n_415),
.Y(n_9859)
);

AOI21xp5_ASAP7_75t_L g9860 ( 
.A1(n_9520),
.A2(n_415),
.B(n_416),
.Y(n_9860)
);

AOI22x1_ASAP7_75t_L g9861 ( 
.A1(n_9440),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_9861)
);

NAND2xp5_ASAP7_75t_SL g9862 ( 
.A(n_9199),
.B(n_416),
.Y(n_9862)
);

BUFx12f_ASAP7_75t_L g9863 ( 
.A(n_9073),
.Y(n_9863)
);

INVx1_ASAP7_75t_L g9864 ( 
.A(n_9186),
.Y(n_9864)
);

NAND2xp5_ASAP7_75t_L g9865 ( 
.A(n_9467),
.B(n_417),
.Y(n_9865)
);

NAND2xp5_ASAP7_75t_L g9866 ( 
.A(n_9482),
.B(n_418),
.Y(n_9866)
);

INVx1_ASAP7_75t_L g9867 ( 
.A(n_9188),
.Y(n_9867)
);

INVx2_ASAP7_75t_L g9868 ( 
.A(n_9295),
.Y(n_9868)
);

INVx1_ASAP7_75t_L g9869 ( 
.A(n_9189),
.Y(n_9869)
);

INVx6_ASAP7_75t_L g9870 ( 
.A(n_9247),
.Y(n_9870)
);

NOR3xp33_ASAP7_75t_L g9871 ( 
.A(n_9333),
.B(n_418),
.C(n_419),
.Y(n_9871)
);

NAND2xp5_ASAP7_75t_L g9872 ( 
.A(n_9494),
.B(n_418),
.Y(n_9872)
);

AOI21xp5_ASAP7_75t_L g9873 ( 
.A1(n_9595),
.A2(n_420),
.B(n_421),
.Y(n_9873)
);

AOI21xp5_ASAP7_75t_L g9874 ( 
.A1(n_9041),
.A2(n_9509),
.B(n_9585),
.Y(n_9874)
);

NAND2xp5_ASAP7_75t_SL g9875 ( 
.A(n_9039),
.B(n_420),
.Y(n_9875)
);

AOI21xp5_ASAP7_75t_L g9876 ( 
.A1(n_9414),
.A2(n_420),
.B(n_421),
.Y(n_9876)
);

NAND2xp5_ASAP7_75t_L g9877 ( 
.A(n_9501),
.B(n_422),
.Y(n_9877)
);

INVx3_ASAP7_75t_L g9878 ( 
.A(n_9449),
.Y(n_9878)
);

AOI21xp5_ASAP7_75t_L g9879 ( 
.A1(n_9455),
.A2(n_422),
.B(n_423),
.Y(n_9879)
);

NOR2x1p5_ASAP7_75t_SL g9880 ( 
.A(n_9194),
.B(n_423),
.Y(n_9880)
);

OA22x2_ASAP7_75t_L g9881 ( 
.A1(n_9443),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_9881)
);

O2A1O1Ixp33_ASAP7_75t_SL g9882 ( 
.A1(n_9180),
.A2(n_427),
.B(n_424),
.C(n_426),
.Y(n_9882)
);

INVx2_ASAP7_75t_L g9883 ( 
.A(n_9303),
.Y(n_9883)
);

NOR2xp33_ASAP7_75t_L g9884 ( 
.A(n_9159),
.B(n_424),
.Y(n_9884)
);

OAI21xp5_ASAP7_75t_L g9885 ( 
.A1(n_9436),
.A2(n_426),
.B(n_427),
.Y(n_9885)
);

INVx2_ASAP7_75t_L g9886 ( 
.A(n_9314),
.Y(n_9886)
);

OAI21xp33_ASAP7_75t_L g9887 ( 
.A1(n_9572),
.A2(n_426),
.B(n_428),
.Y(n_9887)
);

AOI21xp5_ASAP7_75t_L g9888 ( 
.A1(n_9488),
.A2(n_429),
.B(n_430),
.Y(n_9888)
);

NAND2xp5_ASAP7_75t_L g9889 ( 
.A(n_9513),
.B(n_429),
.Y(n_9889)
);

INVx1_ASAP7_75t_L g9890 ( 
.A(n_9203),
.Y(n_9890)
);

NAND2xp5_ASAP7_75t_SL g9891 ( 
.A(n_9461),
.B(n_432),
.Y(n_9891)
);

AOI21x1_ASAP7_75t_L g9892 ( 
.A1(n_9179),
.A2(n_432),
.B(n_433),
.Y(n_9892)
);

OAI22xp5_ASAP7_75t_L g9893 ( 
.A1(n_9230),
.A2(n_9296),
.B1(n_9373),
.B2(n_9325),
.Y(n_9893)
);

CKINVDCx11_ASAP7_75t_R g9894 ( 
.A(n_9099),
.Y(n_9894)
);

O2A1O1Ixp33_ASAP7_75t_L g9895 ( 
.A1(n_9238),
.A2(n_434),
.B(n_432),
.C(n_433),
.Y(n_9895)
);

AOI21xp5_ASAP7_75t_L g9896 ( 
.A1(n_9575),
.A2(n_433),
.B(n_435),
.Y(n_9896)
);

NAND2xp5_ASAP7_75t_L g9897 ( 
.A(n_9519),
.B(n_435),
.Y(n_9897)
);

AOI22xp5_ASAP7_75t_L g9898 ( 
.A1(n_9218),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_9898)
);

AOI22xp5_ASAP7_75t_L g9899 ( 
.A1(n_9218),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.Y(n_9899)
);

NAND2xp5_ASAP7_75t_L g9900 ( 
.A(n_9026),
.B(n_9212),
.Y(n_9900)
);

AOI21xp5_ASAP7_75t_L g9901 ( 
.A1(n_9221),
.A2(n_437),
.B(n_438),
.Y(n_9901)
);

AOI21xp5_ASAP7_75t_L g9902 ( 
.A1(n_9082),
.A2(n_439),
.B(n_440),
.Y(n_9902)
);

AOI21xp5_ASAP7_75t_L g9903 ( 
.A1(n_9061),
.A2(n_439),
.B(n_441),
.Y(n_9903)
);

INVx1_ASAP7_75t_L g9904 ( 
.A(n_9228),
.Y(n_9904)
);

OAI21xp5_ASAP7_75t_L g9905 ( 
.A1(n_9447),
.A2(n_441),
.B(n_442),
.Y(n_9905)
);

NAND2xp5_ASAP7_75t_SL g9906 ( 
.A(n_9461),
.B(n_441),
.Y(n_9906)
);

OR2x6_ASAP7_75t_L g9907 ( 
.A(n_9473),
.B(n_442),
.Y(n_9907)
);

NAND2xp5_ASAP7_75t_L g9908 ( 
.A(n_9233),
.B(n_442),
.Y(n_9908)
);

INVx1_ASAP7_75t_L g9909 ( 
.A(n_9236),
.Y(n_9909)
);

AOI21x1_ASAP7_75t_L g9910 ( 
.A1(n_9319),
.A2(n_443),
.B(n_444),
.Y(n_9910)
);

NAND2xp5_ASAP7_75t_L g9911 ( 
.A(n_9242),
.B(n_443),
.Y(n_9911)
);

OAI21x1_ASAP7_75t_L g9912 ( 
.A1(n_9305),
.A2(n_444),
.B(n_445),
.Y(n_9912)
);

CKINVDCx5p33_ASAP7_75t_R g9913 ( 
.A(n_9020),
.Y(n_9913)
);

AOI22xp5_ASAP7_75t_L g9914 ( 
.A1(n_9218),
.A2(n_446),
.B1(n_444),
.B2(n_445),
.Y(n_9914)
);

NAND3xp33_ASAP7_75t_L g9915 ( 
.A(n_9254),
.B(n_446),
.C(n_447),
.Y(n_9915)
);

INVx1_ASAP7_75t_L g9916 ( 
.A(n_9243),
.Y(n_9916)
);

NAND2xp5_ASAP7_75t_SL g9917 ( 
.A(n_9497),
.B(n_446),
.Y(n_9917)
);

NAND2xp5_ASAP7_75t_L g9918 ( 
.A(n_9246),
.B(n_447),
.Y(n_9918)
);

CKINVDCx5p33_ASAP7_75t_R g9919 ( 
.A(n_9088),
.Y(n_9919)
);

INVxp67_ASAP7_75t_L g9920 ( 
.A(n_9043),
.Y(n_9920)
);

INVx2_ASAP7_75t_L g9921 ( 
.A(n_9340),
.Y(n_9921)
);

NAND2xp5_ASAP7_75t_SL g9922 ( 
.A(n_9465),
.B(n_447),
.Y(n_9922)
);

NAND2xp5_ASAP7_75t_L g9923 ( 
.A(n_9250),
.B(n_448),
.Y(n_9923)
);

NAND2xp5_ASAP7_75t_SL g9924 ( 
.A(n_9465),
.B(n_448),
.Y(n_9924)
);

NAND2xp5_ASAP7_75t_L g9925 ( 
.A(n_9258),
.B(n_448),
.Y(n_9925)
);

AOI21xp5_ASAP7_75t_L g9926 ( 
.A1(n_9097),
.A2(n_9113),
.B(n_9100),
.Y(n_9926)
);

AOI22xp5_ASAP7_75t_L g9927 ( 
.A1(n_9291),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.Y(n_9927)
);

BUFx6f_ASAP7_75t_L g9928 ( 
.A(n_9022),
.Y(n_9928)
);

BUFx2_ASAP7_75t_L g9929 ( 
.A(n_9060),
.Y(n_9929)
);

OAI21xp5_ASAP7_75t_L g9930 ( 
.A1(n_9375),
.A2(n_450),
.B(n_451),
.Y(n_9930)
);

NAND2xp5_ASAP7_75t_L g9931 ( 
.A(n_9260),
.B(n_450),
.Y(n_9931)
);

NAND2x1p5_ASAP7_75t_L g9932 ( 
.A(n_9132),
.B(n_451),
.Y(n_9932)
);

AOI21xp5_ASAP7_75t_L g9933 ( 
.A1(n_9383),
.A2(n_452),
.B(n_453),
.Y(n_9933)
);

NAND2xp5_ASAP7_75t_L g9934 ( 
.A(n_9262),
.B(n_452),
.Y(n_9934)
);

INVxp67_ASAP7_75t_L g9935 ( 
.A(n_9035),
.Y(n_9935)
);

AOI21x1_ASAP7_75t_L g9936 ( 
.A1(n_9371),
.A2(n_453),
.B(n_454),
.Y(n_9936)
);

INVx2_ASAP7_75t_L g9937 ( 
.A(n_9346),
.Y(n_9937)
);

INVx2_ASAP7_75t_L g9938 ( 
.A(n_9357),
.Y(n_9938)
);

OR2x6_ASAP7_75t_SL g9939 ( 
.A(n_9531),
.B(n_9151),
.Y(n_9939)
);

NOR2x1_ASAP7_75t_L g9940 ( 
.A(n_9499),
.B(n_453),
.Y(n_9940)
);

AOI21xp5_ASAP7_75t_L g9941 ( 
.A1(n_9312),
.A2(n_454),
.B(n_455),
.Y(n_9941)
);

AOI21xp5_ASAP7_75t_L g9942 ( 
.A1(n_9347),
.A2(n_454),
.B(n_455),
.Y(n_9942)
);

AND2x2_ASAP7_75t_L g9943 ( 
.A(n_9358),
.B(n_455),
.Y(n_9943)
);

NAND2xp5_ASAP7_75t_L g9944 ( 
.A(n_9265),
.B(n_456),
.Y(n_9944)
);

INVx2_ASAP7_75t_L g9945 ( 
.A(n_9377),
.Y(n_9945)
);

O2A1O1Ixp33_ASAP7_75t_L g9946 ( 
.A1(n_9280),
.A2(n_458),
.B(n_456),
.C(n_457),
.Y(n_9946)
);

INVx1_ASAP7_75t_SL g9947 ( 
.A(n_9285),
.Y(n_9947)
);

NAND2xp5_ASAP7_75t_L g9948 ( 
.A(n_9271),
.B(n_456),
.Y(n_9948)
);

INVx1_ASAP7_75t_L g9949 ( 
.A(n_9275),
.Y(n_9949)
);

O2A1O1Ixp5_ASAP7_75t_L g9950 ( 
.A1(n_9382),
.A2(n_459),
.B(n_457),
.C(n_458),
.Y(n_9950)
);

O2A1O1Ixp33_ASAP7_75t_L g9951 ( 
.A1(n_9352),
.A2(n_459),
.B(n_457),
.C(n_458),
.Y(n_9951)
);

AND2x2_ASAP7_75t_L g9952 ( 
.A(n_9386),
.B(n_459),
.Y(n_9952)
);

A2O1A1Ixp33_ASAP7_75t_L g9953 ( 
.A1(n_9415),
.A2(n_462),
.B(n_460),
.C(n_461),
.Y(n_9953)
);

NAND2xp5_ASAP7_75t_SL g9954 ( 
.A(n_9506),
.B(n_460),
.Y(n_9954)
);

NAND2xp5_ASAP7_75t_SL g9955 ( 
.A(n_9338),
.B(n_461),
.Y(n_9955)
);

AOI21xp5_ASAP7_75t_L g9956 ( 
.A1(n_9360),
.A2(n_9399),
.B(n_9378),
.Y(n_9956)
);

NAND2xp5_ASAP7_75t_L g9957 ( 
.A(n_9279),
.B(n_461),
.Y(n_9957)
);

CKINVDCx10_ASAP7_75t_R g9958 ( 
.A(n_9197),
.Y(n_9958)
);

AOI21xp5_ASAP7_75t_L g9959 ( 
.A1(n_9555),
.A2(n_462),
.B(n_463),
.Y(n_9959)
);

INVx2_ASAP7_75t_L g9960 ( 
.A(n_9084),
.Y(n_9960)
);

NAND2xp5_ASAP7_75t_SL g9961 ( 
.A(n_9338),
.B(n_462),
.Y(n_9961)
);

INVx2_ASAP7_75t_L g9962 ( 
.A(n_9329),
.Y(n_9962)
);

NAND2xp5_ASAP7_75t_L g9963 ( 
.A(n_9281),
.B(n_463),
.Y(n_9963)
);

INVx1_ASAP7_75t_L g9964 ( 
.A(n_9288),
.Y(n_9964)
);

O2A1O1Ixp33_ASAP7_75t_L g9965 ( 
.A1(n_9225),
.A2(n_466),
.B(n_464),
.C(n_465),
.Y(n_9965)
);

NAND2xp5_ASAP7_75t_L g9966 ( 
.A(n_9290),
.B(n_464),
.Y(n_9966)
);

AOI21xp5_ASAP7_75t_L g9967 ( 
.A1(n_9187),
.A2(n_465),
.B(n_466),
.Y(n_9967)
);

BUFx2_ASAP7_75t_L g9968 ( 
.A(n_9200),
.Y(n_9968)
);

AOI21xp5_ASAP7_75t_L g9969 ( 
.A1(n_9193),
.A2(n_466),
.B(n_467),
.Y(n_9969)
);

A2O1A1Ixp33_ASAP7_75t_L g9970 ( 
.A1(n_9374),
.A2(n_469),
.B(n_467),
.C(n_468),
.Y(n_9970)
);

INVx1_ASAP7_75t_L g9971 ( 
.A(n_9297),
.Y(n_9971)
);

NAND2x1p5_ASAP7_75t_L g9972 ( 
.A(n_9075),
.B(n_468),
.Y(n_9972)
);

OAI22xp5_ASAP7_75t_L g9973 ( 
.A1(n_9332),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_9973)
);

INVx1_ASAP7_75t_L g9974 ( 
.A(n_9299),
.Y(n_9974)
);

OAI22xp5_ASAP7_75t_L g9975 ( 
.A1(n_9205),
.A2(n_9426),
.B1(n_9214),
.B2(n_9582),
.Y(n_9975)
);

AO21x1_ASAP7_75t_L g9976 ( 
.A1(n_9576),
.A2(n_469),
.B(n_470),
.Y(n_9976)
);

AOI21xp5_ASAP7_75t_L g9977 ( 
.A1(n_9195),
.A2(n_470),
.B(n_471),
.Y(n_9977)
);

OAI22xp5_ASAP7_75t_L g9978 ( 
.A1(n_9476),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_9978)
);

OAI22xp5_ASAP7_75t_L g9979 ( 
.A1(n_9476),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_9979)
);

O2A1O1Ixp33_ASAP7_75t_L g9980 ( 
.A1(n_9401),
.A2(n_475),
.B(n_473),
.C(n_474),
.Y(n_9980)
);

NAND2xp5_ASAP7_75t_L g9981 ( 
.A(n_9301),
.B(n_474),
.Y(n_9981)
);

AOI21xp5_ASAP7_75t_L g9982 ( 
.A1(n_9196),
.A2(n_474),
.B(n_476),
.Y(n_9982)
);

AOI21xp5_ASAP7_75t_L g9983 ( 
.A1(n_9217),
.A2(n_476),
.B(n_477),
.Y(n_9983)
);

OAI22xp5_ASAP7_75t_L g9984 ( 
.A1(n_9537),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_9984)
);

NAND2xp5_ASAP7_75t_L g9985 ( 
.A(n_9311),
.B(n_477),
.Y(n_9985)
);

NAND2xp5_ASAP7_75t_SL g9986 ( 
.A(n_9018),
.B(n_9459),
.Y(n_9986)
);

NOR2xp33_ASAP7_75t_L g9987 ( 
.A(n_9403),
.B(n_478),
.Y(n_9987)
);

AND2x4_ASAP7_75t_L g9988 ( 
.A(n_9023),
.B(n_9056),
.Y(n_9988)
);

AOI21xp5_ASAP7_75t_L g9989 ( 
.A1(n_9220),
.A2(n_479),
.B(n_480),
.Y(n_9989)
);

NAND2xp5_ASAP7_75t_L g9990 ( 
.A(n_9315),
.B(n_479),
.Y(n_9990)
);

NAND2xp5_ASAP7_75t_L g9991 ( 
.A(n_9316),
.B(n_480),
.Y(n_9991)
);

O2A1O1Ixp33_ASAP7_75t_L g9992 ( 
.A1(n_9145),
.A2(n_483),
.B(n_481),
.C(n_482),
.Y(n_9992)
);

INVx2_ASAP7_75t_L g9993 ( 
.A(n_9334),
.Y(n_9993)
);

AOI22xp5_ASAP7_75t_L g9994 ( 
.A1(n_9291),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_9994)
);

NAND2xp5_ASAP7_75t_L g9995 ( 
.A(n_9317),
.B(n_482),
.Y(n_9995)
);

NAND2xp5_ASAP7_75t_L g9996 ( 
.A(n_9318),
.B(n_483),
.Y(n_9996)
);

AOI22xp5_ASAP7_75t_L g9997 ( 
.A1(n_9291),
.A2(n_486),
.B1(n_484),
.B2(n_485),
.Y(n_9997)
);

O2A1O1Ixp33_ASAP7_75t_L g9998 ( 
.A1(n_9161),
.A2(n_487),
.B(n_484),
.C(n_485),
.Y(n_9998)
);

AOI22xp33_ASAP7_75t_L g9999 ( 
.A1(n_9591),
.A2(n_488),
.B1(n_485),
.B2(n_487),
.Y(n_9999)
);

OA22x2_ASAP7_75t_L g10000 ( 
.A1(n_9496),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_10000)
);

OAI22xp5_ASAP7_75t_SL g10001 ( 
.A1(n_9361),
.A2(n_9403),
.B1(n_9313),
.B2(n_9321),
.Y(n_10001)
);

INVx11_ASAP7_75t_L g10002 ( 
.A(n_9364),
.Y(n_10002)
);

AOI21xp5_ASAP7_75t_L g10003 ( 
.A1(n_9223),
.A2(n_488),
.B(n_489),
.Y(n_10003)
);

BUFx12f_ASAP7_75t_L g10004 ( 
.A(n_9106),
.Y(n_10004)
);

NAND2xp5_ASAP7_75t_L g10005 ( 
.A(n_9322),
.B(n_489),
.Y(n_10005)
);

A2O1A1Ixp33_ASAP7_75t_L g10006 ( 
.A1(n_9430),
.A2(n_492),
.B(n_490),
.C(n_491),
.Y(n_10006)
);

INVx2_ASAP7_75t_L g10007 ( 
.A(n_9337),
.Y(n_10007)
);

OAI321xp33_ASAP7_75t_L g10008 ( 
.A1(n_9142),
.A2(n_492),
.A3(n_494),
.B1(n_490),
.B2(n_491),
.C(n_493),
.Y(n_10008)
);

INVx1_ASAP7_75t_L g10009 ( 
.A(n_9327),
.Y(n_10009)
);

NOR2xp33_ASAP7_75t_SL g10010 ( 
.A(n_9361),
.B(n_493),
.Y(n_10010)
);

AOI22xp5_ASAP7_75t_L g10011 ( 
.A1(n_9364),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_10011)
);

AOI22x1_ASAP7_75t_L g10012 ( 
.A1(n_9239),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.Y(n_10012)
);

NOR2xp33_ASAP7_75t_L g10013 ( 
.A(n_9309),
.B(n_496),
.Y(n_10013)
);

OAI21xp33_ASAP7_75t_L g10014 ( 
.A1(n_9396),
.A2(n_496),
.B(n_497),
.Y(n_10014)
);

NAND2xp5_ASAP7_75t_L g10015 ( 
.A(n_9370),
.B(n_498),
.Y(n_10015)
);

AND2x4_ASAP7_75t_L g10016 ( 
.A(n_9388),
.B(n_498),
.Y(n_10016)
);

INVx2_ASAP7_75t_L g10017 ( 
.A(n_9344),
.Y(n_10017)
);

INVx1_ASAP7_75t_L g10018 ( 
.A(n_9394),
.Y(n_10018)
);

AOI21xp5_ASAP7_75t_L g10019 ( 
.A1(n_9234),
.A2(n_499),
.B(n_500),
.Y(n_10019)
);

AOI21xp5_ASAP7_75t_L g10020 ( 
.A1(n_9264),
.A2(n_499),
.B(n_500),
.Y(n_10020)
);

NOR2x1_ASAP7_75t_L g10021 ( 
.A(n_9446),
.B(n_500),
.Y(n_10021)
);

AO21x1_ASAP7_75t_L g10022 ( 
.A1(n_9133),
.A2(n_501),
.B(n_502),
.Y(n_10022)
);

AOI21xp5_ASAP7_75t_L g10023 ( 
.A1(n_9270),
.A2(n_501),
.B(n_502),
.Y(n_10023)
);

NAND2xp5_ASAP7_75t_SL g10024 ( 
.A(n_9586),
.B(n_9326),
.Y(n_10024)
);

O2A1O1Ixp33_ASAP7_75t_L g10025 ( 
.A1(n_9162),
.A2(n_503),
.B(n_501),
.C(n_502),
.Y(n_10025)
);

AOI21xp5_ASAP7_75t_L g10026 ( 
.A1(n_9292),
.A2(n_503),
.B(n_504),
.Y(n_10026)
);

NOR2xp33_ASAP7_75t_L g10027 ( 
.A(n_9266),
.B(n_503),
.Y(n_10027)
);

INVx2_ASAP7_75t_L g10028 ( 
.A(n_9349),
.Y(n_10028)
);

BUFx6f_ASAP7_75t_L g10029 ( 
.A(n_9121),
.Y(n_10029)
);

NOR2xp33_ASAP7_75t_L g10030 ( 
.A(n_9466),
.B(n_504),
.Y(n_10030)
);

NOR2xp33_ASAP7_75t_L g10031 ( 
.A(n_9328),
.B(n_505),
.Y(n_10031)
);

BUFx3_ASAP7_75t_L g10032 ( 
.A(n_9276),
.Y(n_10032)
);

INVx2_ASAP7_75t_SL g10033 ( 
.A(n_9277),
.Y(n_10033)
);

BUFx6f_ASAP7_75t_L g10034 ( 
.A(n_9406),
.Y(n_10034)
);

INVx2_ASAP7_75t_L g10035 ( 
.A(n_9354),
.Y(n_10035)
);

AOI22xp33_ASAP7_75t_L g10036 ( 
.A1(n_9432),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_10036)
);

INVx1_ASAP7_75t_L g10037 ( 
.A(n_9398),
.Y(n_10037)
);

AND2x2_ASAP7_75t_L g10038 ( 
.A(n_9417),
.B(n_505),
.Y(n_10038)
);

INVx2_ASAP7_75t_L g10039 ( 
.A(n_9363),
.Y(n_10039)
);

NAND2xp5_ASAP7_75t_L g10040 ( 
.A(n_9140),
.B(n_506),
.Y(n_10040)
);

NAND2xp5_ASAP7_75t_L g10041 ( 
.A(n_9063),
.B(n_506),
.Y(n_10041)
);

INVx2_ASAP7_75t_L g10042 ( 
.A(n_9365),
.Y(n_10042)
);

NAND3xp33_ASAP7_75t_L g10043 ( 
.A(n_9381),
.B(n_507),
.C(n_508),
.Y(n_10043)
);

NAND2xp5_ASAP7_75t_L g10044 ( 
.A(n_9091),
.B(n_509),
.Y(n_10044)
);

NOR2xp33_ASAP7_75t_L g10045 ( 
.A(n_9103),
.B(n_509),
.Y(n_10045)
);

NAND2xp5_ASAP7_75t_L g10046 ( 
.A(n_9207),
.B(n_509),
.Y(n_10046)
);

NAND2xp5_ASAP7_75t_L g10047 ( 
.A(n_9384),
.B(n_9306),
.Y(n_10047)
);

NAND2xp33_ASAP7_75t_SL g10048 ( 
.A(n_9042),
.B(n_510),
.Y(n_10048)
);

A2O1A1Ixp33_ASAP7_75t_L g10049 ( 
.A1(n_9144),
.A2(n_513),
.B(n_511),
.C(n_512),
.Y(n_10049)
);

AOI21xp5_ASAP7_75t_L g10050 ( 
.A1(n_9593),
.A2(n_511),
.B(n_514),
.Y(n_10050)
);

AOI22xp5_ASAP7_75t_L g10051 ( 
.A1(n_9493),
.A2(n_515),
.B1(n_511),
.B2(n_514),
.Y(n_10051)
);

AOI21xp5_ASAP7_75t_L g10052 ( 
.A1(n_9485),
.A2(n_515),
.B(n_516),
.Y(n_10052)
);

NAND2xp5_ASAP7_75t_L g10053 ( 
.A(n_9307),
.B(n_516),
.Y(n_10053)
);

OA22x2_ASAP7_75t_L g10054 ( 
.A1(n_9525),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_10054)
);

AND2x2_ASAP7_75t_L g10055 ( 
.A(n_9463),
.B(n_518),
.Y(n_10055)
);

NAND2xp5_ASAP7_75t_SL g10056 ( 
.A(n_9535),
.B(n_519),
.Y(n_10056)
);

AOI21xp5_ASAP7_75t_L g10057 ( 
.A1(n_9490),
.A2(n_519),
.B(n_520),
.Y(n_10057)
);

INVx1_ASAP7_75t_L g10058 ( 
.A(n_9413),
.Y(n_10058)
);

OAI21x1_ASAP7_75t_L g10059 ( 
.A1(n_9418),
.A2(n_520),
.B(n_521),
.Y(n_10059)
);

O2A1O1Ixp33_ASAP7_75t_L g10060 ( 
.A1(n_9500),
.A2(n_9495),
.B(n_9508),
.C(n_9502),
.Y(n_10060)
);

INVx2_ASAP7_75t_SL g10061 ( 
.A(n_9294),
.Y(n_10061)
);

AOI21xp5_ASAP7_75t_L g10062 ( 
.A1(n_9515),
.A2(n_521),
.B(n_522),
.Y(n_10062)
);

AOI21xp5_ASAP7_75t_L g10063 ( 
.A1(n_9516),
.A2(n_521),
.B(n_522),
.Y(n_10063)
);

O2A1O1Ixp5_ASAP7_75t_L g10064 ( 
.A1(n_9177),
.A2(n_524),
.B(n_522),
.C(n_523),
.Y(n_10064)
);

NAND2xp5_ASAP7_75t_SL g10065 ( 
.A(n_9539),
.B(n_523),
.Y(n_10065)
);

INVx1_ASAP7_75t_L g10066 ( 
.A(n_9422),
.Y(n_10066)
);

AOI21xp5_ASAP7_75t_L g10067 ( 
.A1(n_9522),
.A2(n_523),
.B(n_524),
.Y(n_10067)
);

AND2x2_ASAP7_75t_L g10068 ( 
.A(n_9249),
.B(n_9518),
.Y(n_10068)
);

AOI21xp5_ASAP7_75t_L g10069 ( 
.A1(n_9527),
.A2(n_524),
.B(n_525),
.Y(n_10069)
);

O2A1O1Ixp33_ASAP7_75t_L g10070 ( 
.A1(n_9545),
.A2(n_527),
.B(n_525),
.C(n_526),
.Y(n_10070)
);

INVx2_ASAP7_75t_L g10071 ( 
.A(n_9124),
.Y(n_10071)
);

INVx4_ASAP7_75t_L g10072 ( 
.A(n_9335),
.Y(n_10072)
);

AO32x1_ASAP7_75t_L g10073 ( 
.A1(n_9350),
.A2(n_527),
.A3(n_525),
.B1(n_526),
.B2(n_528),
.Y(n_10073)
);

AOI21xp5_ASAP7_75t_L g10074 ( 
.A1(n_9551),
.A2(n_527),
.B(n_529),
.Y(n_10074)
);

INVx2_ASAP7_75t_L g10075 ( 
.A(n_9135),
.Y(n_10075)
);

INVx2_ASAP7_75t_L g10076 ( 
.A(n_9146),
.Y(n_10076)
);

AOI21xp5_ASAP7_75t_L g10077 ( 
.A1(n_9554),
.A2(n_529),
.B(n_530),
.Y(n_10077)
);

INVx1_ASAP7_75t_L g10078 ( 
.A(n_9427),
.Y(n_10078)
);

INVx2_ASAP7_75t_L g10079 ( 
.A(n_9148),
.Y(n_10079)
);

HB1xp67_ASAP7_75t_L g10080 ( 
.A(n_9589),
.Y(n_10080)
);

INVx2_ASAP7_75t_L g10081 ( 
.A(n_9155),
.Y(n_10081)
);

INVx2_ASAP7_75t_L g10082 ( 
.A(n_9170),
.Y(n_10082)
);

INVx2_ASAP7_75t_L g10083 ( 
.A(n_9173),
.Y(n_10083)
);

NAND2xp5_ASAP7_75t_L g10084 ( 
.A(n_9308),
.B(n_529),
.Y(n_10084)
);

AOI22xp5_ASAP7_75t_L g10085 ( 
.A1(n_9331),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.Y(n_10085)
);

NAND2xp5_ASAP7_75t_L g10086 ( 
.A(n_9086),
.B(n_531),
.Y(n_10086)
);

NOR2xp33_ASAP7_75t_L g10087 ( 
.A(n_9211),
.B(n_531),
.Y(n_10087)
);

AOI22xp33_ASAP7_75t_L g10088 ( 
.A1(n_9421),
.A2(n_534),
.B1(n_532),
.B2(n_533),
.Y(n_10088)
);

INVx2_ASAP7_75t_SL g10089 ( 
.A(n_9231),
.Y(n_10089)
);

AOI21xp5_ASAP7_75t_L g10090 ( 
.A1(n_9565),
.A2(n_533),
.B(n_534),
.Y(n_10090)
);

INVx1_ASAP7_75t_L g10091 ( 
.A(n_9442),
.Y(n_10091)
);

BUFx8_ASAP7_75t_L g10092 ( 
.A(n_9219),
.Y(n_10092)
);

NOR2xp33_ASAP7_75t_L g10093 ( 
.A(n_9210),
.B(n_533),
.Y(n_10093)
);

AOI21xp5_ASAP7_75t_L g10094 ( 
.A1(n_9574),
.A2(n_534),
.B(n_535),
.Y(n_10094)
);

INVx2_ASAP7_75t_L g10095 ( 
.A(n_9181),
.Y(n_10095)
);

OAI21x1_ASAP7_75t_L g10096 ( 
.A1(n_9183),
.A2(n_535),
.B(n_536),
.Y(n_10096)
);

AOI21xp5_ASAP7_75t_L g10097 ( 
.A1(n_9549),
.A2(n_9573),
.B(n_9341),
.Y(n_10097)
);

BUFx2_ASAP7_75t_L g10098 ( 
.A(n_9428),
.Y(n_10098)
);

INVx5_ASAP7_75t_L g10099 ( 
.A(n_9507),
.Y(n_10099)
);

AOI21xp5_ASAP7_75t_L g10100 ( 
.A1(n_9416),
.A2(n_535),
.B(n_536),
.Y(n_10100)
);

BUFx6f_ASAP7_75t_L g10101 ( 
.A(n_9407),
.Y(n_10101)
);

NAND2xp5_ASAP7_75t_SL g10102 ( 
.A(n_9512),
.B(n_536),
.Y(n_10102)
);

BUFx12f_ASAP7_75t_L g10103 ( 
.A(n_9154),
.Y(n_10103)
);

AOI21xp5_ASAP7_75t_L g10104 ( 
.A1(n_9366),
.A2(n_537),
.B(n_538),
.Y(n_10104)
);

NAND2xp5_ASAP7_75t_L g10105 ( 
.A(n_9298),
.B(n_537),
.Y(n_10105)
);

AND2x2_ASAP7_75t_L g10106 ( 
.A(n_9274),
.B(n_537),
.Y(n_10106)
);

INVx2_ASAP7_75t_L g10107 ( 
.A(n_9192),
.Y(n_10107)
);

INVxp67_ASAP7_75t_SL g10108 ( 
.A(n_9420),
.Y(n_10108)
);

INVx3_ASAP7_75t_L g10109 ( 
.A(n_9216),
.Y(n_10109)
);

AOI21xp5_ASAP7_75t_L g10110 ( 
.A1(n_9224),
.A2(n_538),
.B(n_539),
.Y(n_10110)
);

OAI21xp33_ASAP7_75t_L g10111 ( 
.A1(n_9577),
.A2(n_538),
.B(n_539),
.Y(n_10111)
);

OAI22xp5_ASAP7_75t_L g10112 ( 
.A1(n_9324),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_10112)
);

AOI21xp5_ASAP7_75t_L g10113 ( 
.A1(n_9171),
.A2(n_540),
.B(n_541),
.Y(n_10113)
);

NAND2xp5_ASAP7_75t_L g10114 ( 
.A(n_9201),
.B(n_542),
.Y(n_10114)
);

OAI21xp5_ASAP7_75t_L g10115 ( 
.A1(n_9544),
.A2(n_543),
.B(n_544),
.Y(n_10115)
);

AOI21xp5_ASAP7_75t_L g10116 ( 
.A1(n_9439),
.A2(n_543),
.B(n_545),
.Y(n_10116)
);

NAND2xp5_ASAP7_75t_L g10117 ( 
.A(n_9206),
.B(n_543),
.Y(n_10117)
);

BUFx2_ASAP7_75t_L g10118 ( 
.A(n_9237),
.Y(n_10118)
);

AOI22xp5_ASAP7_75t_L g10119 ( 
.A1(n_9547),
.A2(n_9182),
.B1(n_9355),
.B2(n_9559),
.Y(n_10119)
);

NOR2x1_ASAP7_75t_L g10120 ( 
.A(n_9158),
.B(n_9475),
.Y(n_10120)
);

AOI21xp5_ASAP7_75t_L g10121 ( 
.A1(n_9081),
.A2(n_545),
.B(n_546),
.Y(n_10121)
);

NAND2xp5_ASAP7_75t_L g10122 ( 
.A(n_9232),
.B(n_545),
.Y(n_10122)
);

AOI21xp5_ASAP7_75t_L g10123 ( 
.A1(n_9569),
.A2(n_546),
.B(n_547),
.Y(n_10123)
);

AOI21xp5_ASAP7_75t_L g10124 ( 
.A1(n_9561),
.A2(n_546),
.B(n_547),
.Y(n_10124)
);

NAND2xp5_ASAP7_75t_SL g10125 ( 
.A(n_9359),
.B(n_548),
.Y(n_10125)
);

AOI21xp5_ASAP7_75t_L g10126 ( 
.A1(n_9560),
.A2(n_548),
.B(n_549),
.Y(n_10126)
);

NAND2xp5_ASAP7_75t_L g10127 ( 
.A(n_9245),
.B(n_9251),
.Y(n_10127)
);

NAND2xp5_ASAP7_75t_L g10128 ( 
.A(n_9252),
.B(n_548),
.Y(n_10128)
);

AOI21xp5_ASAP7_75t_L g10129 ( 
.A1(n_9257),
.A2(n_549),
.B(n_550),
.Y(n_10129)
);

AOI21xp5_ASAP7_75t_L g10130 ( 
.A1(n_9259),
.A2(n_550),
.B(n_551),
.Y(n_10130)
);

NOR2xp33_ASAP7_75t_R g10131 ( 
.A(n_9404),
.B(n_550),
.Y(n_10131)
);

NAND2xp5_ASAP7_75t_L g10132 ( 
.A(n_9269),
.B(n_551),
.Y(n_10132)
);

INVx1_ASAP7_75t_L g10133 ( 
.A(n_9390),
.Y(n_10133)
);

AO22x1_ASAP7_75t_L g10134 ( 
.A1(n_9532),
.A2(n_9273),
.B1(n_9471),
.B2(n_9402),
.Y(n_10134)
);

INVx1_ASAP7_75t_L g10135 ( 
.A(n_9397),
.Y(n_10135)
);

NAND2xp5_ASAP7_75t_SL g10136 ( 
.A(n_9351),
.B(n_552),
.Y(n_10136)
);

AND2x2_ASAP7_75t_L g10137 ( 
.A(n_9261),
.B(n_552),
.Y(n_10137)
);

AO32x1_ASAP7_75t_L g10138 ( 
.A1(n_9408),
.A2(n_555),
.A3(n_553),
.B1(n_554),
.B2(n_556),
.Y(n_10138)
);

NOR2x1_ASAP7_75t_R g10139 ( 
.A(n_9411),
.B(n_553),
.Y(n_10139)
);

INVx1_ASAP7_75t_L g10140 ( 
.A(n_9412),
.Y(n_10140)
);

INVx3_ASAP7_75t_L g10141 ( 
.A(n_9419),
.Y(n_10141)
);

OAI21xp5_ASAP7_75t_L g10142 ( 
.A1(n_9310),
.A2(n_553),
.B(n_554),
.Y(n_10142)
);

NAND2xp5_ASAP7_75t_SL g10143 ( 
.A(n_9425),
.B(n_554),
.Y(n_10143)
);

NOR2xp33_ASAP7_75t_L g10144 ( 
.A(n_9487),
.B(n_555),
.Y(n_10144)
);

AOI21xp5_ASAP7_75t_L g10145 ( 
.A1(n_9429),
.A2(n_556),
.B(n_557),
.Y(n_10145)
);

AOI21xp5_ASAP7_75t_L g10146 ( 
.A1(n_9435),
.A2(n_556),
.B(n_557),
.Y(n_10146)
);

OA22x2_ASAP7_75t_L g10147 ( 
.A1(n_9437),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_10147)
);

AND2x2_ASAP7_75t_L g10148 ( 
.A(n_9438),
.B(n_558),
.Y(n_10148)
);

OAI21xp5_ASAP7_75t_L g10149 ( 
.A1(n_9107),
.A2(n_559),
.B(n_560),
.Y(n_10149)
);

A2O1A1Ixp33_ASAP7_75t_L g10150 ( 
.A1(n_9107),
.A2(n_561),
.B(n_559),
.C(n_560),
.Y(n_10150)
);

NAND2xp5_ASAP7_75t_L g10151 ( 
.A(n_9671),
.B(n_561),
.Y(n_10151)
);

AOI21xp5_ASAP7_75t_L g10152 ( 
.A1(n_9607),
.A2(n_562),
.B(n_563),
.Y(n_10152)
);

AOI21xp33_ASAP7_75t_L g10153 ( 
.A1(n_9624),
.A2(n_562),
.B(n_563),
.Y(n_10153)
);

NAND2xp5_ASAP7_75t_L g10154 ( 
.A(n_9716),
.B(n_564),
.Y(n_10154)
);

BUFx2_ASAP7_75t_R g10155 ( 
.A(n_9657),
.Y(n_10155)
);

INVx2_ASAP7_75t_L g10156 ( 
.A(n_9960),
.Y(n_10156)
);

INVxp67_ASAP7_75t_SL g10157 ( 
.A(n_9605),
.Y(n_10157)
);

INVx3_ASAP7_75t_L g10158 ( 
.A(n_9808),
.Y(n_10158)
);

AO21x2_ASAP7_75t_L g10159 ( 
.A1(n_9707),
.A2(n_564),
.B(n_565),
.Y(n_10159)
);

AOI21xp5_ASAP7_75t_L g10160 ( 
.A1(n_9647),
.A2(n_564),
.B(n_565),
.Y(n_10160)
);

NAND2xp5_ASAP7_75t_L g10161 ( 
.A(n_9662),
.B(n_565),
.Y(n_10161)
);

INVx2_ASAP7_75t_SL g10162 ( 
.A(n_9775),
.Y(n_10162)
);

NAND2xp5_ASAP7_75t_L g10163 ( 
.A(n_9920),
.B(n_566),
.Y(n_10163)
);

AOI22xp5_ASAP7_75t_L g10164 ( 
.A1(n_9842),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_10164)
);

OAI21x1_ASAP7_75t_SL g10165 ( 
.A1(n_9620),
.A2(n_566),
.B(n_567),
.Y(n_10165)
);

NAND2xp5_ASAP7_75t_L g10166 ( 
.A(n_9935),
.B(n_567),
.Y(n_10166)
);

NAND2xp5_ASAP7_75t_L g10167 ( 
.A(n_9854),
.B(n_568),
.Y(n_10167)
);

INVxp67_ASAP7_75t_SL g10168 ( 
.A(n_9645),
.Y(n_10168)
);

HB1xp67_ASAP7_75t_L g10169 ( 
.A(n_9752),
.Y(n_10169)
);

AOI211x1_ASAP7_75t_L g10170 ( 
.A1(n_10134),
.A2(n_570),
.B(n_568),
.C(n_569),
.Y(n_10170)
);

NAND2xp5_ASAP7_75t_L g10171 ( 
.A(n_9619),
.B(n_569),
.Y(n_10171)
);

INVx2_ASAP7_75t_L g10172 ( 
.A(n_9962),
.Y(n_10172)
);

O2A1O1Ixp5_ASAP7_75t_L g10173 ( 
.A1(n_9783),
.A2(n_571),
.B(n_569),
.C(n_570),
.Y(n_10173)
);

INVx1_ASAP7_75t_L g10174 ( 
.A(n_9630),
.Y(n_10174)
);

NAND2x1p5_ASAP7_75t_L g10175 ( 
.A(n_9676),
.B(n_571),
.Y(n_10175)
);

NAND2xp5_ASAP7_75t_L g10176 ( 
.A(n_9839),
.B(n_571),
.Y(n_10176)
);

NOR2x1_ASAP7_75t_SL g10177 ( 
.A(n_9708),
.B(n_572),
.Y(n_10177)
);

NAND2xp5_ASAP7_75t_L g10178 ( 
.A(n_9682),
.B(n_572),
.Y(n_10178)
);

OAI21x1_ASAP7_75t_L g10179 ( 
.A1(n_9727),
.A2(n_9631),
.B(n_9672),
.Y(n_10179)
);

NAND2xp5_ASAP7_75t_L g10180 ( 
.A(n_10080),
.B(n_572),
.Y(n_10180)
);

NAND2xp5_ASAP7_75t_L g10181 ( 
.A(n_9900),
.B(n_573),
.Y(n_10181)
);

AOI21xp5_ASAP7_75t_L g10182 ( 
.A1(n_9773),
.A2(n_573),
.B(n_574),
.Y(n_10182)
);

AOI21xp5_ASAP7_75t_L g10183 ( 
.A1(n_9874),
.A2(n_574),
.B(n_575),
.Y(n_10183)
);

AOI21xp5_ASAP7_75t_L g10184 ( 
.A1(n_9802),
.A2(n_574),
.B(n_575),
.Y(n_10184)
);

OAI21x1_ASAP7_75t_L g10185 ( 
.A1(n_9613),
.A2(n_575),
.B(n_576),
.Y(n_10185)
);

NAND2xp5_ASAP7_75t_L g10186 ( 
.A(n_9648),
.B(n_576),
.Y(n_10186)
);

A2O1A1Ixp33_ASAP7_75t_L g10187 ( 
.A1(n_9731),
.A2(n_578),
.B(n_576),
.C(n_577),
.Y(n_10187)
);

OR2x6_ASAP7_75t_L g10188 ( 
.A(n_9708),
.B(n_578),
.Y(n_10188)
);

NAND2xp5_ASAP7_75t_L g10189 ( 
.A(n_9677),
.B(n_578),
.Y(n_10189)
);

OAI21x1_ASAP7_75t_L g10190 ( 
.A1(n_9640),
.A2(n_579),
.B(n_580),
.Y(n_10190)
);

A2O1A1Ixp33_ASAP7_75t_L g10191 ( 
.A1(n_9632),
.A2(n_582),
.B(n_579),
.C(n_581),
.Y(n_10191)
);

AOI21xp5_ASAP7_75t_L g10192 ( 
.A1(n_9702),
.A2(n_579),
.B(n_581),
.Y(n_10192)
);

OAI21x1_ASAP7_75t_L g10193 ( 
.A1(n_9654),
.A2(n_581),
.B(n_582),
.Y(n_10193)
);

OAI22xp5_ASAP7_75t_L g10194 ( 
.A1(n_9665),
.A2(n_9898),
.B1(n_9914),
.B2(n_9899),
.Y(n_10194)
);

NAND2x1p5_ASAP7_75t_L g10195 ( 
.A(n_9610),
.B(n_582),
.Y(n_10195)
);

AOI21xp5_ASAP7_75t_L g10196 ( 
.A1(n_9710),
.A2(n_583),
.B(n_584),
.Y(n_10196)
);

NAND2xp5_ASAP7_75t_L g10197 ( 
.A(n_9678),
.B(n_583),
.Y(n_10197)
);

OAI21x1_ASAP7_75t_L g10198 ( 
.A1(n_9652),
.A2(n_583),
.B(n_585),
.Y(n_10198)
);

INVx1_ASAP7_75t_L g10199 ( 
.A(n_9721),
.Y(n_10199)
);

AOI21x1_ASAP7_75t_L g10200 ( 
.A1(n_9956),
.A2(n_585),
.B(n_586),
.Y(n_10200)
);

OAI21x1_ASAP7_75t_L g10201 ( 
.A1(n_10096),
.A2(n_585),
.B(n_586),
.Y(n_10201)
);

AOI21x1_ASAP7_75t_L g10202 ( 
.A1(n_9986),
.A2(n_586),
.B(n_588),
.Y(n_10202)
);

NOR2x1_ASAP7_75t_L g10203 ( 
.A(n_9878),
.B(n_588),
.Y(n_10203)
);

NAND2xp5_ASAP7_75t_L g10204 ( 
.A(n_9735),
.B(n_589),
.Y(n_10204)
);

NAND2xp5_ASAP7_75t_L g10205 ( 
.A(n_9746),
.B(n_589),
.Y(n_10205)
);

AOI21x1_ASAP7_75t_L g10206 ( 
.A1(n_9701),
.A2(n_589),
.B(n_590),
.Y(n_10206)
);

AOI21xp5_ASAP7_75t_L g10207 ( 
.A1(n_9629),
.A2(n_590),
.B(n_591),
.Y(n_10207)
);

OAI21xp5_ASAP7_75t_L g10208 ( 
.A1(n_9729),
.A2(n_591),
.B(n_592),
.Y(n_10208)
);

OAI21x1_ASAP7_75t_L g10209 ( 
.A1(n_10059),
.A2(n_592),
.B(n_593),
.Y(n_10209)
);

AOI21xp5_ASAP7_75t_L g10210 ( 
.A1(n_9769),
.A2(n_593),
.B(n_594),
.Y(n_10210)
);

OAI21x1_ASAP7_75t_L g10211 ( 
.A1(n_9912),
.A2(n_9650),
.B(n_9718),
.Y(n_10211)
);

OAI21x1_ASAP7_75t_SL g10212 ( 
.A1(n_9885),
.A2(n_594),
.B(n_595),
.Y(n_10212)
);

NAND2xp5_ASAP7_75t_L g10213 ( 
.A(n_9754),
.B(n_594),
.Y(n_10213)
);

OAI21x1_ASAP7_75t_L g10214 ( 
.A1(n_9724),
.A2(n_595),
.B(n_596),
.Y(n_10214)
);

AOI21xp5_ASAP7_75t_L g10215 ( 
.A1(n_9689),
.A2(n_595),
.B(n_596),
.Y(n_10215)
);

NAND2xp5_ASAP7_75t_L g10216 ( 
.A(n_9761),
.B(n_596),
.Y(n_10216)
);

A2O1A1Ixp33_ASAP7_75t_L g10217 ( 
.A1(n_9887),
.A2(n_599),
.B(n_597),
.C(n_598),
.Y(n_10217)
);

AOI22xp5_ASAP7_75t_L g10218 ( 
.A1(n_9698),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_10218)
);

OAI21x1_ASAP7_75t_L g10219 ( 
.A1(n_9644),
.A2(n_597),
.B(n_599),
.Y(n_10219)
);

BUFx12f_ASAP7_75t_L g10220 ( 
.A(n_9615),
.Y(n_10220)
);

BUFx3_ASAP7_75t_L g10221 ( 
.A(n_9870),
.Y(n_10221)
);

NAND2xp5_ASAP7_75t_L g10222 ( 
.A(n_9774),
.B(n_600),
.Y(n_10222)
);

A2O1A1Ixp33_ASAP7_75t_L g10223 ( 
.A1(n_9792),
.A2(n_602),
.B(n_600),
.C(n_601),
.Y(n_10223)
);

AOI21xp5_ASAP7_75t_L g10224 ( 
.A1(n_9875),
.A2(n_9653),
.B(n_9641),
.Y(n_10224)
);

AOI21xp5_ASAP7_75t_L g10225 ( 
.A1(n_9772),
.A2(n_600),
.B(n_601),
.Y(n_10225)
);

NAND2xp5_ASAP7_75t_L g10226 ( 
.A(n_9810),
.B(n_601),
.Y(n_10226)
);

AO21x2_ASAP7_75t_L g10227 ( 
.A1(n_10143),
.A2(n_602),
.B(n_603),
.Y(n_10227)
);

OAI21xp5_ASAP7_75t_L g10228 ( 
.A1(n_9825),
.A2(n_602),
.B(n_603),
.Y(n_10228)
);

AO31x2_ASAP7_75t_L g10229 ( 
.A1(n_9929),
.A2(n_605),
.A3(n_603),
.B(n_604),
.Y(n_10229)
);

OAI21x1_ASAP7_75t_L g10230 ( 
.A1(n_9737),
.A2(n_604),
.B(n_605),
.Y(n_10230)
);

AOI21xp5_ASAP7_75t_L g10231 ( 
.A1(n_9725),
.A2(n_10149),
.B(n_9663),
.Y(n_10231)
);

INVx2_ASAP7_75t_L g10232 ( 
.A(n_9993),
.Y(n_10232)
);

INVx2_ASAP7_75t_L g10233 ( 
.A(n_10007),
.Y(n_10233)
);

INVx1_ASAP7_75t_L g10234 ( 
.A(n_9827),
.Y(n_10234)
);

CKINVDCx5p33_ASAP7_75t_R g10235 ( 
.A(n_9612),
.Y(n_10235)
);

HB1xp67_ASAP7_75t_L g10236 ( 
.A(n_9848),
.Y(n_10236)
);

AND2x2_ASAP7_75t_L g10237 ( 
.A(n_10068),
.B(n_604),
.Y(n_10237)
);

INVx1_ASAP7_75t_L g10238 ( 
.A(n_9864),
.Y(n_10238)
);

AND2x2_ASAP7_75t_L g10239 ( 
.A(n_9968),
.B(n_606),
.Y(n_10239)
);

INVxp67_ASAP7_75t_SL g10240 ( 
.A(n_9628),
.Y(n_10240)
);

BUFx4_ASAP7_75t_SL g10241 ( 
.A(n_9713),
.Y(n_10241)
);

OAI21x1_ASAP7_75t_L g10242 ( 
.A1(n_9858),
.A2(n_606),
.B(n_607),
.Y(n_10242)
);

AOI21x1_ASAP7_75t_L g10243 ( 
.A1(n_9770),
.A2(n_606),
.B(n_607),
.Y(n_10243)
);

A2O1A1Ixp33_ASAP7_75t_L g10244 ( 
.A1(n_10070),
.A2(n_610),
.B(n_608),
.C(n_609),
.Y(n_10244)
);

AOI21xp5_ASAP7_75t_L g10245 ( 
.A1(n_9782),
.A2(n_608),
.B(n_609),
.Y(n_10245)
);

AO21x2_ASAP7_75t_L g10246 ( 
.A1(n_9926),
.A2(n_610),
.B(n_611),
.Y(n_10246)
);

OAI21x1_ASAP7_75t_L g10247 ( 
.A1(n_9892),
.A2(n_610),
.B(n_611),
.Y(n_10247)
);

AOI21xp5_ASAP7_75t_L g10248 ( 
.A1(n_9786),
.A2(n_612),
.B(n_613),
.Y(n_10248)
);

NAND2xp5_ASAP7_75t_L g10249 ( 
.A(n_9867),
.B(n_9869),
.Y(n_10249)
);

INVx2_ASAP7_75t_L g10250 ( 
.A(n_10017),
.Y(n_10250)
);

BUFx6f_ASAP7_75t_L g10251 ( 
.A(n_9646),
.Y(n_10251)
);

OAI21x1_ASAP7_75t_L g10252 ( 
.A1(n_9788),
.A2(n_612),
.B(n_613),
.Y(n_10252)
);

AOI21xp5_ASAP7_75t_L g10253 ( 
.A1(n_9688),
.A2(n_612),
.B(n_613),
.Y(n_10253)
);

OA22x2_ASAP7_75t_L g10254 ( 
.A1(n_9913),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_10254)
);

NAND3xp33_ASAP7_75t_SL g10255 ( 
.A(n_10131),
.B(n_615),
.C(n_616),
.Y(n_10255)
);

BUFx6f_ASAP7_75t_L g10256 ( 
.A(n_9646),
.Y(n_10256)
);

AOI21xp33_ASAP7_75t_L g10257 ( 
.A1(n_10060),
.A2(n_9951),
.B(n_9748),
.Y(n_10257)
);

OAI21x1_ASAP7_75t_L g10258 ( 
.A1(n_9813),
.A2(n_616),
.B(n_617),
.Y(n_10258)
);

HB1xp67_ASAP7_75t_L g10259 ( 
.A(n_9890),
.Y(n_10259)
);

OAI21x1_ASAP7_75t_SL g10260 ( 
.A1(n_9905),
.A2(n_9976),
.B(n_9711),
.Y(n_10260)
);

NAND2xp5_ASAP7_75t_L g10261 ( 
.A(n_9904),
.B(n_618),
.Y(n_10261)
);

OAI21x1_ASAP7_75t_L g10262 ( 
.A1(n_9856),
.A2(n_618),
.B(n_619),
.Y(n_10262)
);

AO21x1_ASAP7_75t_L g10263 ( 
.A1(n_10045),
.A2(n_618),
.B(n_619),
.Y(n_10263)
);

AOI21x1_ASAP7_75t_L g10264 ( 
.A1(n_9908),
.A2(n_9918),
.B(n_9911),
.Y(n_10264)
);

OA22x2_ASAP7_75t_L g10265 ( 
.A1(n_10118),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_10265)
);

AO31x2_ASAP7_75t_L g10266 ( 
.A1(n_9751),
.A2(n_622),
.A3(n_620),
.B(n_621),
.Y(n_10266)
);

NOR2x1_ASAP7_75t_R g10267 ( 
.A(n_9870),
.B(n_620),
.Y(n_10267)
);

NAND2xp5_ASAP7_75t_L g10268 ( 
.A(n_9909),
.B(n_621),
.Y(n_10268)
);

A2O1A1Ixp33_ASAP7_75t_L g10269 ( 
.A1(n_10111),
.A2(n_625),
.B(n_623),
.C(n_624),
.Y(n_10269)
);

NAND2xp5_ASAP7_75t_L g10270 ( 
.A(n_9916),
.B(n_623),
.Y(n_10270)
);

NOR2xp33_ASAP7_75t_R g10271 ( 
.A(n_9732),
.B(n_9621),
.Y(n_10271)
);

OAI21x1_ASAP7_75t_L g10272 ( 
.A1(n_9910),
.A2(n_623),
.B(n_624),
.Y(n_10272)
);

OAI21xp5_ASAP7_75t_L g10273 ( 
.A1(n_9687),
.A2(n_9690),
.B(n_9816),
.Y(n_10273)
);

OAI21x1_ASAP7_75t_L g10274 ( 
.A1(n_9936),
.A2(n_625),
.B(n_626),
.Y(n_10274)
);

BUFx6f_ASAP7_75t_L g10275 ( 
.A(n_9705),
.Y(n_10275)
);

AOI21x1_ASAP7_75t_L g10276 ( 
.A1(n_9923),
.A2(n_625),
.B(n_626),
.Y(n_10276)
);

NOR2x1_ASAP7_75t_SL g10277 ( 
.A(n_9907),
.B(n_627),
.Y(n_10277)
);

NAND3xp33_ASAP7_75t_L g10278 ( 
.A(n_9753),
.B(n_627),
.C(n_628),
.Y(n_10278)
);

OAI21x1_ASAP7_75t_L g10279 ( 
.A1(n_9831),
.A2(n_627),
.B(n_628),
.Y(n_10279)
);

OA21x2_ASAP7_75t_L g10280 ( 
.A1(n_9949),
.A2(n_628),
.B(n_629),
.Y(n_10280)
);

A2O1A1Ixp33_ASAP7_75t_L g10281 ( 
.A1(n_9965),
.A2(n_631),
.B(n_629),
.C(n_630),
.Y(n_10281)
);

OAI22xp33_ASAP7_75t_L g10282 ( 
.A1(n_9927),
.A2(n_631),
.B1(n_629),
.B2(n_630),
.Y(n_10282)
);

AND2x6_ASAP7_75t_L g10283 ( 
.A(n_10120),
.B(n_630),
.Y(n_10283)
);

AOI21x1_ASAP7_75t_L g10284 ( 
.A1(n_9925),
.A2(n_631),
.B(n_632),
.Y(n_10284)
);

CKINVDCx5p33_ASAP7_75t_R g10285 ( 
.A(n_9814),
.Y(n_10285)
);

OAI21x1_ASAP7_75t_L g10286 ( 
.A1(n_9840),
.A2(n_632),
.B(n_633),
.Y(n_10286)
);

A2O1A1Ixp33_ASAP7_75t_L g10287 ( 
.A1(n_9680),
.A2(n_635),
.B(n_633),
.C(n_634),
.Y(n_10287)
);

INVx4_ASAP7_75t_L g10288 ( 
.A(n_9622),
.Y(n_10288)
);

OAI21xp33_ASAP7_75t_L g10289 ( 
.A1(n_9692),
.A2(n_634),
.B(n_635),
.Y(n_10289)
);

NAND3xp33_ASAP7_75t_L g10290 ( 
.A(n_9970),
.B(n_636),
.C(n_637),
.Y(n_10290)
);

A2O1A1Ixp33_ASAP7_75t_L g10291 ( 
.A1(n_10014),
.A2(n_638),
.B(n_636),
.C(n_637),
.Y(n_10291)
);

INVx3_ASAP7_75t_SL g10292 ( 
.A(n_9728),
.Y(n_10292)
);

OAI21xp5_ASAP7_75t_L g10293 ( 
.A1(n_10006),
.A2(n_10150),
.B(n_9609),
.Y(n_10293)
);

OAI21x1_ASAP7_75t_L g10294 ( 
.A1(n_9661),
.A2(n_637),
.B(n_638),
.Y(n_10294)
);

A2O1A1Ixp33_ASAP7_75t_L g10295 ( 
.A1(n_10144),
.A2(n_640),
.B(n_638),
.C(n_639),
.Y(n_10295)
);

NOR2xp67_ASAP7_75t_L g10296 ( 
.A(n_10099),
.B(n_639),
.Y(n_10296)
);

NAND3xp33_ASAP7_75t_L g10297 ( 
.A(n_9861),
.B(n_640),
.C(n_641),
.Y(n_10297)
);

OAI21x1_ASAP7_75t_L g10298 ( 
.A1(n_9902),
.A2(n_642),
.B(n_643),
.Y(n_10298)
);

A2O1A1Ixp33_ASAP7_75t_L g10299 ( 
.A1(n_10030),
.A2(n_644),
.B(n_642),
.C(n_643),
.Y(n_10299)
);

OAI21xp5_ASAP7_75t_L g10300 ( 
.A1(n_9953),
.A2(n_642),
.B(n_643),
.Y(n_10300)
);

AOI21xp5_ASAP7_75t_L g10301 ( 
.A1(n_9673),
.A2(n_645),
.B(n_646),
.Y(n_10301)
);

AOI21xp5_ASAP7_75t_L g10302 ( 
.A1(n_9673),
.A2(n_645),
.B(n_646),
.Y(n_10302)
);

OAI21x1_ASAP7_75t_L g10303 ( 
.A1(n_10097),
.A2(n_645),
.B(n_646),
.Y(n_10303)
);

AOI21xp5_ASAP7_75t_L g10304 ( 
.A1(n_9797),
.A2(n_647),
.B(n_648),
.Y(n_10304)
);

OAI21x1_ASAP7_75t_L g10305 ( 
.A1(n_10121),
.A2(n_648),
.B(n_649),
.Y(n_10305)
);

OAI21xp5_ASAP7_75t_L g10306 ( 
.A1(n_9795),
.A2(n_9830),
.B(n_9759),
.Y(n_10306)
);

OAI21x1_ASAP7_75t_L g10307 ( 
.A1(n_9931),
.A2(n_648),
.B(n_649),
.Y(n_10307)
);

NAND2xp5_ASAP7_75t_L g10308 ( 
.A(n_9964),
.B(n_649),
.Y(n_10308)
);

NAND2xp5_ASAP7_75t_L g10309 ( 
.A(n_9971),
.B(n_650),
.Y(n_10309)
);

AOI22xp5_ASAP7_75t_L g10310 ( 
.A1(n_9614),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.Y(n_10310)
);

NAND2xp5_ASAP7_75t_L g10311 ( 
.A(n_9974),
.B(n_651),
.Y(n_10311)
);

OAI21xp5_ASAP7_75t_L g10312 ( 
.A1(n_9695),
.A2(n_651),
.B(n_652),
.Y(n_10312)
);

A2O1A1Ixp33_ASAP7_75t_L g10313 ( 
.A1(n_10115),
.A2(n_655),
.B(n_653),
.C(n_654),
.Y(n_10313)
);

OAI21x1_ASAP7_75t_L g10314 ( 
.A1(n_9934),
.A2(n_654),
.B(n_655),
.Y(n_10314)
);

NAND2xp5_ASAP7_75t_L g10315 ( 
.A(n_10009),
.B(n_654),
.Y(n_10315)
);

OAI21x1_ASAP7_75t_L g10316 ( 
.A1(n_9944),
.A2(n_656),
.B(n_657),
.Y(n_10316)
);

OAI21x1_ASAP7_75t_L g10317 ( 
.A1(n_9948),
.A2(n_656),
.B(n_657),
.Y(n_10317)
);

NOR2xp67_ASAP7_75t_L g10318 ( 
.A(n_10099),
.B(n_658),
.Y(n_10318)
);

AOI221xp5_ASAP7_75t_L g10319 ( 
.A1(n_9651),
.A2(n_660),
.B1(n_658),
.B2(n_659),
.C(n_661),
.Y(n_10319)
);

OAI21x1_ASAP7_75t_L g10320 ( 
.A1(n_9957),
.A2(n_658),
.B(n_659),
.Y(n_10320)
);

AOI22xp5_ASAP7_75t_L g10321 ( 
.A1(n_9675),
.A2(n_9801),
.B1(n_9893),
.B2(n_9975),
.Y(n_10321)
);

INVxp67_ASAP7_75t_L g10322 ( 
.A(n_10098),
.Y(n_10322)
);

OAI21xp5_ASAP7_75t_L g10323 ( 
.A1(n_9617),
.A2(n_660),
.B(n_662),
.Y(n_10323)
);

AND2x4_ASAP7_75t_L g10324 ( 
.A(n_9988),
.B(n_663),
.Y(n_10324)
);

NOR2xp67_ASAP7_75t_SL g10325 ( 
.A(n_10099),
.B(n_9808),
.Y(n_10325)
);

INVxp67_ASAP7_75t_L g10326 ( 
.A(n_10061),
.Y(n_10326)
);

OAI22xp5_ASAP7_75t_L g10327 ( 
.A1(n_9994),
.A2(n_665),
.B1(n_663),
.B2(n_664),
.Y(n_10327)
);

AND2x2_ASAP7_75t_L g10328 ( 
.A(n_10032),
.B(n_664),
.Y(n_10328)
);

AOI22xp5_ASAP7_75t_SL g10329 ( 
.A1(n_9919),
.A2(n_666),
.B1(n_664),
.B2(n_665),
.Y(n_10329)
);

AOI22xp5_ASAP7_75t_L g10330 ( 
.A1(n_10010),
.A2(n_667),
.B1(n_665),
.B2(n_666),
.Y(n_10330)
);

INVx1_ASAP7_75t_L g10331 ( 
.A(n_10018),
.Y(n_10331)
);

INVx1_ASAP7_75t_L g10332 ( 
.A(n_10037),
.Y(n_10332)
);

AOI21xp5_ASAP7_75t_L g10333 ( 
.A1(n_9797),
.A2(n_667),
.B(n_668),
.Y(n_10333)
);

INVx2_ASAP7_75t_L g10334 ( 
.A(n_10028),
.Y(n_10334)
);

AND2x2_ASAP7_75t_L g10335 ( 
.A(n_9939),
.B(n_667),
.Y(n_10335)
);

AOI22xp5_ASAP7_75t_L g10336 ( 
.A1(n_9871),
.A2(n_10001),
.B1(n_9618),
.B2(n_9668),
.Y(n_10336)
);

OAI21x1_ASAP7_75t_L g10337 ( 
.A1(n_9963),
.A2(n_668),
.B(n_669),
.Y(n_10337)
);

AO21x1_ASAP7_75t_L g10338 ( 
.A1(n_9978),
.A2(n_9979),
.B(n_9966),
.Y(n_10338)
);

OAI21x1_ASAP7_75t_L g10339 ( 
.A1(n_9981),
.A2(n_668),
.B(n_669),
.Y(n_10339)
);

OR2x6_ASAP7_75t_L g10340 ( 
.A(n_9907),
.B(n_670),
.Y(n_10340)
);

AOI21x1_ASAP7_75t_L g10341 ( 
.A1(n_9985),
.A2(n_670),
.B(n_671),
.Y(n_10341)
);

OAI21x1_ASAP7_75t_L g10342 ( 
.A1(n_9990),
.A2(n_670),
.B(n_672),
.Y(n_10342)
);

AOI21xp5_ASAP7_75t_L g10343 ( 
.A1(n_9821),
.A2(n_672),
.B(n_673),
.Y(n_10343)
);

NAND2x1_ASAP7_75t_L g10344 ( 
.A(n_9747),
.B(n_673),
.Y(n_10344)
);

NAND2xp5_ASAP7_75t_L g10345 ( 
.A(n_10108),
.B(n_673),
.Y(n_10345)
);

AOI21xp5_ASAP7_75t_L g10346 ( 
.A1(n_10138),
.A2(n_674),
.B(n_675),
.Y(n_10346)
);

NAND3xp33_ASAP7_75t_L g10347 ( 
.A(n_9736),
.B(n_9764),
.C(n_9757),
.Y(n_10347)
);

AOI21xp5_ASAP7_75t_L g10348 ( 
.A1(n_10138),
.A2(n_674),
.B(n_675),
.Y(n_10348)
);

NAND2xp5_ASAP7_75t_L g10349 ( 
.A(n_9947),
.B(n_675),
.Y(n_10349)
);

NAND3xp33_ASAP7_75t_L g10350 ( 
.A(n_9766),
.B(n_676),
.C(n_677),
.Y(n_10350)
);

AOI21xp5_ASAP7_75t_L g10351 ( 
.A1(n_9930),
.A2(n_676),
.B(n_678),
.Y(n_10351)
);

OAI21x1_ASAP7_75t_SL g10352 ( 
.A1(n_9997),
.A2(n_678),
.B(n_679),
.Y(n_10352)
);

OAI22x1_ASAP7_75t_L g10353 ( 
.A1(n_10119),
.A2(n_680),
.B1(n_678),
.B2(n_679),
.Y(n_10353)
);

AOI221xp5_ASAP7_75t_L g10354 ( 
.A1(n_9755),
.A2(n_682),
.B1(n_680),
.B2(n_681),
.C(n_683),
.Y(n_10354)
);

AOI21x1_ASAP7_75t_L g10355 ( 
.A1(n_9991),
.A2(n_681),
.B(n_682),
.Y(n_10355)
);

AND2x2_ASAP7_75t_L g10356 ( 
.A(n_9683),
.B(n_683),
.Y(n_10356)
);

OAI21x1_ASAP7_75t_L g10357 ( 
.A1(n_9995),
.A2(n_10005),
.B(n_9996),
.Y(n_10357)
);

OAI22xp5_ASAP7_75t_L g10358 ( 
.A1(n_9633),
.A2(n_685),
.B1(n_683),
.B2(n_684),
.Y(n_10358)
);

OAI21x1_ASAP7_75t_L g10359 ( 
.A1(n_9822),
.A2(n_684),
.B(n_686),
.Y(n_10359)
);

INVx3_ASAP7_75t_L g10360 ( 
.A(n_9705),
.Y(n_10360)
);

AND3x4_ASAP7_75t_L g10361 ( 
.A(n_9940),
.B(n_684),
.C(n_686),
.Y(n_10361)
);

AOI21xp5_ASAP7_75t_L g10362 ( 
.A1(n_10024),
.A2(n_687),
.B(n_688),
.Y(n_10362)
);

OAI21x1_ASAP7_75t_L g10363 ( 
.A1(n_10114),
.A2(n_687),
.B(n_688),
.Y(n_10363)
);

INVx2_ASAP7_75t_L g10364 ( 
.A(n_10035),
.Y(n_10364)
);

OAI21xp5_ASAP7_75t_L g10365 ( 
.A1(n_9846),
.A2(n_687),
.B(n_688),
.Y(n_10365)
);

BUFx12f_ASAP7_75t_L g10366 ( 
.A(n_9684),
.Y(n_10366)
);

OR2x2_ASAP7_75t_L g10367 ( 
.A(n_10047),
.B(n_689),
.Y(n_10367)
);

AOI21xp5_ASAP7_75t_L g10368 ( 
.A1(n_9733),
.A2(n_689),
.B(n_690),
.Y(n_10368)
);

AND2x4_ASAP7_75t_L g10369 ( 
.A(n_9793),
.B(n_689),
.Y(n_10369)
);

INVx2_ASAP7_75t_L g10370 ( 
.A(n_10039),
.Y(n_10370)
);

OR2x2_ASAP7_75t_L g10371 ( 
.A(n_9625),
.B(n_690),
.Y(n_10371)
);

OAI21x1_ASAP7_75t_L g10372 ( 
.A1(n_10117),
.A2(n_690),
.B(n_691),
.Y(n_10372)
);

OAI21x1_ASAP7_75t_L g10373 ( 
.A1(n_10122),
.A2(n_691),
.B(n_692),
.Y(n_10373)
);

BUFx3_ASAP7_75t_L g10374 ( 
.A(n_9722),
.Y(n_10374)
);

AOI21xp5_ASAP7_75t_L g10375 ( 
.A1(n_9844),
.A2(n_691),
.B(n_692),
.Y(n_10375)
);

AO21x1_ASAP7_75t_L g10376 ( 
.A1(n_9649),
.A2(n_692),
.B(n_693),
.Y(n_10376)
);

NAND2xp5_ASAP7_75t_L g10377 ( 
.A(n_9709),
.B(n_693),
.Y(n_10377)
);

BUFx2_ASAP7_75t_L g10378 ( 
.A(n_9730),
.Y(n_10378)
);

OA22x2_ASAP7_75t_L g10379 ( 
.A1(n_10011),
.A2(n_10051),
.B1(n_10085),
.B2(n_9849),
.Y(n_10379)
);

OAI21x1_ASAP7_75t_L g10380 ( 
.A1(n_10128),
.A2(n_693),
.B(n_694),
.Y(n_10380)
);

OAI21xp5_ASAP7_75t_L g10381 ( 
.A1(n_9681),
.A2(n_694),
.B(n_695),
.Y(n_10381)
);

A2O1A1Ixp33_ASAP7_75t_L g10382 ( 
.A1(n_10048),
.A2(n_10142),
.B(n_9946),
.C(n_9719),
.Y(n_10382)
);

INVx4_ASAP7_75t_L g10383 ( 
.A(n_9622),
.Y(n_10383)
);

NAND2xp5_ASAP7_75t_L g10384 ( 
.A(n_9809),
.B(n_9712),
.Y(n_10384)
);

OAI21xp5_ASAP7_75t_L g10385 ( 
.A1(n_9693),
.A2(n_694),
.B(n_695),
.Y(n_10385)
);

AOI21xp5_ASAP7_75t_L g10386 ( 
.A1(n_10073),
.A2(n_695),
.B(n_696),
.Y(n_10386)
);

INVx3_ASAP7_75t_L g10387 ( 
.A(n_9730),
.Y(n_10387)
);

OA21x2_ASAP7_75t_L g10388 ( 
.A1(n_9659),
.A2(n_696),
.B(n_697),
.Y(n_10388)
);

NAND2xp5_ASAP7_75t_L g10389 ( 
.A(n_9832),
.B(n_696),
.Y(n_10389)
);

NAND2xp5_ASAP7_75t_L g10390 ( 
.A(n_9660),
.B(n_697),
.Y(n_10390)
);

NOR2xp33_ASAP7_75t_SL g10391 ( 
.A(n_9863),
.B(n_697),
.Y(n_10391)
);

INVx4_ASAP7_75t_L g10392 ( 
.A(n_10004),
.Y(n_10392)
);

OAI21x1_ASAP7_75t_L g10393 ( 
.A1(n_10132),
.A2(n_698),
.B(n_699),
.Y(n_10393)
);

AOI21xp5_ASAP7_75t_L g10394 ( 
.A1(n_10073),
.A2(n_698),
.B(n_699),
.Y(n_10394)
);

OAI22x1_ASAP7_75t_L g10395 ( 
.A1(n_9604),
.A2(n_700),
.B1(n_698),
.B2(n_699),
.Y(n_10395)
);

INVx1_ASAP7_75t_L g10396 ( 
.A(n_10058),
.Y(n_10396)
);

AOI21xp5_ASAP7_75t_L g10397 ( 
.A1(n_10008),
.A2(n_700),
.B(n_702),
.Y(n_10397)
);

O2A1O1Ixp33_ASAP7_75t_L g10398 ( 
.A1(n_9778),
.A2(n_704),
.B(n_702),
.C(n_703),
.Y(n_10398)
);

NAND2xp5_ASAP7_75t_L g10399 ( 
.A(n_10041),
.B(n_9694),
.Y(n_10399)
);

OAI22xp5_ASAP7_75t_L g10400 ( 
.A1(n_9686),
.A2(n_704),
.B1(n_702),
.B2(n_703),
.Y(n_10400)
);

INVx2_ASAP7_75t_L g10401 ( 
.A(n_10042),
.Y(n_10401)
);

OAI21x1_ASAP7_75t_L g10402 ( 
.A1(n_9903),
.A2(n_703),
.B(n_705),
.Y(n_10402)
);

OAI21x1_ASAP7_75t_SL g10403 ( 
.A1(n_10022),
.A2(n_705),
.B(n_706),
.Y(n_10403)
);

AOI21x1_ASAP7_75t_L g10404 ( 
.A1(n_9819),
.A2(n_705),
.B(n_706),
.Y(n_10404)
);

A2O1A1Ixp33_ASAP7_75t_L g10405 ( 
.A1(n_9763),
.A2(n_708),
.B(n_706),
.C(n_707),
.Y(n_10405)
);

NAND2xp5_ASAP7_75t_L g10406 ( 
.A(n_9715),
.B(n_9706),
.Y(n_10406)
);

OAI21x1_ASAP7_75t_L g10407 ( 
.A1(n_9850),
.A2(n_707),
.B(n_708),
.Y(n_10407)
);

OAI21x1_ASAP7_75t_L g10408 ( 
.A1(n_9851),
.A2(n_707),
.B(n_708),
.Y(n_10408)
);

OAI22xp5_ASAP7_75t_L g10409 ( 
.A1(n_9771),
.A2(n_711),
.B1(n_709),
.B2(n_710),
.Y(n_10409)
);

OAI22xp5_ASAP7_75t_L g10410 ( 
.A1(n_10036),
.A2(n_712),
.B1(n_709),
.B2(n_710),
.Y(n_10410)
);

OAI21x1_ASAP7_75t_L g10411 ( 
.A1(n_9853),
.A2(n_710),
.B(n_712),
.Y(n_10411)
);

OAI21xp33_ASAP7_75t_SL g10412 ( 
.A1(n_10002),
.A2(n_712),
.B(n_713),
.Y(n_10412)
);

AND2x2_ASAP7_75t_L g10413 ( 
.A(n_10033),
.B(n_713),
.Y(n_10413)
);

NAND2xp5_ASAP7_75t_SL g10414 ( 
.A(n_10101),
.B(n_713),
.Y(n_10414)
);

OAI21x1_ASAP7_75t_L g10415 ( 
.A1(n_9857),
.A2(n_714),
.B(n_715),
.Y(n_10415)
);

CKINVDCx5p33_ASAP7_75t_R g10416 ( 
.A(n_9894),
.Y(n_10416)
);

AOI21xp5_ASAP7_75t_L g10417 ( 
.A1(n_9855),
.A2(n_715),
.B(n_716),
.Y(n_10417)
);

OAI21xp5_ASAP7_75t_L g10418 ( 
.A1(n_9860),
.A2(n_717),
.B(n_718),
.Y(n_10418)
);

NAND2xp5_ASAP7_75t_L g10419 ( 
.A(n_9723),
.B(n_9806),
.Y(n_10419)
);

O2A1O1Ixp5_ASAP7_75t_L g10420 ( 
.A1(n_9824),
.A2(n_719),
.B(n_717),
.C(n_718),
.Y(n_10420)
);

AO21x1_ASAP7_75t_L g10421 ( 
.A1(n_9917),
.A2(n_717),
.B(n_719),
.Y(n_10421)
);

INVx2_ASAP7_75t_L g10422 ( 
.A(n_10066),
.Y(n_10422)
);

OAI21x1_ASAP7_75t_L g10423 ( 
.A1(n_10129),
.A2(n_719),
.B(n_720),
.Y(n_10423)
);

OAI21x1_ASAP7_75t_L g10424 ( 
.A1(n_10130),
.A2(n_720),
.B(n_721),
.Y(n_10424)
);

NAND2x1p5_ASAP7_75t_L g10425 ( 
.A(n_9634),
.B(n_720),
.Y(n_10425)
);

AND2x2_ASAP7_75t_L g10426 ( 
.A(n_9696),
.B(n_721),
.Y(n_10426)
);

AOI21xp5_ASAP7_75t_L g10427 ( 
.A1(n_9933),
.A2(n_721),
.B(n_722),
.Y(n_10427)
);

BUFx12f_ASAP7_75t_L g10428 ( 
.A(n_10092),
.Y(n_10428)
);

INVx1_ASAP7_75t_L g10429 ( 
.A(n_10078),
.Y(n_10429)
);

NAND2xp5_ASAP7_75t_L g10430 ( 
.A(n_9608),
.B(n_722),
.Y(n_10430)
);

OAI21xp5_ASAP7_75t_L g10431 ( 
.A1(n_9636),
.A2(n_722),
.B(n_723),
.Y(n_10431)
);

NAND2xp5_ASAP7_75t_L g10432 ( 
.A(n_9611),
.B(n_9623),
.Y(n_10432)
);

AOI21x1_ASAP7_75t_L g10433 ( 
.A1(n_9656),
.A2(n_723),
.B(n_724),
.Y(n_10433)
);

AOI21xp5_ASAP7_75t_L g10434 ( 
.A1(n_9959),
.A2(n_723),
.B(n_724),
.Y(n_10434)
);

AOI22xp5_ASAP7_75t_L g10435 ( 
.A1(n_9749),
.A2(n_726),
.B1(n_724),
.B2(n_725),
.Y(n_10435)
);

AND2x4_ASAP7_75t_L g10436 ( 
.A(n_9637),
.B(n_725),
.Y(n_10436)
);

AND2x4_ASAP7_75t_L g10437 ( 
.A(n_10091),
.B(n_726),
.Y(n_10437)
);

AOI21xp5_ASAP7_75t_SL g10438 ( 
.A1(n_10139),
.A2(n_726),
.B(n_727),
.Y(n_10438)
);

INVx1_ASAP7_75t_L g10439 ( 
.A(n_10133),
.Y(n_10439)
);

AND2x2_ASAP7_75t_L g10440 ( 
.A(n_9697),
.B(n_727),
.Y(n_10440)
);

OAI21x1_ASAP7_75t_L g10441 ( 
.A1(n_10145),
.A2(n_728),
.B(n_729),
.Y(n_10441)
);

INVx2_ASAP7_75t_L g10442 ( 
.A(n_9616),
.Y(n_10442)
);

INVx2_ASAP7_75t_SL g10443 ( 
.A(n_10029),
.Y(n_10443)
);

AND2x4_ASAP7_75t_L g10444 ( 
.A(n_10141),
.B(n_728),
.Y(n_10444)
);

OAI21xp5_ASAP7_75t_L g10445 ( 
.A1(n_9691),
.A2(n_728),
.B(n_729),
.Y(n_10445)
);

AND2x2_ASAP7_75t_L g10446 ( 
.A(n_9833),
.B(n_730),
.Y(n_10446)
);

A2O1A1Ixp33_ASAP7_75t_L g10447 ( 
.A1(n_9873),
.A2(n_10124),
.B(n_10043),
.C(n_10057),
.Y(n_10447)
);

OAI21x1_ASAP7_75t_L g10448 ( 
.A1(n_10146),
.A2(n_730),
.B(n_731),
.Y(n_10448)
);

AO31x2_ASAP7_75t_L g10449 ( 
.A1(n_10135),
.A2(n_733),
.A3(n_731),
.B(n_732),
.Y(n_10449)
);

BUFx2_ASAP7_75t_L g10450 ( 
.A(n_9841),
.Y(n_10450)
);

OAI21x1_ASAP7_75t_L g10451 ( 
.A1(n_9627),
.A2(n_731),
.B(n_732),
.Y(n_10451)
);

NAND2xp5_ASAP7_75t_L g10452 ( 
.A(n_9635),
.B(n_9670),
.Y(n_10452)
);

AOI221xp5_ASAP7_75t_SL g10453 ( 
.A1(n_10113),
.A2(n_734),
.B1(n_732),
.B2(n_733),
.C(n_735),
.Y(n_10453)
);

NAND2xp5_ASAP7_75t_L g10454 ( 
.A(n_9720),
.B(n_734),
.Y(n_10454)
);

OR2x6_ASAP7_75t_L g10455 ( 
.A(n_9928),
.B(n_735),
.Y(n_10455)
);

AOI21xp33_ASAP7_75t_L g10456 ( 
.A1(n_9807),
.A2(n_736),
.B(n_737),
.Y(n_10456)
);

INVx4_ASAP7_75t_L g10457 ( 
.A(n_9765),
.Y(n_10457)
);

OAI21x1_ASAP7_75t_L g10458 ( 
.A1(n_10012),
.A2(n_736),
.B(n_738),
.Y(n_10458)
);

NOR2xp33_ASAP7_75t_R g10459 ( 
.A(n_9787),
.B(n_736),
.Y(n_10459)
);

AOI21xp5_ASAP7_75t_L g10460 ( 
.A1(n_10110),
.A2(n_738),
.B(n_739),
.Y(n_10460)
);

INVx2_ASAP7_75t_L g10461 ( 
.A(n_9626),
.Y(n_10461)
);

INVx1_ASAP7_75t_SL g10462 ( 
.A(n_10034),
.Y(n_10462)
);

AOI21x1_ASAP7_75t_L g10463 ( 
.A1(n_9664),
.A2(n_738),
.B(n_739),
.Y(n_10463)
);

OAI22x1_ASAP7_75t_L g10464 ( 
.A1(n_10102),
.A2(n_741),
.B1(n_739),
.B2(n_740),
.Y(n_10464)
);

AOI21xp5_ASAP7_75t_L g10465 ( 
.A1(n_10049),
.A2(n_740),
.B(n_741),
.Y(n_10465)
);

INVx3_ASAP7_75t_L g10466 ( 
.A(n_10029),
.Y(n_10466)
);

AOI21xp5_ASAP7_75t_L g10467 ( 
.A1(n_9915),
.A2(n_741),
.B(n_742),
.Y(n_10467)
);

NAND2xp5_ASAP7_75t_L g10468 ( 
.A(n_9674),
.B(n_742),
.Y(n_10468)
);

AO21x2_ASAP7_75t_L g10469 ( 
.A1(n_9739),
.A2(n_742),
.B(n_743),
.Y(n_10469)
);

NAND2xp5_ASAP7_75t_SL g10470 ( 
.A(n_10101),
.B(n_743),
.Y(n_10470)
);

A2O1A1Ixp33_ASAP7_75t_L g10471 ( 
.A1(n_10052),
.A2(n_746),
.B(n_744),
.C(n_745),
.Y(n_10471)
);

NOR2xp67_ASAP7_75t_L g10472 ( 
.A(n_9781),
.B(n_744),
.Y(n_10472)
);

AOI22xp33_ASAP7_75t_L g10473 ( 
.A1(n_9796),
.A2(n_746),
.B1(n_744),
.B2(n_745),
.Y(n_10473)
);

AOI21xp5_ASAP7_75t_L g10474 ( 
.A1(n_9779),
.A2(n_745),
.B(n_747),
.Y(n_10474)
);

OAI21x1_ASAP7_75t_L g10475 ( 
.A1(n_9843),
.A2(n_747),
.B(n_748),
.Y(n_10475)
);

AOI21xp5_ASAP7_75t_L g10476 ( 
.A1(n_9980),
.A2(n_747),
.B(n_748),
.Y(n_10476)
);

NAND2xp5_ASAP7_75t_L g10477 ( 
.A(n_9703),
.B(n_748),
.Y(n_10477)
);

INVx2_ASAP7_75t_L g10478 ( 
.A(n_9639),
.Y(n_10478)
);

NOR2xp33_ASAP7_75t_L g10479 ( 
.A(n_9790),
.B(n_749),
.Y(n_10479)
);

AOI22xp33_ASAP7_75t_L g10480 ( 
.A1(n_9796),
.A2(n_751),
.B1(n_749),
.B2(n_750),
.Y(n_10480)
);

AOI21x1_ASAP7_75t_L g10481 ( 
.A1(n_9667),
.A2(n_750),
.B(n_751),
.Y(n_10481)
);

INVx3_ASAP7_75t_L g10482 ( 
.A(n_9928),
.Y(n_10482)
);

NAND2xp5_ASAP7_75t_SL g10483 ( 
.A(n_10034),
.B(n_750),
.Y(n_10483)
);

INVx2_ASAP7_75t_L g10484 ( 
.A(n_9658),
.Y(n_10484)
);

AOI21xp5_ASAP7_75t_L g10485 ( 
.A1(n_9882),
.A2(n_751),
.B(n_752),
.Y(n_10485)
);

NAND2xp5_ASAP7_75t_L g10486 ( 
.A(n_9704),
.B(n_752),
.Y(n_10486)
);

INVx3_ASAP7_75t_L g10487 ( 
.A(n_9765),
.Y(n_10487)
);

OAI21x1_ASAP7_75t_SL g10488 ( 
.A1(n_9679),
.A2(n_752),
.B(n_753),
.Y(n_10488)
);

A2O1A1Ixp33_ASAP7_75t_L g10489 ( 
.A1(n_10062),
.A2(n_755),
.B(n_753),
.C(n_754),
.Y(n_10489)
);

NAND2xp5_ASAP7_75t_L g10490 ( 
.A(n_9638),
.B(n_753),
.Y(n_10490)
);

BUFx2_ASAP7_75t_L g10491 ( 
.A(n_10016),
.Y(n_10491)
);

BUFx4f_ASAP7_75t_L g10492 ( 
.A(n_9780),
.Y(n_10492)
);

OAI21x1_ASAP7_75t_L g10493 ( 
.A1(n_9950),
.A2(n_754),
.B(n_755),
.Y(n_10493)
);

OAI21x1_ASAP7_75t_L g10494 ( 
.A1(n_9967),
.A2(n_754),
.B(n_756),
.Y(n_10494)
);

NAND2xp33_ASAP7_75t_SL g10495 ( 
.A(n_9655),
.B(n_756),
.Y(n_10495)
);

NAND2x1p5_ASAP7_75t_L g10496 ( 
.A(n_9780),
.B(n_756),
.Y(n_10496)
);

AND2x6_ASAP7_75t_L g10497 ( 
.A(n_9791),
.B(n_757),
.Y(n_10497)
);

NAND2xp5_ASAP7_75t_L g10498 ( 
.A(n_9758),
.B(n_757),
.Y(n_10498)
);

AOI21xp5_ASAP7_75t_L g10499 ( 
.A1(n_10112),
.A2(n_757),
.B(n_758),
.Y(n_10499)
);

INVx1_ASAP7_75t_L g10500 ( 
.A(n_10140),
.Y(n_10500)
);

INVx3_ASAP7_75t_L g10501 ( 
.A(n_10072),
.Y(n_10501)
);

INVx1_ASAP7_75t_L g10502 ( 
.A(n_9685),
.Y(n_10502)
);

OAI22xp5_ASAP7_75t_L g10503 ( 
.A1(n_9606),
.A2(n_760),
.B1(n_758),
.B2(n_759),
.Y(n_10503)
);

AOI21x1_ASAP7_75t_L g10504 ( 
.A1(n_9738),
.A2(n_758),
.B(n_759),
.Y(n_10504)
);

NAND2xp5_ASAP7_75t_L g10505 ( 
.A(n_9762),
.B(n_9767),
.Y(n_10505)
);

HB1xp67_ASAP7_75t_L g10506 ( 
.A(n_10015),
.Y(n_10506)
);

NAND2xp5_ASAP7_75t_L g10507 ( 
.A(n_9768),
.B(n_759),
.Y(n_10507)
);

INVx2_ASAP7_75t_L g10508 ( 
.A(n_9714),
.Y(n_10508)
);

NOR2x1_ASAP7_75t_SL g10509 ( 
.A(n_9798),
.B(n_760),
.Y(n_10509)
);

AND3x2_ASAP7_75t_L g10510 ( 
.A(n_9987),
.B(n_761),
.C(n_762),
.Y(n_10510)
);

OAI21xp5_ASAP7_75t_L g10511 ( 
.A1(n_9969),
.A2(n_761),
.B(n_762),
.Y(n_10511)
);

BUFx12f_ASAP7_75t_L g10512 ( 
.A(n_10103),
.Y(n_10512)
);

AO21x1_ASAP7_75t_L g10513 ( 
.A1(n_9954),
.A2(n_761),
.B(n_762),
.Y(n_10513)
);

OAI21xp5_ASAP7_75t_L g10514 ( 
.A1(n_9977),
.A2(n_763),
.B(n_764),
.Y(n_10514)
);

INVx1_ASAP7_75t_L g10515 ( 
.A(n_9717),
.Y(n_10515)
);

OR2x2_ASAP7_75t_L g10516 ( 
.A(n_10040),
.B(n_763),
.Y(n_10516)
);

AOI21xp5_ASAP7_75t_SL g10517 ( 
.A1(n_9642),
.A2(n_764),
.B(n_765),
.Y(n_10517)
);

BUFx6f_ASAP7_75t_L g10518 ( 
.A(n_10089),
.Y(n_10518)
);

HB1xp67_ASAP7_75t_L g10519 ( 
.A(n_9865),
.Y(n_10519)
);

BUFx3_ASAP7_75t_L g10520 ( 
.A(n_10109),
.Y(n_10520)
);

OAI21x1_ASAP7_75t_L g10521 ( 
.A1(n_9982),
.A2(n_9989),
.B(n_9983),
.Y(n_10521)
);

AOI21xp5_ASAP7_75t_SL g10522 ( 
.A1(n_9643),
.A2(n_764),
.B(n_765),
.Y(n_10522)
);

AOI21xp5_ASAP7_75t_L g10523 ( 
.A1(n_9984),
.A2(n_765),
.B(n_766),
.Y(n_10523)
);

AO31x2_ASAP7_75t_L g10524 ( 
.A1(n_9726),
.A2(n_768),
.A3(n_766),
.B(n_767),
.Y(n_10524)
);

AND3x1_ASAP7_75t_SL g10525 ( 
.A(n_9958),
.B(n_766),
.C(n_768),
.Y(n_10525)
);

AND2x6_ASAP7_75t_L g10526 ( 
.A(n_10021),
.B(n_768),
.Y(n_10526)
);

OAI21x1_ASAP7_75t_L g10527 ( 
.A1(n_10003),
.A2(n_769),
.B(n_770),
.Y(n_10527)
);

AOI21x1_ASAP7_75t_L g10528 ( 
.A1(n_9744),
.A2(n_769),
.B(n_770),
.Y(n_10528)
);

INVx8_ASAP7_75t_L g10529 ( 
.A(n_9798),
.Y(n_10529)
);

NAND2xp5_ASAP7_75t_L g10530 ( 
.A(n_9866),
.B(n_769),
.Y(n_10530)
);

OAI21x1_ASAP7_75t_L g10531 ( 
.A1(n_10019),
.A2(n_770),
.B(n_771),
.Y(n_10531)
);

AOI21xp5_ASAP7_75t_L g10532 ( 
.A1(n_9699),
.A2(n_772),
.B(n_773),
.Y(n_10532)
);

AOI21xp5_ASAP7_75t_L g10533 ( 
.A1(n_9750),
.A2(n_772),
.B(n_773),
.Y(n_10533)
);

INVx3_ASAP7_75t_L g10534 ( 
.A(n_9666),
.Y(n_10534)
);

NOR2x1_ASAP7_75t_SL g10535 ( 
.A(n_9803),
.B(n_772),
.Y(n_10535)
);

AO21x1_ASAP7_75t_L g10536 ( 
.A1(n_9794),
.A2(n_773),
.B(n_774),
.Y(n_10536)
);

INVx1_ASAP7_75t_L g10537 ( 
.A(n_9734),
.Y(n_10537)
);

BUFx3_ASAP7_75t_L g10538 ( 
.A(n_9796),
.Y(n_10538)
);

OAI22xp5_ASAP7_75t_L g10539 ( 
.A1(n_10088),
.A2(n_776),
.B1(n_774),
.B2(n_775),
.Y(n_10539)
);

INVx3_ASAP7_75t_L g10540 ( 
.A(n_10148),
.Y(n_10540)
);

INVx2_ASAP7_75t_L g10541 ( 
.A(n_9741),
.Y(n_10541)
);

AND2x4_ASAP7_75t_L g10542 ( 
.A(n_9742),
.B(n_775),
.Y(n_10542)
);

AOI21xp5_ASAP7_75t_L g10543 ( 
.A1(n_9669),
.A2(n_775),
.B(n_776),
.Y(n_10543)
);

BUFx2_ASAP7_75t_R g10544 ( 
.A(n_10056),
.Y(n_10544)
);

INVx3_ASAP7_75t_SL g10545 ( 
.A(n_10125),
.Y(n_10545)
);

OAI21x1_ASAP7_75t_L g10546 ( 
.A1(n_10020),
.A2(n_777),
.B(n_778),
.Y(n_10546)
);

NAND2xp5_ASAP7_75t_L g10547 ( 
.A(n_9872),
.B(n_9877),
.Y(n_10547)
);

OAI21x1_ASAP7_75t_L g10548 ( 
.A1(n_10023),
.A2(n_777),
.B(n_779),
.Y(n_10548)
);

AOI21xp5_ASAP7_75t_L g10549 ( 
.A1(n_10123),
.A2(n_779),
.B(n_780),
.Y(n_10549)
);

INVx3_ASAP7_75t_L g10550 ( 
.A(n_9932),
.Y(n_10550)
);

OAI21x1_ASAP7_75t_L g10551 ( 
.A1(n_10026),
.A2(n_779),
.B(n_780),
.Y(n_10551)
);

NOR2xp33_ASAP7_75t_SL g10552 ( 
.A(n_9823),
.B(n_780),
.Y(n_10552)
);

OAI21x1_ASAP7_75t_L g10553 ( 
.A1(n_9889),
.A2(n_781),
.B(n_782),
.Y(n_10553)
);

NAND2xp5_ASAP7_75t_SL g10554 ( 
.A(n_10000),
.B(n_782),
.Y(n_10554)
);

INVx2_ASAP7_75t_L g10555 ( 
.A(n_9785),
.Y(n_10555)
);

NAND2xp5_ASAP7_75t_L g10556 ( 
.A(n_9897),
.B(n_783),
.Y(n_10556)
);

NAND2xp5_ASAP7_75t_L g10557 ( 
.A(n_9776),
.B(n_783),
.Y(n_10557)
);

NAND2xp5_ASAP7_75t_L g10558 ( 
.A(n_9777),
.B(n_783),
.Y(n_10558)
);

AND2x2_ASAP7_75t_L g10559 ( 
.A(n_9829),
.B(n_784),
.Y(n_10559)
);

AOI21xp5_ASAP7_75t_L g10560 ( 
.A1(n_10126),
.A2(n_784),
.B(n_785),
.Y(n_10560)
);

AOI21xp5_ASAP7_75t_L g10561 ( 
.A1(n_9700),
.A2(n_785),
.B(n_786),
.Y(n_10561)
);

NAND2xp5_ASAP7_75t_L g10562 ( 
.A(n_9784),
.B(n_786),
.Y(n_10562)
);

NAND2xp5_ASAP7_75t_L g10563 ( 
.A(n_9804),
.B(n_786),
.Y(n_10563)
);

NAND2xp5_ASAP7_75t_L g10564 ( 
.A(n_9805),
.B(n_787),
.Y(n_10564)
);

AOI21xp5_ASAP7_75t_L g10565 ( 
.A1(n_9745),
.A2(n_788),
.B(n_789),
.Y(n_10565)
);

HB1xp67_ASAP7_75t_L g10566 ( 
.A(n_9838),
.Y(n_10566)
);

A2O1A1Ixp33_ASAP7_75t_L g10567 ( 
.A1(n_10063),
.A2(n_791),
.B(n_788),
.C(n_790),
.Y(n_10567)
);

AOI21xp5_ASAP7_75t_L g10568 ( 
.A1(n_9895),
.A2(n_788),
.B(n_790),
.Y(n_10568)
);

O2A1O1Ixp5_ASAP7_75t_L g10569 ( 
.A1(n_9760),
.A2(n_9789),
.B(n_9906),
.C(n_9891),
.Y(n_10569)
);

INVx1_ASAP7_75t_L g10570 ( 
.A(n_9847),
.Y(n_10570)
);

NAND2xp5_ASAP7_75t_L g10571 ( 
.A(n_9815),
.B(n_792),
.Y(n_10571)
);

AOI21xp5_ASAP7_75t_L g10572 ( 
.A1(n_9973),
.A2(n_792),
.B(n_793),
.Y(n_10572)
);

AOI21xp33_ASAP7_75t_L g10573 ( 
.A1(n_9992),
.A2(n_792),
.B(n_793),
.Y(n_10573)
);

AOI21xp5_ASAP7_75t_L g10574 ( 
.A1(n_9998),
.A2(n_793),
.B(n_794),
.Y(n_10574)
);

NOR2xp33_ASAP7_75t_SL g10575 ( 
.A(n_10031),
.B(n_794),
.Y(n_10575)
);

NAND2xp5_ASAP7_75t_L g10576 ( 
.A(n_9817),
.B(n_9818),
.Y(n_10576)
);

NAND2xp5_ASAP7_75t_L g10577 ( 
.A(n_9835),
.B(n_794),
.Y(n_10577)
);

AND2x4_ASAP7_75t_L g10578 ( 
.A(n_9868),
.B(n_795),
.Y(n_10578)
);

INVx4_ASAP7_75t_L g10579 ( 
.A(n_9972),
.Y(n_10579)
);

NAND2xp5_ASAP7_75t_L g10580 ( 
.A(n_9836),
.B(n_795),
.Y(n_10580)
);

NAND2xp5_ASAP7_75t_L g10581 ( 
.A(n_9837),
.B(n_796),
.Y(n_10581)
);

AO31x2_ASAP7_75t_L g10582 ( 
.A1(n_9883),
.A2(n_799),
.A3(n_797),
.B(n_798),
.Y(n_10582)
);

INVx3_ASAP7_75t_L g10583 ( 
.A(n_9886),
.Y(n_10583)
);

NOR2xp67_ASAP7_75t_L g10584 ( 
.A(n_9845),
.B(n_797),
.Y(n_10584)
);

NAND2xp5_ASAP7_75t_L g10585 ( 
.A(n_9859),
.B(n_797),
.Y(n_10585)
);

AOI221xp5_ASAP7_75t_SL g10586 ( 
.A1(n_9941),
.A2(n_800),
.B1(n_798),
.B2(n_799),
.C(n_801),
.Y(n_10586)
);

AOI22xp33_ASAP7_75t_L g10587 ( 
.A1(n_10054),
.A2(n_800),
.B1(n_798),
.B2(n_799),
.Y(n_10587)
);

AO31x2_ASAP7_75t_L g10588 ( 
.A1(n_9921),
.A2(n_802),
.A3(n_800),
.B(n_801),
.Y(n_10588)
);

INVx2_ASAP7_75t_L g10589 ( 
.A(n_9937),
.Y(n_10589)
);

AND2x2_ASAP7_75t_L g10590 ( 
.A(n_9943),
.B(n_801),
.Y(n_10590)
);

OAI21x1_ASAP7_75t_L g10591 ( 
.A1(n_9876),
.A2(n_802),
.B(n_803),
.Y(n_10591)
);

AOI21xp5_ASAP7_75t_L g10592 ( 
.A1(n_10025),
.A2(n_802),
.B(n_803),
.Y(n_10592)
);

AND2x2_ASAP7_75t_L g10593 ( 
.A(n_9952),
.B(n_803),
.Y(n_10593)
);

OAI21x1_ASAP7_75t_L g10594 ( 
.A1(n_9879),
.A2(n_804),
.B(n_805),
.Y(n_10594)
);

NAND2xp5_ASAP7_75t_SL g10595 ( 
.A(n_10147),
.B(n_804),
.Y(n_10595)
);

BUFx12f_ASAP7_75t_L g10596 ( 
.A(n_10106),
.Y(n_10596)
);

AOI21x1_ASAP7_75t_L g10597 ( 
.A1(n_9922),
.A2(n_9924),
.B(n_9862),
.Y(n_10597)
);

NAND2xp5_ASAP7_75t_L g10598 ( 
.A(n_10053),
.B(n_804),
.Y(n_10598)
);

INVx2_ASAP7_75t_L g10599 ( 
.A(n_9938),
.Y(n_10599)
);

AOI21xp5_ASAP7_75t_L g10600 ( 
.A1(n_9888),
.A2(n_805),
.B(n_806),
.Y(n_10600)
);

OAI21x1_ASAP7_75t_L g10601 ( 
.A1(n_9896),
.A2(n_806),
.B(n_807),
.Y(n_10601)
);

INVx5_ASAP7_75t_L g10602 ( 
.A(n_10137),
.Y(n_10602)
);

OAI22x1_ASAP7_75t_L g10603 ( 
.A1(n_9834),
.A2(n_808),
.B1(n_806),
.B2(n_807),
.Y(n_10603)
);

NAND2xp5_ASAP7_75t_L g10604 ( 
.A(n_10084),
.B(n_807),
.Y(n_10604)
);

AOI21xp5_ASAP7_75t_L g10605 ( 
.A1(n_10136),
.A2(n_808),
.B(n_809),
.Y(n_10605)
);

INVx1_ASAP7_75t_L g10606 ( 
.A(n_9945),
.Y(n_10606)
);

AOI21xp5_ASAP7_75t_L g10607 ( 
.A1(n_9901),
.A2(n_808),
.B(n_809),
.Y(n_10607)
);

OAI21x1_ASAP7_75t_L g10608 ( 
.A1(n_9740),
.A2(n_809),
.B(n_810),
.Y(n_10608)
);

NAND2xp5_ASAP7_75t_SL g10609 ( 
.A(n_10013),
.B(n_810),
.Y(n_10609)
);

NAND2xp5_ASAP7_75t_L g10610 ( 
.A(n_10086),
.B(n_810),
.Y(n_10610)
);

NAND2xp5_ASAP7_75t_L g10611 ( 
.A(n_10044),
.B(n_811),
.Y(n_10611)
);

AOI21xp5_ASAP7_75t_L g10612 ( 
.A1(n_9743),
.A2(n_811),
.B(n_812),
.Y(n_10612)
);

INVx3_ASAP7_75t_L g10613 ( 
.A(n_10071),
.Y(n_10613)
);

AO31x2_ASAP7_75t_L g10614 ( 
.A1(n_10075),
.A2(n_814),
.A3(n_812),
.B(n_813),
.Y(n_10614)
);

NAND2xp5_ASAP7_75t_L g10615 ( 
.A(n_10105),
.B(n_813),
.Y(n_10615)
);

NOR2xp33_ASAP7_75t_L g10616 ( 
.A(n_9828),
.B(n_813),
.Y(n_10616)
);

OAI21x1_ASAP7_75t_L g10617 ( 
.A1(n_9756),
.A2(n_10064),
.B(n_9942),
.Y(n_10617)
);

OAI21x1_ASAP7_75t_SL g10618 ( 
.A1(n_10116),
.A2(n_814),
.B(n_815),
.Y(n_10618)
);

INVx2_ASAP7_75t_L g10619 ( 
.A(n_10076),
.Y(n_10619)
);

OAI21xp5_ASAP7_75t_L g10620 ( 
.A1(n_10067),
.A2(n_814),
.B(n_815),
.Y(n_10620)
);

AO221x1_ASAP7_75t_L g10621 ( 
.A1(n_9880),
.A2(n_818),
.B1(n_816),
.B2(n_817),
.C(n_819),
.Y(n_10621)
);

OAI21xp5_ASAP7_75t_L g10622 ( 
.A1(n_10069),
.A2(n_816),
.B(n_817),
.Y(n_10622)
);

INVx2_ASAP7_75t_SL g10623 ( 
.A(n_10038),
.Y(n_10623)
);

OAI21xp33_ASAP7_75t_L g10624 ( 
.A1(n_10074),
.A2(n_816),
.B(n_818),
.Y(n_10624)
);

NAND2xp5_ASAP7_75t_L g10625 ( 
.A(n_10055),
.B(n_818),
.Y(n_10625)
);

AOI21xp5_ASAP7_75t_L g10626 ( 
.A1(n_10077),
.A2(n_819),
.B(n_820),
.Y(n_10626)
);

NAND2xp5_ASAP7_75t_SL g10627 ( 
.A(n_9881),
.B(n_819),
.Y(n_10627)
);

NAND2xp5_ASAP7_75t_L g10628 ( 
.A(n_10027),
.B(n_820),
.Y(n_10628)
);

NAND2xp5_ASAP7_75t_L g10629 ( 
.A(n_9826),
.B(n_821),
.Y(n_10629)
);

INVx1_ASAP7_75t_L g10630 ( 
.A(n_10127),
.Y(n_10630)
);

NAND2xp5_ASAP7_75t_L g10631 ( 
.A(n_9852),
.B(n_821),
.Y(n_10631)
);

AOI21xp5_ASAP7_75t_L g10632 ( 
.A1(n_10090),
.A2(n_821),
.B(n_822),
.Y(n_10632)
);

INVx1_ASAP7_75t_L g10633 ( 
.A(n_10079),
.Y(n_10633)
);

NAND2xp5_ASAP7_75t_L g10634 ( 
.A(n_9884),
.B(n_822),
.Y(n_10634)
);

AOI22xp5_ASAP7_75t_L g10635 ( 
.A1(n_10065),
.A2(n_9961),
.B1(n_9955),
.B2(n_9999),
.Y(n_10635)
);

OAI21x1_ASAP7_75t_L g10636 ( 
.A1(n_10094),
.A2(n_823),
.B(n_824),
.Y(n_10636)
);

OAI21x1_ASAP7_75t_L g10637 ( 
.A1(n_10100),
.A2(n_823),
.B(n_824),
.Y(n_10637)
);

A2O1A1Ixp33_ASAP7_75t_L g10638 ( 
.A1(n_10104),
.A2(n_10050),
.B(n_9800),
.C(n_9811),
.Y(n_10638)
);

NAND2x1p5_ASAP7_75t_L g10639 ( 
.A(n_10081),
.B(n_823),
.Y(n_10639)
);

NAND2x1p5_ASAP7_75t_L g10640 ( 
.A(n_10082),
.B(n_825),
.Y(n_10640)
);

NAND2xp5_ASAP7_75t_SL g10641 ( 
.A(n_10046),
.B(n_825),
.Y(n_10641)
);

INVx1_ASAP7_75t_L g10642 ( 
.A(n_10083),
.Y(n_10642)
);

NAND2x1p5_ASAP7_75t_L g10643 ( 
.A(n_10095),
.B(n_826),
.Y(n_10643)
);

INVx2_ASAP7_75t_L g10644 ( 
.A(n_10107),
.Y(n_10644)
);

AOI21x1_ASAP7_75t_L g10645 ( 
.A1(n_9799),
.A2(n_826),
.B(n_827),
.Y(n_10645)
);

INVx2_ASAP7_75t_L g10646 ( 
.A(n_10093),
.Y(n_10646)
);

INVx1_ASAP7_75t_L g10647 ( 
.A(n_10087),
.Y(n_10647)
);

AOI221x1_ASAP7_75t_L g10648 ( 
.A1(n_10479),
.A2(n_9820),
.B1(n_9812),
.B2(n_829),
.C(n_827),
.Y(n_10648)
);

AOI21xp5_ASAP7_75t_L g10649 ( 
.A1(n_10231),
.A2(n_827),
.B(n_828),
.Y(n_10649)
);

AOI21xp5_ASAP7_75t_L g10650 ( 
.A1(n_10224),
.A2(n_828),
.B(n_830),
.Y(n_10650)
);

NAND3x1_ASAP7_75t_L g10651 ( 
.A(n_10335),
.B(n_828),
.C(n_830),
.Y(n_10651)
);

INVx1_ASAP7_75t_L g10652 ( 
.A(n_10236),
.Y(n_10652)
);

OAI21x1_ASAP7_75t_L g10653 ( 
.A1(n_10179),
.A2(n_831),
.B(n_832),
.Y(n_10653)
);

BUFx6f_ASAP7_75t_L g10654 ( 
.A(n_10275),
.Y(n_10654)
);

AOI21xp5_ASAP7_75t_L g10655 ( 
.A1(n_10273),
.A2(n_831),
.B(n_832),
.Y(n_10655)
);

INVx1_ASAP7_75t_L g10656 ( 
.A(n_10259),
.Y(n_10656)
);

NAND2xp5_ASAP7_75t_L g10657 ( 
.A(n_10157),
.B(n_832),
.Y(n_10657)
);

BUFx2_ASAP7_75t_L g10658 ( 
.A(n_10450),
.Y(n_10658)
);

OAI22xp5_ASAP7_75t_L g10659 ( 
.A1(n_10321),
.A2(n_10336),
.B1(n_10480),
.B2(n_10473),
.Y(n_10659)
);

INVx3_ASAP7_75t_L g10660 ( 
.A(n_10275),
.Y(n_10660)
);

AOI21xp5_ASAP7_75t_L g10661 ( 
.A1(n_10184),
.A2(n_833),
.B(n_834),
.Y(n_10661)
);

OAI21xp5_ASAP7_75t_L g10662 ( 
.A1(n_10228),
.A2(n_833),
.B(n_834),
.Y(n_10662)
);

OAI21x1_ASAP7_75t_L g10663 ( 
.A1(n_10264),
.A2(n_833),
.B(n_835),
.Y(n_10663)
);

AO31x2_ASAP7_75t_L g10664 ( 
.A1(n_10338),
.A2(n_837),
.A3(n_835),
.B(n_836),
.Y(n_10664)
);

NAND2xp5_ASAP7_75t_L g10665 ( 
.A(n_10169),
.B(n_835),
.Y(n_10665)
);

O2A1O1Ixp5_ASAP7_75t_SL g10666 ( 
.A1(n_10506),
.A2(n_839),
.B(n_837),
.C(n_838),
.Y(n_10666)
);

INVx2_ASAP7_75t_L g10667 ( 
.A(n_10422),
.Y(n_10667)
);

NOR2xp33_ASAP7_75t_SL g10668 ( 
.A(n_10155),
.B(n_837),
.Y(n_10668)
);

AOI21xp33_ASAP7_75t_L g10669 ( 
.A1(n_10260),
.A2(n_838),
.B(n_839),
.Y(n_10669)
);

AOI21xp33_ASAP7_75t_L g10670 ( 
.A1(n_10246),
.A2(n_840),
.B(n_841),
.Y(n_10670)
);

OR2x6_ASAP7_75t_L g10671 ( 
.A(n_10538),
.B(n_10529),
.Y(n_10671)
);

OAI21x1_ASAP7_75t_L g10672 ( 
.A1(n_10357),
.A2(n_841),
.B(n_842),
.Y(n_10672)
);

AO21x2_ASAP7_75t_L g10673 ( 
.A1(n_10186),
.A2(n_841),
.B(n_842),
.Y(n_10673)
);

NAND2xp5_ASAP7_75t_L g10674 ( 
.A(n_10240),
.B(n_842),
.Y(n_10674)
);

AOI21xp5_ASAP7_75t_L g10675 ( 
.A1(n_10293),
.A2(n_843),
.B(n_844),
.Y(n_10675)
);

OAI21x1_ASAP7_75t_SL g10676 ( 
.A1(n_10177),
.A2(n_843),
.B(n_844),
.Y(n_10676)
);

AO21x1_ASAP7_75t_L g10677 ( 
.A1(n_10552),
.A2(n_844),
.B(n_845),
.Y(n_10677)
);

OAI21x1_ASAP7_75t_L g10678 ( 
.A1(n_10211),
.A2(n_10200),
.B(n_10252),
.Y(n_10678)
);

AND2x2_ASAP7_75t_L g10679 ( 
.A(n_10322),
.B(n_10168),
.Y(n_10679)
);

OAI21x1_ASAP7_75t_L g10680 ( 
.A1(n_10258),
.A2(n_845),
.B(n_846),
.Y(n_10680)
);

NAND2x1p5_ASAP7_75t_L g10681 ( 
.A(n_10325),
.B(n_845),
.Y(n_10681)
);

NAND2xp5_ASAP7_75t_SL g10682 ( 
.A(n_10602),
.B(n_846),
.Y(n_10682)
);

O2A1O1Ixp33_ASAP7_75t_L g10683 ( 
.A1(n_10299),
.A2(n_849),
.B(n_847),
.C(n_848),
.Y(n_10683)
);

OAI21xp5_ASAP7_75t_L g10684 ( 
.A1(n_10183),
.A2(n_847),
.B(n_848),
.Y(n_10684)
);

OAI21xp5_ASAP7_75t_L g10685 ( 
.A1(n_10182),
.A2(n_847),
.B(n_849),
.Y(n_10685)
);

OAI21xp5_ASAP7_75t_L g10686 ( 
.A1(n_10210),
.A2(n_10207),
.B(n_10160),
.Y(n_10686)
);

AND2x2_ASAP7_75t_L g10687 ( 
.A(n_10534),
.B(n_849),
.Y(n_10687)
);

NAND2xp5_ASAP7_75t_L g10688 ( 
.A(n_10174),
.B(n_850),
.Y(n_10688)
);

INVx1_ASAP7_75t_SL g10689 ( 
.A(n_10271),
.Y(n_10689)
);

OAI21x1_ASAP7_75t_L g10690 ( 
.A1(n_10262),
.A2(n_850),
.B(n_851),
.Y(n_10690)
);

INVxp67_ASAP7_75t_SL g10691 ( 
.A(n_10326),
.Y(n_10691)
);

NOR4xp25_ASAP7_75t_L g10692 ( 
.A(n_10289),
.B(n_853),
.C(n_851),
.D(n_852),
.Y(n_10692)
);

AOI221xp5_ASAP7_75t_L g10693 ( 
.A1(n_10257),
.A2(n_854),
.B1(n_852),
.B2(n_853),
.C(n_855),
.Y(n_10693)
);

OAI21x1_ASAP7_75t_L g10694 ( 
.A1(n_10167),
.A2(n_852),
.B(n_854),
.Y(n_10694)
);

NAND2xp5_ASAP7_75t_L g10695 ( 
.A(n_10519),
.B(n_856),
.Y(n_10695)
);

INVx3_ASAP7_75t_L g10696 ( 
.A(n_10457),
.Y(n_10696)
);

OAI21x1_ASAP7_75t_L g10697 ( 
.A1(n_10521),
.A2(n_856),
.B(n_857),
.Y(n_10697)
);

INVx1_ASAP7_75t_L g10698 ( 
.A(n_10249),
.Y(n_10698)
);

AOI211x1_ASAP7_75t_L g10699 ( 
.A1(n_10263),
.A2(n_858),
.B(n_856),
.C(n_857),
.Y(n_10699)
);

OAI21x1_ASAP7_75t_L g10700 ( 
.A1(n_10165),
.A2(n_857),
.B(n_858),
.Y(n_10700)
);

NAND2xp5_ASAP7_75t_L g10701 ( 
.A(n_10199),
.B(n_858),
.Y(n_10701)
);

INVx3_ASAP7_75t_L g10702 ( 
.A(n_10221),
.Y(n_10702)
);

AOI22xp5_ASAP7_75t_L g10703 ( 
.A1(n_10283),
.A2(n_861),
.B1(n_859),
.B2(n_860),
.Y(n_10703)
);

OA21x2_ASAP7_75t_L g10704 ( 
.A1(n_10189),
.A2(n_859),
.B(n_860),
.Y(n_10704)
);

NOR2x1_ASAP7_75t_R g10705 ( 
.A(n_10220),
.B(n_861),
.Y(n_10705)
);

INVx1_ASAP7_75t_L g10706 ( 
.A(n_10234),
.Y(n_10706)
);

OAI21x1_ASAP7_75t_L g10707 ( 
.A1(n_10206),
.A2(n_861),
.B(n_862),
.Y(n_10707)
);

INVx1_ASAP7_75t_L g10708 ( 
.A(n_10238),
.Y(n_10708)
);

OAI21x1_ASAP7_75t_L g10709 ( 
.A1(n_10276),
.A2(n_863),
.B(n_864),
.Y(n_10709)
);

OR2x6_ASAP7_75t_L g10710 ( 
.A(n_10529),
.B(n_863),
.Y(n_10710)
);

INVx2_ASAP7_75t_L g10711 ( 
.A(n_10156),
.Y(n_10711)
);

AOI21xp5_ASAP7_75t_SL g10712 ( 
.A1(n_10277),
.A2(n_864),
.B(n_865),
.Y(n_10712)
);

AO21x2_ASAP7_75t_L g10713 ( 
.A1(n_10197),
.A2(n_865),
.B(n_866),
.Y(n_10713)
);

INVx1_ASAP7_75t_L g10714 ( 
.A(n_10331),
.Y(n_10714)
);

AOI21xp5_ASAP7_75t_L g10715 ( 
.A1(n_10194),
.A2(n_866),
.B(n_867),
.Y(n_10715)
);

AOI211x1_ASAP7_75t_L g10716 ( 
.A1(n_10255),
.A2(n_870),
.B(n_868),
.C(n_869),
.Y(n_10716)
);

AOI21x1_ASAP7_75t_L g10717 ( 
.A1(n_10463),
.A2(n_868),
.B(n_869),
.Y(n_10717)
);

OAI21x1_ASAP7_75t_L g10718 ( 
.A1(n_10284),
.A2(n_868),
.B(n_869),
.Y(n_10718)
);

NAND2xp5_ASAP7_75t_SL g10719 ( 
.A(n_10602),
.B(n_870),
.Y(n_10719)
);

NAND2xp5_ASAP7_75t_L g10720 ( 
.A(n_10332),
.B(n_870),
.Y(n_10720)
);

AND2x2_ASAP7_75t_L g10721 ( 
.A(n_10491),
.B(n_871),
.Y(n_10721)
);

NAND2xp5_ASAP7_75t_L g10722 ( 
.A(n_10396),
.B(n_871),
.Y(n_10722)
);

OAI22xp5_ASAP7_75t_L g10723 ( 
.A1(n_10218),
.A2(n_873),
.B1(n_871),
.B2(n_872),
.Y(n_10723)
);

NAND2xp5_ASAP7_75t_L g10724 ( 
.A(n_10429),
.B(n_873),
.Y(n_10724)
);

A2O1A1Ixp33_ASAP7_75t_L g10725 ( 
.A1(n_10215),
.A2(n_876),
.B(n_874),
.C(n_875),
.Y(n_10725)
);

OAI21x1_ASAP7_75t_L g10726 ( 
.A1(n_10341),
.A2(n_874),
.B(n_875),
.Y(n_10726)
);

NAND2xp5_ASAP7_75t_L g10727 ( 
.A(n_10432),
.B(n_874),
.Y(n_10727)
);

OAI21x1_ASAP7_75t_L g10728 ( 
.A1(n_10355),
.A2(n_875),
.B(n_877),
.Y(n_10728)
);

INVx1_ASAP7_75t_L g10729 ( 
.A(n_10439),
.Y(n_10729)
);

AND2x2_ASAP7_75t_L g10730 ( 
.A(n_10623),
.B(n_877),
.Y(n_10730)
);

NAND2xp5_ASAP7_75t_L g10731 ( 
.A(n_10576),
.B(n_879),
.Y(n_10731)
);

AOI221xp5_ASAP7_75t_L g10732 ( 
.A1(n_10503),
.A2(n_881),
.B1(n_879),
.B2(n_880),
.C(n_882),
.Y(n_10732)
);

AOI21xp5_ASAP7_75t_L g10733 ( 
.A1(n_10225),
.A2(n_879),
.B(n_880),
.Y(n_10733)
);

AND2x2_ASAP7_75t_L g10734 ( 
.A(n_10378),
.B(n_10520),
.Y(n_10734)
);

OA21x2_ASAP7_75t_L g10735 ( 
.A1(n_10204),
.A2(n_880),
.B(n_881),
.Y(n_10735)
);

AOI21xp5_ASAP7_75t_L g10736 ( 
.A1(n_10191),
.A2(n_882),
.B(n_883),
.Y(n_10736)
);

NAND2xp5_ASAP7_75t_L g10737 ( 
.A(n_10399),
.B(n_883),
.Y(n_10737)
);

AOI21xp5_ASAP7_75t_L g10738 ( 
.A1(n_10245),
.A2(n_884),
.B(n_885),
.Y(n_10738)
);

O2A1O1Ixp33_ASAP7_75t_SL g10739 ( 
.A1(n_10162),
.A2(n_886),
.B(n_884),
.C(n_885),
.Y(n_10739)
);

AOI21xp5_ASAP7_75t_SL g10740 ( 
.A1(n_10280),
.A2(n_886),
.B(n_887),
.Y(n_10740)
);

OAI21x1_ASAP7_75t_L g10741 ( 
.A1(n_10481),
.A2(n_10303),
.B(n_10185),
.Y(n_10741)
);

AOI21xp5_ASAP7_75t_L g10742 ( 
.A1(n_10300),
.A2(n_887),
.B(n_888),
.Y(n_10742)
);

OAI21x1_ASAP7_75t_L g10743 ( 
.A1(n_10202),
.A2(n_888),
.B(n_889),
.Y(n_10743)
);

BUFx12f_ASAP7_75t_L g10744 ( 
.A(n_10235),
.Y(n_10744)
);

INVx2_ASAP7_75t_SL g10745 ( 
.A(n_10241),
.Y(n_10745)
);

OAI21x1_ASAP7_75t_L g10746 ( 
.A1(n_10171),
.A2(n_10243),
.B(n_10433),
.Y(n_10746)
);

NAND2xp5_ASAP7_75t_L g10747 ( 
.A(n_10384),
.B(n_889),
.Y(n_10747)
);

INVx1_ASAP7_75t_L g10748 ( 
.A(n_10500),
.Y(n_10748)
);

NAND2xp5_ASAP7_75t_L g10749 ( 
.A(n_10452),
.B(n_889),
.Y(n_10749)
);

OAI21x1_ASAP7_75t_L g10750 ( 
.A1(n_10205),
.A2(n_890),
.B(n_891),
.Y(n_10750)
);

NAND3xp33_ASAP7_75t_SL g10751 ( 
.A(n_10361),
.B(n_890),
.C(n_891),
.Y(n_10751)
);

AND2x4_ASAP7_75t_L g10752 ( 
.A(n_10540),
.B(n_890),
.Y(n_10752)
);

OAI21xp5_ASAP7_75t_L g10753 ( 
.A1(n_10152),
.A2(n_891),
.B(n_892),
.Y(n_10753)
);

HB1xp67_ASAP7_75t_L g10754 ( 
.A(n_10151),
.Y(n_10754)
);

AOI21x1_ASAP7_75t_L g10755 ( 
.A1(n_10404),
.A2(n_893),
.B(n_894),
.Y(n_10755)
);

AND2x4_ASAP7_75t_L g10756 ( 
.A(n_10443),
.B(n_893),
.Y(n_10756)
);

AOI21xp5_ASAP7_75t_L g10757 ( 
.A1(n_10382),
.A2(n_895),
.B(n_896),
.Y(n_10757)
);

OAI21x1_ASAP7_75t_L g10758 ( 
.A1(n_10213),
.A2(n_895),
.B(n_896),
.Y(n_10758)
);

AOI21xp5_ASAP7_75t_L g10759 ( 
.A1(n_10281),
.A2(n_895),
.B(n_896),
.Y(n_10759)
);

NAND2xp5_ASAP7_75t_L g10760 ( 
.A(n_10505),
.B(n_897),
.Y(n_10760)
);

INVx5_ASAP7_75t_L g10761 ( 
.A(n_10366),
.Y(n_10761)
);

OAI21x1_ASAP7_75t_L g10762 ( 
.A1(n_10216),
.A2(n_10226),
.B(n_10222),
.Y(n_10762)
);

AO31x2_ASAP7_75t_L g10763 ( 
.A1(n_10376),
.A2(n_899),
.A3(n_897),
.B(n_898),
.Y(n_10763)
);

INVx1_ASAP7_75t_L g10764 ( 
.A(n_10630),
.Y(n_10764)
);

AOI21xp5_ASAP7_75t_L g10765 ( 
.A1(n_10217),
.A2(n_898),
.B(n_900),
.Y(n_10765)
);

NAND2xp5_ASAP7_75t_L g10766 ( 
.A(n_10547),
.B(n_898),
.Y(n_10766)
);

OAI21x1_ASAP7_75t_L g10767 ( 
.A1(n_10261),
.A2(n_900),
.B(n_901),
.Y(n_10767)
);

AOI21xp5_ASAP7_75t_L g10768 ( 
.A1(n_10447),
.A2(n_900),
.B(n_901),
.Y(n_10768)
);

BUFx2_ASAP7_75t_L g10769 ( 
.A(n_10466),
.Y(n_10769)
);

AOI21xp5_ASAP7_75t_L g10770 ( 
.A1(n_10313),
.A2(n_901),
.B(n_902),
.Y(n_10770)
);

BUFx3_ASAP7_75t_L g10771 ( 
.A(n_10428),
.Y(n_10771)
);

INVx1_ASAP7_75t_L g10772 ( 
.A(n_10172),
.Y(n_10772)
);

INVx1_ASAP7_75t_L g10773 ( 
.A(n_10232),
.Y(n_10773)
);

NAND2xp5_ASAP7_75t_SL g10774 ( 
.A(n_10518),
.B(n_902),
.Y(n_10774)
);

OA21x2_ASAP7_75t_L g10775 ( 
.A1(n_10268),
.A2(n_903),
.B(n_904),
.Y(n_10775)
);

BUFx2_ASAP7_75t_L g10776 ( 
.A(n_10158),
.Y(n_10776)
);

A2O1A1Ixp33_ASAP7_75t_L g10777 ( 
.A1(n_10329),
.A2(n_905),
.B(n_903),
.C(n_904),
.Y(n_10777)
);

OAI22xp5_ASAP7_75t_L g10778 ( 
.A1(n_10310),
.A2(n_906),
.B1(n_903),
.B2(n_905),
.Y(n_10778)
);

OAI21x1_ASAP7_75t_L g10779 ( 
.A1(n_10270),
.A2(n_906),
.B(n_907),
.Y(n_10779)
);

OAI21xp5_ASAP7_75t_L g10780 ( 
.A1(n_10173),
.A2(n_907),
.B(n_908),
.Y(n_10780)
);

INVx3_ASAP7_75t_SL g10781 ( 
.A(n_10285),
.Y(n_10781)
);

OAI21xp5_ASAP7_75t_L g10782 ( 
.A1(n_10438),
.A2(n_10347),
.B(n_10295),
.Y(n_10782)
);

OA21x2_ASAP7_75t_L g10783 ( 
.A1(n_10308),
.A2(n_907),
.B(n_908),
.Y(n_10783)
);

NOR2xp33_ASAP7_75t_R g10784 ( 
.A(n_10416),
.B(n_909),
.Y(n_10784)
);

BUFx6f_ASAP7_75t_L g10785 ( 
.A(n_10251),
.Y(n_10785)
);

AO31x2_ASAP7_75t_L g10786 ( 
.A1(n_10353),
.A2(n_911),
.A3(n_909),
.B(n_910),
.Y(n_10786)
);

BUFx2_ASAP7_75t_L g10787 ( 
.A(n_10374),
.Y(n_10787)
);

NAND2xp5_ASAP7_75t_L g10788 ( 
.A(n_10178),
.B(n_909),
.Y(n_10788)
);

NAND2xp5_ASAP7_75t_L g10789 ( 
.A(n_10181),
.B(n_910),
.Y(n_10789)
);

INVx1_ASAP7_75t_L g10790 ( 
.A(n_10233),
.Y(n_10790)
);

OAI21x1_ASAP7_75t_L g10791 ( 
.A1(n_10309),
.A2(n_910),
.B(n_911),
.Y(n_10791)
);

OAI21x1_ASAP7_75t_L g10792 ( 
.A1(n_10311),
.A2(n_912),
.B(n_913),
.Y(n_10792)
);

NAND2xp5_ASAP7_75t_L g10793 ( 
.A(n_10161),
.B(n_912),
.Y(n_10793)
);

INVx1_ASAP7_75t_L g10794 ( 
.A(n_10250),
.Y(n_10794)
);

INVx1_ASAP7_75t_L g10795 ( 
.A(n_10334),
.Y(n_10795)
);

OA21x2_ASAP7_75t_L g10796 ( 
.A1(n_10315),
.A2(n_913),
.B(n_914),
.Y(n_10796)
);

INVx1_ASAP7_75t_L g10797 ( 
.A(n_10364),
.Y(n_10797)
);

NAND2xp5_ASAP7_75t_L g10798 ( 
.A(n_10166),
.B(n_914),
.Y(n_10798)
);

HB1xp67_ASAP7_75t_L g10799 ( 
.A(n_10180),
.Y(n_10799)
);

NOR2xp33_ASAP7_75t_L g10800 ( 
.A(n_10292),
.B(n_915),
.Y(n_10800)
);

NAND2xp5_ASAP7_75t_L g10801 ( 
.A(n_10367),
.B(n_915),
.Y(n_10801)
);

OAI21xp33_ASAP7_75t_L g10802 ( 
.A1(n_10164),
.A2(n_916),
.B(n_917),
.Y(n_10802)
);

OAI21x1_ASAP7_75t_L g10803 ( 
.A1(n_10209),
.A2(n_916),
.B(n_917),
.Y(n_10803)
);

OAI21x1_ASAP7_75t_L g10804 ( 
.A1(n_10190),
.A2(n_916),
.B(n_918),
.Y(n_10804)
);

NAND2xp5_ASAP7_75t_L g10805 ( 
.A(n_10345),
.B(n_918),
.Y(n_10805)
);

A2O1A1Ixp33_ASAP7_75t_L g10806 ( 
.A1(n_10192),
.A2(n_921),
.B(n_919),
.C(n_920),
.Y(n_10806)
);

NAND2xp5_ASAP7_75t_SL g10807 ( 
.A(n_10518),
.B(n_919),
.Y(n_10807)
);

NAND2xp5_ASAP7_75t_L g10808 ( 
.A(n_10437),
.B(n_919),
.Y(n_10808)
);

NOR4xp25_ASAP7_75t_L g10809 ( 
.A(n_10627),
.B(n_922),
.C(n_920),
.D(n_921),
.Y(n_10809)
);

A2O1A1Ixp33_ASAP7_75t_L g10810 ( 
.A1(n_10624),
.A2(n_923),
.B(n_920),
.C(n_922),
.Y(n_10810)
);

INVx4_ASAP7_75t_L g10811 ( 
.A(n_10492),
.Y(n_10811)
);

AOI21xp5_ASAP7_75t_L g10812 ( 
.A1(n_10187),
.A2(n_10351),
.B(n_10269),
.Y(n_10812)
);

AO31x2_ASAP7_75t_L g10813 ( 
.A1(n_10421),
.A2(n_925),
.A3(n_923),
.B(n_924),
.Y(n_10813)
);

AND2x2_ASAP7_75t_L g10814 ( 
.A(n_10501),
.B(n_923),
.Y(n_10814)
);

AOI21x1_ASAP7_75t_L g10815 ( 
.A1(n_10472),
.A2(n_924),
.B(n_925),
.Y(n_10815)
);

AOI21xp5_ASAP7_75t_L g10816 ( 
.A1(n_10223),
.A2(n_926),
.B(n_927),
.Y(n_10816)
);

NOR2xp33_ASAP7_75t_SL g10817 ( 
.A(n_10392),
.B(n_926),
.Y(n_10817)
);

NAND2xp5_ASAP7_75t_L g10818 ( 
.A(n_10154),
.B(n_926),
.Y(n_10818)
);

OAI21x1_ASAP7_75t_L g10819 ( 
.A1(n_10193),
.A2(n_927),
.B(n_928),
.Y(n_10819)
);

OAI21x1_ASAP7_75t_SL g10820 ( 
.A1(n_10509),
.A2(n_928),
.B(n_929),
.Y(n_10820)
);

OR2x6_ASAP7_75t_L g10821 ( 
.A(n_10188),
.B(n_929),
.Y(n_10821)
);

NAND2xp5_ASAP7_75t_L g10822 ( 
.A(n_10176),
.B(n_930),
.Y(n_10822)
);

NAND2xp5_ASAP7_75t_L g10823 ( 
.A(n_10163),
.B(n_930),
.Y(n_10823)
);

OAI21x1_ASAP7_75t_L g10824 ( 
.A1(n_10617),
.A2(n_930),
.B(n_931),
.Y(n_10824)
);

NOR4xp25_ASAP7_75t_L g10825 ( 
.A(n_10554),
.B(n_933),
.C(n_931),
.D(n_932),
.Y(n_10825)
);

INVx2_ASAP7_75t_SL g10826 ( 
.A(n_10487),
.Y(n_10826)
);

OAI21x1_ASAP7_75t_L g10827 ( 
.A1(n_10201),
.A2(n_10372),
.B(n_10363),
.Y(n_10827)
);

AOI21xp5_ASAP7_75t_L g10828 ( 
.A1(n_10244),
.A2(n_931),
.B(n_932),
.Y(n_10828)
);

OR2x6_ASAP7_75t_L g10829 ( 
.A(n_10188),
.B(n_933),
.Y(n_10829)
);

AOI21xp5_ASAP7_75t_L g10830 ( 
.A1(n_10306),
.A2(n_933),
.B(n_934),
.Y(n_10830)
);

BUFx12f_ASAP7_75t_L g10831 ( 
.A(n_10512),
.Y(n_10831)
);

NAND2xp5_ASAP7_75t_L g10832 ( 
.A(n_10388),
.B(n_934),
.Y(n_10832)
);

OAI21xp5_ASAP7_75t_L g10833 ( 
.A1(n_10297),
.A2(n_10290),
.B(n_10397),
.Y(n_10833)
);

AOI21xp5_ASAP7_75t_L g10834 ( 
.A1(n_10417),
.A2(n_934),
.B(n_935),
.Y(n_10834)
);

OAI21xp5_ASAP7_75t_L g10835 ( 
.A1(n_10278),
.A2(n_935),
.B(n_936),
.Y(n_10835)
);

OR2x2_ASAP7_75t_L g10836 ( 
.A(n_10419),
.B(n_935),
.Y(n_10836)
);

OAI22xp5_ASAP7_75t_L g10837 ( 
.A1(n_10379),
.A2(n_938),
.B1(n_936),
.B2(n_937),
.Y(n_10837)
);

AOI21xp5_ASAP7_75t_L g10838 ( 
.A1(n_10381),
.A2(n_936),
.B(n_937),
.Y(n_10838)
);

NAND2xp5_ASAP7_75t_L g10839 ( 
.A(n_10566),
.B(n_937),
.Y(n_10839)
);

NAND3xp33_ASAP7_75t_L g10840 ( 
.A(n_10453),
.B(n_10586),
.C(n_10638),
.Y(n_10840)
);

AND2x2_ASAP7_75t_L g10841 ( 
.A(n_10647),
.B(n_938),
.Y(n_10841)
);

NAND3x1_ASAP7_75t_L g10842 ( 
.A(n_10616),
.B(n_938),
.C(n_940),
.Y(n_10842)
);

OR2x6_ASAP7_75t_L g10843 ( 
.A(n_10340),
.B(n_940),
.Y(n_10843)
);

NAND2xp5_ASAP7_75t_L g10844 ( 
.A(n_10406),
.B(n_940),
.Y(n_10844)
);

INVx1_ASAP7_75t_L g10845 ( 
.A(n_10370),
.Y(n_10845)
);

NAND2xp5_ASAP7_75t_L g10846 ( 
.A(n_10469),
.B(n_941),
.Y(n_10846)
);

BUFx3_ASAP7_75t_L g10847 ( 
.A(n_10596),
.Y(n_10847)
);

A2O1A1Ixp33_ASAP7_75t_L g10848 ( 
.A1(n_10368),
.A2(n_943),
.B(n_941),
.C(n_942),
.Y(n_10848)
);

AOI21xp33_ASAP7_75t_L g10849 ( 
.A1(n_10159),
.A2(n_941),
.B(n_942),
.Y(n_10849)
);

INVx2_ASAP7_75t_L g10850 ( 
.A(n_10401),
.Y(n_10850)
);

INVx1_ASAP7_75t_SL g10851 ( 
.A(n_10462),
.Y(n_10851)
);

INVx1_ASAP7_75t_L g10852 ( 
.A(n_10502),
.Y(n_10852)
);

AOI221xp5_ASAP7_75t_SL g10853 ( 
.A1(n_10603),
.A2(n_944),
.B1(n_942),
.B2(n_943),
.C(n_945),
.Y(n_10853)
);

NAND3xp33_ASAP7_75t_L g10854 ( 
.A(n_10350),
.B(n_943),
.C(n_944),
.Y(n_10854)
);

AO21x2_ASAP7_75t_L g10855 ( 
.A1(n_10488),
.A2(n_944),
.B(n_945),
.Y(n_10855)
);

AND2x4_ASAP7_75t_L g10856 ( 
.A(n_10583),
.B(n_10613),
.Y(n_10856)
);

AOI21xp5_ASAP7_75t_L g10857 ( 
.A1(n_10385),
.A2(n_945),
.B(n_946),
.Y(n_10857)
);

INVx2_ASAP7_75t_L g10858 ( 
.A(n_10442),
.Y(n_10858)
);

AOI21xp5_ASAP7_75t_L g10859 ( 
.A1(n_10291),
.A2(n_946),
.B(n_947),
.Y(n_10859)
);

AOI21xp5_ASAP7_75t_L g10860 ( 
.A1(n_10248),
.A2(n_946),
.B(n_947),
.Y(n_10860)
);

INVx2_ASAP7_75t_L g10861 ( 
.A(n_10461),
.Y(n_10861)
);

AOI21xp5_ASAP7_75t_L g10862 ( 
.A1(n_10465),
.A2(n_948),
.B(n_949),
.Y(n_10862)
);

NAND3xp33_ASAP7_75t_L g10863 ( 
.A(n_10511),
.B(n_948),
.C(n_950),
.Y(n_10863)
);

NAND2xp5_ASAP7_75t_SL g10864 ( 
.A(n_10288),
.B(n_10383),
.Y(n_10864)
);

OAI21x1_ASAP7_75t_L g10865 ( 
.A1(n_10373),
.A2(n_948),
.B(n_950),
.Y(n_10865)
);

OAI21x1_ASAP7_75t_L g10866 ( 
.A1(n_10380),
.A2(n_950),
.B(n_951),
.Y(n_10866)
);

OAI21xp5_ASAP7_75t_L g10867 ( 
.A1(n_10569),
.A2(n_951),
.B(n_952),
.Y(n_10867)
);

A2O1A1Ixp33_ASAP7_75t_L g10868 ( 
.A1(n_10398),
.A2(n_953),
.B(n_951),
.C(n_952),
.Y(n_10868)
);

OAI21x1_ASAP7_75t_L g10869 ( 
.A1(n_10393),
.A2(n_953),
.B(n_954),
.Y(n_10869)
);

INVx1_ASAP7_75t_L g10870 ( 
.A(n_10515),
.Y(n_10870)
);

AOI221x1_ASAP7_75t_L g10871 ( 
.A1(n_10495),
.A2(n_955),
.B1(n_953),
.B2(n_954),
.C(n_956),
.Y(n_10871)
);

AO31x2_ASAP7_75t_L g10872 ( 
.A1(n_10536),
.A2(n_956),
.A3(n_954),
.B(n_955),
.Y(n_10872)
);

AOI21xp5_ASAP7_75t_L g10873 ( 
.A1(n_10153),
.A2(n_955),
.B(n_956),
.Y(n_10873)
);

NOR2xp33_ASAP7_75t_L g10874 ( 
.A(n_10629),
.B(n_957),
.Y(n_10874)
);

OAI21x1_ASAP7_75t_L g10875 ( 
.A1(n_10307),
.A2(n_957),
.B(n_958),
.Y(n_10875)
);

AOI21xp5_ASAP7_75t_L g10876 ( 
.A1(n_10208),
.A2(n_957),
.B(n_958),
.Y(n_10876)
);

INVx2_ASAP7_75t_L g10877 ( 
.A(n_10478),
.Y(n_10877)
);

INVx1_ASAP7_75t_L g10878 ( 
.A(n_10537),
.Y(n_10878)
);

A2O1A1Ixp33_ASAP7_75t_L g10879 ( 
.A1(n_10620),
.A2(n_960),
.B(n_958),
.C(n_959),
.Y(n_10879)
);

NAND2xp5_ASAP7_75t_L g10880 ( 
.A(n_10237),
.B(n_959),
.Y(n_10880)
);

NAND2xp5_ASAP7_75t_L g10881 ( 
.A(n_10377),
.B(n_960),
.Y(n_10881)
);

AOI21xp5_ASAP7_75t_L g10882 ( 
.A1(n_10418),
.A2(n_960),
.B(n_961),
.Y(n_10882)
);

OAI21x1_ASAP7_75t_L g10883 ( 
.A1(n_10314),
.A2(n_961),
.B(n_962),
.Y(n_10883)
);

AOI221xp5_ASAP7_75t_SL g10884 ( 
.A1(n_10282),
.A2(n_10395),
.B1(n_10327),
.B2(n_10454),
.C(n_10287),
.Y(n_10884)
);

INVx2_ASAP7_75t_L g10885 ( 
.A(n_10484),
.Y(n_10885)
);

OAI21xp5_ASAP7_75t_L g10886 ( 
.A1(n_10343),
.A2(n_962),
.B(n_963),
.Y(n_10886)
);

INVx3_ASAP7_75t_L g10887 ( 
.A(n_10360),
.Y(n_10887)
);

INVx2_ASAP7_75t_L g10888 ( 
.A(n_10508),
.Y(n_10888)
);

OAI22xp5_ASAP7_75t_L g10889 ( 
.A1(n_10340),
.A2(n_965),
.B1(n_963),
.B2(n_964),
.Y(n_10889)
);

NOR2xp67_ASAP7_75t_SL g10890 ( 
.A(n_10517),
.B(n_963),
.Y(n_10890)
);

AOI211x1_ASAP7_75t_L g10891 ( 
.A1(n_10323),
.A2(n_966),
.B(n_964),
.C(n_965),
.Y(n_10891)
);

NAND2xp5_ASAP7_75t_L g10892 ( 
.A(n_10498),
.B(n_10507),
.Y(n_10892)
);

BUFx6f_ASAP7_75t_L g10893 ( 
.A(n_10251),
.Y(n_10893)
);

NOR4xp25_ASAP7_75t_L g10894 ( 
.A(n_10595),
.B(n_966),
.C(n_964),
.D(n_965),
.Y(n_10894)
);

NOR2xp33_ASAP7_75t_L g10895 ( 
.A(n_10256),
.B(n_966),
.Y(n_10895)
);

AND2x2_ASAP7_75t_L g10896 ( 
.A(n_10446),
.B(n_967),
.Y(n_10896)
);

NOR2xp33_ASAP7_75t_SL g10897 ( 
.A(n_10544),
.B(n_967),
.Y(n_10897)
);

NAND2xp5_ASAP7_75t_L g10898 ( 
.A(n_10530),
.B(n_967),
.Y(n_10898)
);

OAI21x1_ASAP7_75t_L g10899 ( 
.A1(n_10316),
.A2(n_968),
.B(n_969),
.Y(n_10899)
);

BUFx3_ASAP7_75t_L g10900 ( 
.A(n_10256),
.Y(n_10900)
);

NAND2xp5_ASAP7_75t_L g10901 ( 
.A(n_10556),
.B(n_968),
.Y(n_10901)
);

AOI21xp5_ASAP7_75t_L g10902 ( 
.A1(n_10405),
.A2(n_968),
.B(n_969),
.Y(n_10902)
);

OR2x6_ASAP7_75t_L g10903 ( 
.A(n_10455),
.B(n_969),
.Y(n_10903)
);

INVx6_ASAP7_75t_L g10904 ( 
.A(n_10324),
.Y(n_10904)
);

OAI22xp5_ASAP7_75t_L g10905 ( 
.A1(n_10330),
.A2(n_973),
.B1(n_970),
.B2(n_971),
.Y(n_10905)
);

INVxp33_ASAP7_75t_L g10906 ( 
.A(n_10267),
.Y(n_10906)
);

AOI221x1_ASAP7_75t_L g10907 ( 
.A1(n_10390),
.A2(n_973),
.B1(n_970),
.B2(n_971),
.C(n_974),
.Y(n_10907)
);

OAI21x1_ASAP7_75t_L g10908 ( 
.A1(n_10317),
.A2(n_970),
.B(n_973),
.Y(n_10908)
);

O2A1O1Ixp5_ASAP7_75t_L g10909 ( 
.A1(n_10609),
.A2(n_976),
.B(n_974),
.C(n_975),
.Y(n_10909)
);

AOI21x1_ASAP7_75t_L g10910 ( 
.A1(n_10344),
.A2(n_974),
.B(n_975),
.Y(n_10910)
);

OAI21x1_ASAP7_75t_L g10911 ( 
.A1(n_10320),
.A2(n_975),
.B(n_976),
.Y(n_10911)
);

AOI21xp5_ASAP7_75t_L g10912 ( 
.A1(n_10253),
.A2(n_10312),
.B(n_10420),
.Y(n_10912)
);

INVx1_ASAP7_75t_L g10913 ( 
.A(n_10570),
.Y(n_10913)
);

AOI221x1_ASAP7_75t_L g10914 ( 
.A1(n_10430),
.A2(n_10558),
.B1(n_10563),
.B2(n_10562),
.C(n_10557),
.Y(n_10914)
);

NAND2xp5_ASAP7_75t_L g10915 ( 
.A(n_10468),
.B(n_976),
.Y(n_10915)
);

BUFx6f_ASAP7_75t_L g10916 ( 
.A(n_10387),
.Y(n_10916)
);

INVx3_ASAP7_75t_L g10917 ( 
.A(n_10482),
.Y(n_10917)
);

A2O1A1Ixp33_ASAP7_75t_L g10918 ( 
.A1(n_10622),
.A2(n_979),
.B(n_977),
.C(n_978),
.Y(n_10918)
);

AOI21x1_ASAP7_75t_L g10919 ( 
.A1(n_10597),
.A2(n_977),
.B(n_978),
.Y(n_10919)
);

OA21x2_ASAP7_75t_L g10920 ( 
.A1(n_10606),
.A2(n_977),
.B(n_978),
.Y(n_10920)
);

OA21x2_ASAP7_75t_L g10921 ( 
.A1(n_10633),
.A2(n_979),
.B(n_980),
.Y(n_10921)
);

AOI21x1_ASAP7_75t_L g10922 ( 
.A1(n_10296),
.A2(n_979),
.B(n_980),
.Y(n_10922)
);

BUFx8_ASAP7_75t_L g10923 ( 
.A(n_10239),
.Y(n_10923)
);

NAND3xp33_ASAP7_75t_L g10924 ( 
.A(n_10514),
.B(n_981),
.C(n_982),
.Y(n_10924)
);

AO32x2_ASAP7_75t_L g10925 ( 
.A1(n_10409),
.A2(n_983),
.A3(n_981),
.B1(n_982),
.B2(n_984),
.Y(n_10925)
);

AOI21xp5_ASAP7_75t_L g10926 ( 
.A1(n_10499),
.A2(n_982),
.B(n_983),
.Y(n_10926)
);

OAI21xp5_ASAP7_75t_SL g10927 ( 
.A1(n_10445),
.A2(n_983),
.B(n_984),
.Y(n_10927)
);

AOI221xp5_ASAP7_75t_L g10928 ( 
.A1(n_10170),
.A2(n_986),
.B1(n_984),
.B2(n_985),
.C(n_987),
.Y(n_10928)
);

CKINVDCx20_ASAP7_75t_R g10929 ( 
.A(n_10459),
.Y(n_10929)
);

OAI21xp5_ASAP7_75t_L g10930 ( 
.A1(n_10265),
.A2(n_10489),
.B(n_10471),
.Y(n_10930)
);

CKINVDCx11_ASAP7_75t_R g10931 ( 
.A(n_10545),
.Y(n_10931)
);

NAND2xp5_ASAP7_75t_L g10932 ( 
.A(n_10477),
.B(n_985),
.Y(n_10932)
);

OAI21x1_ASAP7_75t_L g10933 ( 
.A1(n_10337),
.A2(n_985),
.B(n_986),
.Y(n_10933)
);

AOI21xp5_ASAP7_75t_L g10934 ( 
.A1(n_10523),
.A2(n_986),
.B(n_987),
.Y(n_10934)
);

AOI21xp5_ASAP7_75t_L g10935 ( 
.A1(n_10474),
.A2(n_10568),
.B(n_10476),
.Y(n_10935)
);

A2O1A1Ixp33_ASAP7_75t_L g10936 ( 
.A1(n_10365),
.A2(n_990),
.B(n_987),
.C(n_989),
.Y(n_10936)
);

AOI21xp5_ASAP7_75t_L g10937 ( 
.A1(n_10574),
.A2(n_989),
.B(n_990),
.Y(n_10937)
);

INVx1_ASAP7_75t_L g10938 ( 
.A(n_10642),
.Y(n_10938)
);

OAI21x1_ASAP7_75t_L g10939 ( 
.A1(n_10339),
.A2(n_989),
.B(n_990),
.Y(n_10939)
);

AND2x4_ASAP7_75t_L g10940 ( 
.A(n_10542),
.B(n_991),
.Y(n_10940)
);

BUFx6f_ASAP7_75t_L g10941 ( 
.A(n_10444),
.Y(n_10941)
);

HB1xp67_ASAP7_75t_L g10942 ( 
.A(n_10349),
.Y(n_10942)
);

NAND2xp5_ASAP7_75t_L g10943 ( 
.A(n_10486),
.B(n_991),
.Y(n_10943)
);

O2A1O1Ixp5_ASAP7_75t_L g10944 ( 
.A1(n_10483),
.A2(n_993),
.B(n_991),
.C(n_992),
.Y(n_10944)
);

AOI21xp5_ASAP7_75t_L g10945 ( 
.A1(n_10592),
.A2(n_992),
.B(n_993),
.Y(n_10945)
);

AOI22xp33_ASAP7_75t_L g10946 ( 
.A1(n_10254),
.A2(n_994),
.B1(n_992),
.B2(n_993),
.Y(n_10946)
);

AOI21xp5_ASAP7_75t_L g10947 ( 
.A1(n_10467),
.A2(n_994),
.B(n_995),
.Y(n_10947)
);

BUFx3_ASAP7_75t_L g10948 ( 
.A(n_10436),
.Y(n_10948)
);

INVx2_ASAP7_75t_L g10949 ( 
.A(n_10541),
.Y(n_10949)
);

OAI21x1_ASAP7_75t_L g10950 ( 
.A1(n_10342),
.A2(n_995),
.B(n_996),
.Y(n_10950)
);

AOI21xp5_ASAP7_75t_L g10951 ( 
.A1(n_10375),
.A2(n_996),
.B(n_997),
.Y(n_10951)
);

OAI21x1_ASAP7_75t_L g10952 ( 
.A1(n_10553),
.A2(n_996),
.B(n_997),
.Y(n_10952)
);

AND2x6_ASAP7_75t_L g10953 ( 
.A(n_10203),
.B(n_10578),
.Y(n_10953)
);

INVx1_ASAP7_75t_L g10954 ( 
.A(n_10555),
.Y(n_10954)
);

NOR2xp33_ASAP7_75t_SL g10955 ( 
.A(n_10579),
.B(n_997),
.Y(n_10955)
);

NAND2xp5_ASAP7_75t_L g10956 ( 
.A(n_10564),
.B(n_998),
.Y(n_10956)
);

AO32x2_ASAP7_75t_L g10957 ( 
.A1(n_10400),
.A2(n_1000),
.A3(n_998),
.B1(n_999),
.B2(n_1001),
.Y(n_10957)
);

NAND2xp5_ASAP7_75t_L g10958 ( 
.A(n_10571),
.B(n_999),
.Y(n_10958)
);

A2O1A1Ixp33_ASAP7_75t_L g10959 ( 
.A1(n_10626),
.A2(n_1001),
.B(n_999),
.C(n_1000),
.Y(n_10959)
);

NOR2xp33_ASAP7_75t_L g10960 ( 
.A(n_10516),
.B(n_1000),
.Y(n_10960)
);

OAI21x1_ASAP7_75t_L g10961 ( 
.A1(n_10230),
.A2(n_1001),
.B(n_1002),
.Y(n_10961)
);

CKINVDCx5p33_ASAP7_75t_R g10962 ( 
.A(n_10646),
.Y(n_10962)
);

AO21x1_ASAP7_75t_L g10963 ( 
.A1(n_10391),
.A2(n_1002),
.B(n_1003),
.Y(n_10963)
);

AOI22xp5_ASAP7_75t_L g10964 ( 
.A1(n_10283),
.A2(n_1005),
.B1(n_1003),
.B2(n_1004),
.Y(n_10964)
);

AOI21xp5_ASAP7_75t_L g10965 ( 
.A1(n_10427),
.A2(n_10434),
.B(n_10572),
.Y(n_10965)
);

OAI22xp33_ASAP7_75t_L g10966 ( 
.A1(n_10575),
.A2(n_10635),
.B1(n_10435),
.B2(n_10455),
.Y(n_10966)
);

A2O1A1Ixp33_ASAP7_75t_L g10967 ( 
.A1(n_10632),
.A2(n_1005),
.B(n_1003),
.C(n_1004),
.Y(n_10967)
);

BUFx6f_ASAP7_75t_L g10968 ( 
.A(n_10369),
.Y(n_10968)
);

NOR2x1_ASAP7_75t_L g10969 ( 
.A(n_10577),
.B(n_1004),
.Y(n_10969)
);

OAI21xp5_ASAP7_75t_L g10970 ( 
.A1(n_10567),
.A2(n_1005),
.B(n_1006),
.Y(n_10970)
);

OAI22x1_ASAP7_75t_L g10971 ( 
.A1(n_10195),
.A2(n_1008),
.B1(n_1006),
.B2(n_1007),
.Y(n_10971)
);

AOI22xp33_ASAP7_75t_L g10972 ( 
.A1(n_10621),
.A2(n_1008),
.B1(n_1006),
.B2(n_1007),
.Y(n_10972)
);

AO31x2_ASAP7_75t_L g10973 ( 
.A1(n_10513),
.A2(n_1009),
.A3(n_1007),
.B(n_1008),
.Y(n_10973)
);

INVx2_ASAP7_75t_L g10974 ( 
.A(n_10589),
.Y(n_10974)
);

AND2x4_ASAP7_75t_L g10975 ( 
.A(n_10599),
.B(n_1009),
.Y(n_10975)
);

AND2x4_ASAP7_75t_L g10976 ( 
.A(n_10619),
.B(n_1010),
.Y(n_10976)
);

AOI221x1_ASAP7_75t_L g10977 ( 
.A1(n_10580),
.A2(n_1012),
.B1(n_1010),
.B2(n_1011),
.C(n_1013),
.Y(n_10977)
);

INVx1_ASAP7_75t_L g10978 ( 
.A(n_10644),
.Y(n_10978)
);

OAI21x1_ASAP7_75t_L g10979 ( 
.A1(n_10247),
.A2(n_10274),
.B(n_10272),
.Y(n_10979)
);

INVx2_ASAP7_75t_SL g10980 ( 
.A(n_10328),
.Y(n_10980)
);

A2O1A1Ixp33_ASAP7_75t_L g10981 ( 
.A1(n_10584),
.A2(n_1012),
.B(n_1010),
.C(n_1011),
.Y(n_10981)
);

AND2x4_ASAP7_75t_L g10982 ( 
.A(n_10550),
.B(n_1012),
.Y(n_10982)
);

AOI21xp5_ASAP7_75t_L g10983 ( 
.A1(n_10561),
.A2(n_1013),
.B(n_1014),
.Y(n_10983)
);

AND2x2_ASAP7_75t_L g10984 ( 
.A(n_10356),
.B(n_1014),
.Y(n_10984)
);

HB1xp67_ASAP7_75t_L g10985 ( 
.A(n_10229),
.Y(n_10985)
);

NOR4xp25_ASAP7_75t_L g10986 ( 
.A(n_10628),
.B(n_1016),
.C(n_1014),
.D(n_1015),
.Y(n_10986)
);

AND2x4_ASAP7_75t_L g10987 ( 
.A(n_10283),
.B(n_1015),
.Y(n_10987)
);

OAI21x1_ASAP7_75t_L g10988 ( 
.A1(n_10451),
.A2(n_1015),
.B(n_1016),
.Y(n_10988)
);

AND2x2_ASAP7_75t_L g10989 ( 
.A(n_10559),
.B(n_1016),
.Y(n_10989)
);

INVx1_ASAP7_75t_L g10990 ( 
.A(n_10524),
.Y(n_10990)
);

AND2x2_ASAP7_75t_L g10991 ( 
.A(n_10590),
.B(n_1017),
.Y(n_10991)
);

NAND2xp5_ASAP7_75t_SL g10992 ( 
.A(n_10318),
.B(n_10412),
.Y(n_10992)
);

OAI21xp5_ASAP7_75t_L g10993 ( 
.A1(n_10386),
.A2(n_1017),
.B(n_1018),
.Y(n_10993)
);

AOI211x1_ASAP7_75t_L g10994 ( 
.A1(n_10631),
.A2(n_1020),
.B(n_1018),
.C(n_1019),
.Y(n_10994)
);

NAND2xp5_ASAP7_75t_L g10995 ( 
.A(n_10581),
.B(n_1019),
.Y(n_10995)
);

AOI21xp33_ASAP7_75t_L g10996 ( 
.A1(n_10403),
.A2(n_1020),
.B(n_1021),
.Y(n_10996)
);

AO21x1_ASAP7_75t_L g10997 ( 
.A1(n_10634),
.A2(n_10585),
.B(n_10389),
.Y(n_10997)
);

NAND2xp5_ASAP7_75t_SL g10998 ( 
.A(n_10639),
.B(n_1021),
.Y(n_10998)
);

OAI21xp5_ASAP7_75t_L g10999 ( 
.A1(n_10394),
.A2(n_1021),
.B(n_1022),
.Y(n_10999)
);

OAI21xp5_ASAP7_75t_L g11000 ( 
.A1(n_10526),
.A2(n_1022),
.B(n_1023),
.Y(n_11000)
);

BUFx2_ASAP7_75t_L g11001 ( 
.A(n_10413),
.Y(n_11001)
);

AO31x2_ASAP7_75t_L g11002 ( 
.A1(n_10346),
.A2(n_1024),
.A3(n_1022),
.B(n_1023),
.Y(n_11002)
);

INVx1_ASAP7_75t_L g11003 ( 
.A(n_10524),
.Y(n_11003)
);

NOR2x1_ASAP7_75t_L g11004 ( 
.A(n_10490),
.B(n_1023),
.Y(n_11004)
);

NAND2xp5_ASAP7_75t_L g11005 ( 
.A(n_10526),
.B(n_1024),
.Y(n_11005)
);

OAI22xp33_ASAP7_75t_L g11006 ( 
.A1(n_10640),
.A2(n_1026),
.B1(n_1024),
.B2(n_1025),
.Y(n_11006)
);

AO31x2_ASAP7_75t_L g11007 ( 
.A1(n_10348),
.A2(n_1027),
.A3(n_1025),
.B(n_1026),
.Y(n_11007)
);

AOI211x1_ASAP7_75t_L g11008 ( 
.A1(n_10641),
.A2(n_1028),
.B(n_1025),
.C(n_1027),
.Y(n_11008)
);

NAND2xp5_ASAP7_75t_L g11009 ( 
.A(n_10526),
.B(n_1028),
.Y(n_11009)
);

NAND2xp5_ASAP7_75t_L g11010 ( 
.A(n_10371),
.B(n_1028),
.Y(n_11010)
);

BUFx2_ASAP7_75t_L g11011 ( 
.A(n_10496),
.Y(n_11011)
);

AOI221x1_ASAP7_75t_L g11012 ( 
.A1(n_10464),
.A2(n_1031),
.B1(n_1029),
.B2(n_1030),
.C(n_1032),
.Y(n_11012)
);

INVxp67_ASAP7_75t_L g11013 ( 
.A(n_10615),
.Y(n_11013)
);

OR2x6_ASAP7_75t_L g11014 ( 
.A(n_10643),
.B(n_1029),
.Y(n_11014)
);

BUFx3_ASAP7_75t_L g11015 ( 
.A(n_10175),
.Y(n_11015)
);

NAND2xp5_ASAP7_75t_L g11016 ( 
.A(n_10598),
.B(n_1030),
.Y(n_11016)
);

HB1xp67_ASAP7_75t_L g11017 ( 
.A(n_10229),
.Y(n_11017)
);

INVx5_ASAP7_75t_L g11018 ( 
.A(n_10497),
.Y(n_11018)
);

OAI21xp5_ASAP7_75t_L g11019 ( 
.A1(n_10301),
.A2(n_1030),
.B(n_1033),
.Y(n_11019)
);

AOI21xp5_ASAP7_75t_L g11020 ( 
.A1(n_10565),
.A2(n_1033),
.B(n_1034),
.Y(n_11020)
);

OAI21xp5_ASAP7_75t_L g11021 ( 
.A1(n_10302),
.A2(n_1034),
.B(n_1035),
.Y(n_11021)
);

O2A1O1Ixp33_ASAP7_75t_SL g11022 ( 
.A1(n_10414),
.A2(n_1037),
.B(n_1035),
.C(n_1036),
.Y(n_11022)
);

INVx1_ASAP7_75t_SL g11023 ( 
.A(n_10625),
.Y(n_11023)
);

NAND2xp5_ASAP7_75t_SL g11024 ( 
.A(n_10604),
.B(n_1035),
.Y(n_11024)
);

NAND2xp5_ASAP7_75t_L g11025 ( 
.A(n_10610),
.B(n_1036),
.Y(n_11025)
);

OAI21x1_ASAP7_75t_L g11026 ( 
.A1(n_10198),
.A2(n_1036),
.B(n_1037),
.Y(n_11026)
);

NAND2xp5_ASAP7_75t_L g11027 ( 
.A(n_10611),
.B(n_1038),
.Y(n_11027)
);

NAND2x1p5_ASAP7_75t_L g11028 ( 
.A(n_10470),
.B(n_1038),
.Y(n_11028)
);

NAND2xp5_ASAP7_75t_SL g11029 ( 
.A(n_10425),
.B(n_1039),
.Y(n_11029)
);

AOI21xp5_ASAP7_75t_L g11030 ( 
.A1(n_10600),
.A2(n_1039),
.B(n_1040),
.Y(n_11030)
);

INVx3_ASAP7_75t_L g11031 ( 
.A(n_10497),
.Y(n_11031)
);

INVx1_ASAP7_75t_L g11032 ( 
.A(n_10582),
.Y(n_11032)
);

OAI21xp5_ASAP7_75t_L g11033 ( 
.A1(n_10304),
.A2(n_1039),
.B(n_1040),
.Y(n_11033)
);

A2O1A1Ixp33_ASAP7_75t_L g11034 ( 
.A1(n_10196),
.A2(n_1042),
.B(n_1040),
.C(n_1041),
.Y(n_11034)
);

BUFx6f_ASAP7_75t_L g11035 ( 
.A(n_10497),
.Y(n_11035)
);

NAND3xp33_ASAP7_75t_L g11036 ( 
.A(n_10354),
.B(n_1041),
.C(n_1042),
.Y(n_11036)
);

NAND2xp5_ASAP7_75t_L g11037 ( 
.A(n_10426),
.B(n_1041),
.Y(n_11037)
);

INVx1_ASAP7_75t_L g11038 ( 
.A(n_10582),
.Y(n_11038)
);

AOI21xp5_ASAP7_75t_L g11039 ( 
.A1(n_10549),
.A2(n_1042),
.B(n_1043),
.Y(n_11039)
);

OAI21x1_ASAP7_75t_L g11040 ( 
.A1(n_10504),
.A2(n_1043),
.B(n_1044),
.Y(n_11040)
);

BUFx10_ASAP7_75t_L g11041 ( 
.A(n_10510),
.Y(n_11041)
);

NOR2xp67_ASAP7_75t_SL g11042 ( 
.A(n_10522),
.B(n_1043),
.Y(n_11042)
);

CKINVDCx5p33_ASAP7_75t_R g11043 ( 
.A(n_10593),
.Y(n_11043)
);

INVx1_ASAP7_75t_L g11044 ( 
.A(n_10588),
.Y(n_11044)
);

BUFx2_ASAP7_75t_L g11045 ( 
.A(n_10440),
.Y(n_11045)
);

NAND2xp5_ASAP7_75t_L g11046 ( 
.A(n_10588),
.B(n_1044),
.Y(n_11046)
);

AO32x2_ASAP7_75t_L g11047 ( 
.A1(n_10358),
.A2(n_1046),
.A3(n_1044),
.B1(n_1045),
.B2(n_1047),
.Y(n_11047)
);

INVx1_ASAP7_75t_L g11048 ( 
.A(n_10614),
.Y(n_11048)
);

NAND2xp5_ASAP7_75t_L g11049 ( 
.A(n_10614),
.B(n_1045),
.Y(n_11049)
);

AOI211x1_ASAP7_75t_L g11050 ( 
.A1(n_10431),
.A2(n_1049),
.B(n_1047),
.C(n_1048),
.Y(n_11050)
);

OAI21x1_ASAP7_75t_L g11051 ( 
.A1(n_10528),
.A2(n_1047),
.B(n_1048),
.Y(n_11051)
);

NAND3xp33_ASAP7_75t_L g11052 ( 
.A(n_10319),
.B(n_1048),
.C(n_1049),
.Y(n_11052)
);

NOR2xp33_ASAP7_75t_L g11053 ( 
.A(n_10535),
.B(n_1049),
.Y(n_11053)
);

NOR4xp25_ASAP7_75t_L g11054 ( 
.A(n_10587),
.B(n_1052),
.C(n_1050),
.D(n_1051),
.Y(n_11054)
);

OAI21x1_ASAP7_75t_L g11055 ( 
.A1(n_10242),
.A2(n_1050),
.B(n_1053),
.Y(n_11055)
);

OAI21x1_ASAP7_75t_L g11056 ( 
.A1(n_10214),
.A2(n_1053),
.B(n_1054),
.Y(n_11056)
);

BUFx6f_ASAP7_75t_L g11057 ( 
.A(n_10636),
.Y(n_11057)
);

INVx2_ASAP7_75t_L g11058 ( 
.A(n_10449),
.Y(n_11058)
);

INVx2_ASAP7_75t_L g11059 ( 
.A(n_10449),
.Y(n_11059)
);

NAND3x1_ASAP7_75t_L g11060 ( 
.A(n_10525),
.B(n_1053),
.C(n_1054),
.Y(n_11060)
);

A2O1A1Ixp33_ASAP7_75t_L g11061 ( 
.A1(n_10485),
.A2(n_1057),
.B(n_1055),
.C(n_1056),
.Y(n_11061)
);

NAND3x1_ASAP7_75t_L g11062 ( 
.A(n_10362),
.B(n_1055),
.C(n_1056),
.Y(n_11062)
);

AO31x2_ASAP7_75t_L g11063 ( 
.A1(n_10333),
.A2(n_1057),
.A3(n_1055),
.B(n_1056),
.Y(n_11063)
);

NOR2xp67_ASAP7_75t_L g11064 ( 
.A(n_10533),
.B(n_1057),
.Y(n_11064)
);

INVx2_ASAP7_75t_L g11065 ( 
.A(n_10227),
.Y(n_11065)
);

NAND2xp5_ASAP7_75t_SL g11066 ( 
.A(n_10212),
.B(n_1058),
.Y(n_11066)
);

CKINVDCx5p33_ASAP7_75t_R g11067 ( 
.A(n_10532),
.Y(n_11067)
);

AOI21xp5_ASAP7_75t_L g11068 ( 
.A1(n_10560),
.A2(n_1058),
.B(n_1059),
.Y(n_11068)
);

OAI21x1_ASAP7_75t_L g11069 ( 
.A1(n_10279),
.A2(n_1058),
.B(n_1059),
.Y(n_11069)
);

CKINVDCx5p33_ASAP7_75t_R g11070 ( 
.A(n_10605),
.Y(n_11070)
);

NAND2xp5_ASAP7_75t_L g11071 ( 
.A(n_10266),
.B(n_10402),
.Y(n_11071)
);

AO31x2_ASAP7_75t_L g11072 ( 
.A1(n_10410),
.A2(n_10539),
.A3(n_10460),
.B(n_10543),
.Y(n_11072)
);

OAI21x1_ASAP7_75t_L g11073 ( 
.A1(n_10286),
.A2(n_1059),
.B(n_1060),
.Y(n_11073)
);

AND2x4_ASAP7_75t_L g11074 ( 
.A(n_10637),
.B(n_1060),
.Y(n_11074)
);

AOI221x1_ASAP7_75t_L g11075 ( 
.A1(n_10352),
.A2(n_1062),
.B1(n_1060),
.B2(n_1061),
.C(n_1063),
.Y(n_11075)
);

INVx1_ASAP7_75t_L g11076 ( 
.A(n_10266),
.Y(n_11076)
);

NAND2xp5_ASAP7_75t_L g11077 ( 
.A(n_10359),
.B(n_1061),
.Y(n_11077)
);

OAI21x1_ASAP7_75t_L g11078 ( 
.A1(n_10645),
.A2(n_1062),
.B(n_1063),
.Y(n_11078)
);

AOI21xp5_ASAP7_75t_L g11079 ( 
.A1(n_10456),
.A2(n_1062),
.B(n_1063),
.Y(n_11079)
);

BUFx2_ASAP7_75t_L g11080 ( 
.A(n_10219),
.Y(n_11080)
);

CKINVDCx6p67_ASAP7_75t_R g11081 ( 
.A(n_10618),
.Y(n_11081)
);

NAND2xp33_ASAP7_75t_R g11082 ( 
.A(n_10494),
.B(n_1064),
.Y(n_11082)
);

NOR2xp33_ASAP7_75t_L g11083 ( 
.A(n_10573),
.B(n_1064),
.Y(n_11083)
);

NAND3xp33_ASAP7_75t_L g11084 ( 
.A(n_10607),
.B(n_1064),
.C(n_1065),
.Y(n_11084)
);

AND2x6_ASAP7_75t_L g11085 ( 
.A(n_11035),
.B(n_10527),
.Y(n_11085)
);

CKINVDCx9p33_ASAP7_75t_R g11086 ( 
.A(n_10787),
.Y(n_11086)
);

NAND2xp5_ASAP7_75t_L g11087 ( 
.A(n_10698),
.B(n_10298),
.Y(n_11087)
);

INVx1_ASAP7_75t_L g11088 ( 
.A(n_10652),
.Y(n_11088)
);

INVx2_ASAP7_75t_L g11089 ( 
.A(n_10667),
.Y(n_11089)
);

INVx1_ASAP7_75t_SL g11090 ( 
.A(n_10931),
.Y(n_11090)
);

AO21x2_ASAP7_75t_L g11091 ( 
.A1(n_11076),
.A2(n_10612),
.B(n_10475),
.Y(n_11091)
);

INVx1_ASAP7_75t_L g11092 ( 
.A(n_10656),
.Y(n_11092)
);

BUFx8_ASAP7_75t_L g11093 ( 
.A(n_10831),
.Y(n_11093)
);

INVx3_ASAP7_75t_L g11094 ( 
.A(n_10671),
.Y(n_11094)
);

INVx1_ASAP7_75t_L g11095 ( 
.A(n_10764),
.Y(n_11095)
);

OAI21x1_ASAP7_75t_L g11096 ( 
.A1(n_11058),
.A2(n_10546),
.B(n_10531),
.Y(n_11096)
);

OAI21x1_ASAP7_75t_L g11097 ( 
.A1(n_11059),
.A2(n_10551),
.B(n_10548),
.Y(n_11097)
);

OAI21x1_ASAP7_75t_L g11098 ( 
.A1(n_11065),
.A2(n_10408),
.B(n_10407),
.Y(n_11098)
);

OAI21x1_ASAP7_75t_L g11099 ( 
.A1(n_10990),
.A2(n_10415),
.B(n_10411),
.Y(n_11099)
);

AO31x2_ASAP7_75t_L g11100 ( 
.A1(n_11080),
.A2(n_10458),
.A3(n_10493),
.B(n_1068),
.Y(n_11100)
);

INVx3_ASAP7_75t_L g11101 ( 
.A(n_10671),
.Y(n_11101)
);

BUFx2_ASAP7_75t_L g11102 ( 
.A(n_10658),
.Y(n_11102)
);

BUFx3_ASAP7_75t_L g11103 ( 
.A(n_10744),
.Y(n_11103)
);

AND2x2_ASAP7_75t_L g11104 ( 
.A(n_10679),
.B(n_10608),
.Y(n_11104)
);

OAI21x1_ASAP7_75t_L g11105 ( 
.A1(n_11003),
.A2(n_10424),
.B(n_10423),
.Y(n_11105)
);

BUFx3_ASAP7_75t_L g11106 ( 
.A(n_10761),
.Y(n_11106)
);

BUFx8_ASAP7_75t_L g11107 ( 
.A(n_10771),
.Y(n_11107)
);

INVx1_ASAP7_75t_SL g11108 ( 
.A(n_10784),
.Y(n_11108)
);

OAI21x1_ASAP7_75t_L g11109 ( 
.A1(n_11032),
.A2(n_10448),
.B(n_10441),
.Y(n_11109)
);

AOI21x1_ASAP7_75t_L g11110 ( 
.A1(n_10985),
.A2(n_10594),
.B(n_10591),
.Y(n_11110)
);

AND2x4_ASAP7_75t_L g11111 ( 
.A(n_10734),
.B(n_10601),
.Y(n_11111)
);

AND2x2_ASAP7_75t_L g11112 ( 
.A(n_10691),
.B(n_10294),
.Y(n_11112)
);

HB1xp67_ASAP7_75t_L g11113 ( 
.A(n_10754),
.Y(n_11113)
);

OA21x2_ASAP7_75t_L g11114 ( 
.A1(n_10762),
.A2(n_10305),
.B(n_1066),
.Y(n_11114)
);

INVx2_ASAP7_75t_L g11115 ( 
.A(n_10711),
.Y(n_11115)
);

AND2x4_ASAP7_75t_L g11116 ( 
.A(n_10856),
.B(n_1066),
.Y(n_11116)
);

OAI21x1_ASAP7_75t_L g11117 ( 
.A1(n_11038),
.A2(n_1067),
.B(n_1068),
.Y(n_11117)
);

BUFx3_ASAP7_75t_L g11118 ( 
.A(n_10761),
.Y(n_11118)
);

AND2x2_ASAP7_75t_L g11119 ( 
.A(n_10769),
.B(n_1067),
.Y(n_11119)
);

INVx3_ASAP7_75t_SL g11120 ( 
.A(n_10781),
.Y(n_11120)
);

INVx1_ASAP7_75t_L g11121 ( 
.A(n_10706),
.Y(n_11121)
);

OAI21x1_ASAP7_75t_L g11122 ( 
.A1(n_11044),
.A2(n_1068),
.B(n_1069),
.Y(n_11122)
);

AO21x1_ASAP7_75t_L g11123 ( 
.A1(n_10657),
.A2(n_1069),
.B(n_1070),
.Y(n_11123)
);

INVx8_ASAP7_75t_L g11124 ( 
.A(n_10710),
.Y(n_11124)
);

OAI22xp5_ASAP7_75t_L g11125 ( 
.A1(n_11018),
.A2(n_1072),
.B1(n_1070),
.B2(n_1071),
.Y(n_11125)
);

OAI22xp5_ASAP7_75t_L g11126 ( 
.A1(n_11018),
.A2(n_1074),
.B1(n_1071),
.B2(n_1072),
.Y(n_11126)
);

NAND3xp33_ASAP7_75t_L g11127 ( 
.A(n_10840),
.B(n_1071),
.C(n_1072),
.Y(n_11127)
);

OAI21x1_ASAP7_75t_L g11128 ( 
.A1(n_11048),
.A2(n_1074),
.B(n_1075),
.Y(n_11128)
);

AO21x2_ASAP7_75t_L g11129 ( 
.A1(n_11017),
.A2(n_1075),
.B(n_1076),
.Y(n_11129)
);

NAND2xp5_ASAP7_75t_L g11130 ( 
.A(n_10799),
.B(n_1076),
.Y(n_11130)
);

OA21x2_ASAP7_75t_L g11131 ( 
.A1(n_10914),
.A2(n_1076),
.B(n_1077),
.Y(n_11131)
);

INVx1_ASAP7_75t_L g11132 ( 
.A(n_10708),
.Y(n_11132)
);

OAI21x1_ASAP7_75t_SL g11133 ( 
.A1(n_10745),
.A2(n_1077),
.B(n_1078),
.Y(n_11133)
);

OAI21x1_ASAP7_75t_L g11134 ( 
.A1(n_10678),
.A2(n_1077),
.B(n_1078),
.Y(n_11134)
);

INVx1_ASAP7_75t_L g11135 ( 
.A(n_10714),
.Y(n_11135)
);

BUFx6f_ASAP7_75t_L g11136 ( 
.A(n_10847),
.Y(n_11136)
);

NAND2x1p5_ASAP7_75t_L g11137 ( 
.A(n_11035),
.B(n_1079),
.Y(n_11137)
);

BUFx2_ASAP7_75t_R g11138 ( 
.A(n_10948),
.Y(n_11138)
);

INVx3_ASAP7_75t_L g11139 ( 
.A(n_10702),
.Y(n_11139)
);

INVx8_ASAP7_75t_L g11140 ( 
.A(n_10710),
.Y(n_11140)
);

OAI21x1_ASAP7_75t_L g11141 ( 
.A1(n_11071),
.A2(n_1079),
.B(n_1081),
.Y(n_11141)
);

AND2x4_ASAP7_75t_L g11142 ( 
.A(n_10776),
.B(n_1079),
.Y(n_11142)
);

AND2x2_ASAP7_75t_L g11143 ( 
.A(n_11001),
.B(n_1082),
.Y(n_11143)
);

OAI21x1_ASAP7_75t_SL g11144 ( 
.A1(n_10676),
.A2(n_1082),
.B(n_1083),
.Y(n_11144)
);

OAI21x1_ASAP7_75t_L g11145 ( 
.A1(n_10746),
.A2(n_1082),
.B(n_1083),
.Y(n_11145)
);

INVx2_ASAP7_75t_SL g11146 ( 
.A(n_10941),
.Y(n_11146)
);

OA21x2_ASAP7_75t_L g11147 ( 
.A1(n_10674),
.A2(n_1084),
.B(n_1085),
.Y(n_11147)
);

AO31x2_ASAP7_75t_L g11148 ( 
.A1(n_10997),
.A2(n_1086),
.A3(n_1084),
.B(n_1085),
.Y(n_11148)
);

AO21x2_ASAP7_75t_L g11149 ( 
.A1(n_10839),
.A2(n_1086),
.B(n_1087),
.Y(n_11149)
);

OAI21x1_ASAP7_75t_L g11150 ( 
.A1(n_11046),
.A2(n_1087),
.B(n_1088),
.Y(n_11150)
);

OAI21x1_ASAP7_75t_L g11151 ( 
.A1(n_11049),
.A2(n_1087),
.B(n_1088),
.Y(n_11151)
);

OAI21x1_ASAP7_75t_L g11152 ( 
.A1(n_10919),
.A2(n_1090),
.B(n_1091),
.Y(n_11152)
);

NOR2xp33_ASAP7_75t_L g11153 ( 
.A(n_10689),
.B(n_1090),
.Y(n_11153)
);

OAI21x1_ASAP7_75t_L g11154 ( 
.A1(n_10827),
.A2(n_1090),
.B(n_1091),
.Y(n_11154)
);

NAND2x1p5_ASAP7_75t_L g11155 ( 
.A(n_10682),
.B(n_1091),
.Y(n_11155)
);

BUFx2_ASAP7_75t_L g11156 ( 
.A(n_10696),
.Y(n_11156)
);

OR2x6_ASAP7_75t_L g11157 ( 
.A(n_10811),
.B(n_1092),
.Y(n_11157)
);

OAI21x1_ASAP7_75t_L g11158 ( 
.A1(n_10741),
.A2(n_10653),
.B(n_10887),
.Y(n_11158)
);

OAI21x1_ASAP7_75t_L g11159 ( 
.A1(n_10663),
.A2(n_1092),
.B(n_1093),
.Y(n_11159)
);

NAND2x1p5_ASAP7_75t_L g11160 ( 
.A(n_10719),
.B(n_1092),
.Y(n_11160)
);

NAND2x1p5_ASAP7_75t_L g11161 ( 
.A(n_11031),
.B(n_1093),
.Y(n_11161)
);

BUFx5_ASAP7_75t_L g11162 ( 
.A(n_10900),
.Y(n_11162)
);

INVx8_ASAP7_75t_L g11163 ( 
.A(n_10843),
.Y(n_11163)
);

INVx2_ASAP7_75t_L g11164 ( 
.A(n_10850),
.Y(n_11164)
);

OA21x2_ASAP7_75t_L g11165 ( 
.A1(n_10665),
.A2(n_1093),
.B(n_1094),
.Y(n_11165)
);

AND2x4_ASAP7_75t_L g11166 ( 
.A(n_10826),
.B(n_1094),
.Y(n_11166)
);

INVx1_ASAP7_75t_L g11167 ( 
.A(n_10729),
.Y(n_11167)
);

OA21x2_ASAP7_75t_L g11168 ( 
.A1(n_10748),
.A2(n_10870),
.B(n_10852),
.Y(n_11168)
);

OAI21x1_ASAP7_75t_L g11169 ( 
.A1(n_10701),
.A2(n_1094),
.B(n_1095),
.Y(n_11169)
);

AO21x2_ASAP7_75t_L g11170 ( 
.A1(n_10720),
.A2(n_1095),
.B(n_1096),
.Y(n_11170)
);

NAND3xp33_ASAP7_75t_L g11171 ( 
.A(n_10782),
.B(n_1096),
.C(n_1097),
.Y(n_11171)
);

OA21x2_ASAP7_75t_L g11172 ( 
.A1(n_10878),
.A2(n_1096),
.B(n_1097),
.Y(n_11172)
);

NAND3xp33_ASAP7_75t_L g11173 ( 
.A(n_10649),
.B(n_1097),
.C(n_1098),
.Y(n_11173)
);

AND2x2_ASAP7_75t_L g11174 ( 
.A(n_10980),
.B(n_1098),
.Y(n_11174)
);

INVxp67_ASAP7_75t_L g11175 ( 
.A(n_10942),
.Y(n_11175)
);

OAI21x1_ASAP7_75t_L g11176 ( 
.A1(n_10722),
.A2(n_10724),
.B(n_10917),
.Y(n_11176)
);

OAI21x1_ASAP7_75t_SL g11177 ( 
.A1(n_10677),
.A2(n_1099),
.B(n_1100),
.Y(n_11177)
);

OAI21x1_ASAP7_75t_L g11178 ( 
.A1(n_10688),
.A2(n_1099),
.B(n_1100),
.Y(n_11178)
);

INVx1_ASAP7_75t_L g11179 ( 
.A(n_10913),
.Y(n_11179)
);

OAI21x1_ASAP7_75t_L g11180 ( 
.A1(n_10717),
.A2(n_1099),
.B(n_1101),
.Y(n_11180)
);

OA21x2_ASAP7_75t_L g11181 ( 
.A1(n_10938),
.A2(n_1101),
.B(n_1102),
.Y(n_11181)
);

NAND2xp5_ASAP7_75t_L g11182 ( 
.A(n_11013),
.B(n_1101),
.Y(n_11182)
);

INVx2_ASAP7_75t_L g11183 ( 
.A(n_10858),
.Y(n_11183)
);

OAI21x1_ASAP7_75t_L g11184 ( 
.A1(n_10672),
.A2(n_1102),
.B(n_1103),
.Y(n_11184)
);

OAI21x1_ASAP7_75t_L g11185 ( 
.A1(n_10755),
.A2(n_1104),
.B(n_1105),
.Y(n_11185)
);

HB1xp67_ASAP7_75t_L g11186 ( 
.A(n_11045),
.Y(n_11186)
);

INVx4_ASAP7_75t_L g11187 ( 
.A(n_10785),
.Y(n_11187)
);

AND2x4_ASAP7_75t_L g11188 ( 
.A(n_10851),
.B(n_1104),
.Y(n_11188)
);

INVx1_ASAP7_75t_L g11189 ( 
.A(n_10772),
.Y(n_11189)
);

CKINVDCx5p33_ASAP7_75t_R g11190 ( 
.A(n_10929),
.Y(n_11190)
);

AND2x4_ASAP7_75t_SL g11191 ( 
.A(n_10785),
.B(n_1104),
.Y(n_11191)
);

INVx4_ASAP7_75t_L g11192 ( 
.A(n_10893),
.Y(n_11192)
);

AND2x4_ASAP7_75t_L g11193 ( 
.A(n_10660),
.B(n_1105),
.Y(n_11193)
);

BUFx3_ASAP7_75t_L g11194 ( 
.A(n_10923),
.Y(n_11194)
);

INVx6_ASAP7_75t_L g11195 ( 
.A(n_10968),
.Y(n_11195)
);

AO21x1_ASAP7_75t_L g11196 ( 
.A1(n_10987),
.A2(n_1106),
.B(n_1107),
.Y(n_11196)
);

INVx1_ASAP7_75t_L g11197 ( 
.A(n_10773),
.Y(n_11197)
);

NOR2xp33_ASAP7_75t_L g11198 ( 
.A(n_10906),
.B(n_10892),
.Y(n_11198)
);

AO21x2_ASAP7_75t_L g11199 ( 
.A1(n_10695),
.A2(n_1106),
.B(n_1107),
.Y(n_11199)
);

BUFx6f_ASAP7_75t_L g11200 ( 
.A(n_10893),
.Y(n_11200)
);

AO21x2_ASAP7_75t_L g11201 ( 
.A1(n_10832),
.A2(n_1107),
.B(n_1108),
.Y(n_11201)
);

INVx2_ASAP7_75t_L g11202 ( 
.A(n_10861),
.Y(n_11202)
);

INVx1_ASAP7_75t_L g11203 ( 
.A(n_10790),
.Y(n_11203)
);

OA21x2_ASAP7_75t_L g11204 ( 
.A1(n_10794),
.A2(n_1108),
.B(n_1109),
.Y(n_11204)
);

NOR2x1_ASAP7_75t_SL g11205 ( 
.A(n_10821),
.B(n_1108),
.Y(n_11205)
);

NOR2xp67_ASAP7_75t_L g11206 ( 
.A(n_10800),
.B(n_1109),
.Y(n_11206)
);

OAI21x1_ASAP7_75t_SL g11207 ( 
.A1(n_10963),
.A2(n_1110),
.B(n_1111),
.Y(n_11207)
);

AOI221xp5_ASAP7_75t_L g11208 ( 
.A1(n_10986),
.A2(n_1112),
.B1(n_1110),
.B2(n_1111),
.C(n_1113),
.Y(n_11208)
);

OAI21x1_ASAP7_75t_L g11209 ( 
.A1(n_10979),
.A2(n_1110),
.B(n_1111),
.Y(n_11209)
);

INVx6_ASAP7_75t_L g11210 ( 
.A(n_10968),
.Y(n_11210)
);

AND2x6_ASAP7_75t_L g11211 ( 
.A(n_11015),
.B(n_1113),
.Y(n_11211)
);

OAI21x1_ASAP7_75t_SL g11212 ( 
.A1(n_10820),
.A2(n_1113),
.B(n_1114),
.Y(n_11212)
);

AND2x2_ASAP7_75t_L g11213 ( 
.A(n_10941),
.B(n_1114),
.Y(n_11213)
);

OA21x2_ASAP7_75t_L g11214 ( 
.A1(n_10795),
.A2(n_1114),
.B(n_1115),
.Y(n_11214)
);

BUFx2_ASAP7_75t_L g11215 ( 
.A(n_10916),
.Y(n_11215)
);

OAI21x1_ASAP7_75t_L g11216 ( 
.A1(n_10697),
.A2(n_1115),
.B(n_1116),
.Y(n_11216)
);

AO21x2_ASAP7_75t_L g11217 ( 
.A1(n_10846),
.A2(n_1116),
.B(n_1117),
.Y(n_11217)
);

AO21x1_ASAP7_75t_L g11218 ( 
.A1(n_10960),
.A2(n_1117),
.B(n_1118),
.Y(n_11218)
);

AOI21x1_ASAP7_75t_L g11219 ( 
.A1(n_10864),
.A2(n_1117),
.B(n_1118),
.Y(n_11219)
);

BUFx3_ASAP7_75t_L g11220 ( 
.A(n_10962),
.Y(n_11220)
);

INVx1_ASAP7_75t_L g11221 ( 
.A(n_10797),
.Y(n_11221)
);

OAI21x1_ASAP7_75t_L g11222 ( 
.A1(n_10824),
.A2(n_1118),
.B(n_1119),
.Y(n_11222)
);

NOR2xp67_ASAP7_75t_L g11223 ( 
.A(n_10760),
.B(n_1119),
.Y(n_11223)
);

INVx1_ASAP7_75t_L g11224 ( 
.A(n_10845),
.Y(n_11224)
);

AO21x2_ASAP7_75t_L g11225 ( 
.A1(n_10749),
.A2(n_1120),
.B(n_1121),
.Y(n_11225)
);

OAI21x1_ASAP7_75t_L g11226 ( 
.A1(n_10750),
.A2(n_1121),
.B(n_1122),
.Y(n_11226)
);

OAI21x1_ASAP7_75t_L g11227 ( 
.A1(n_10758),
.A2(n_1121),
.B(n_1122),
.Y(n_11227)
);

OAI21x1_ASAP7_75t_L g11228 ( 
.A1(n_10767),
.A2(n_1123),
.B(n_1124),
.Y(n_11228)
);

AOI22x1_ASAP7_75t_L g11229 ( 
.A1(n_10768),
.A2(n_1126),
.B1(n_1123),
.B2(n_1124),
.Y(n_11229)
);

BUFx4f_ASAP7_75t_SL g11230 ( 
.A(n_10916),
.Y(n_11230)
);

AND2x4_ASAP7_75t_L g11231 ( 
.A(n_10654),
.B(n_1123),
.Y(n_11231)
);

AO21x2_ASAP7_75t_L g11232 ( 
.A1(n_10766),
.A2(n_1126),
.B(n_1127),
.Y(n_11232)
);

OAI21xp5_ASAP7_75t_L g11233 ( 
.A1(n_10842),
.A2(n_1126),
.B(n_1127),
.Y(n_11233)
);

INVx2_ASAP7_75t_L g11234 ( 
.A(n_10877),
.Y(n_11234)
);

AOI21xp5_ASAP7_75t_L g11235 ( 
.A1(n_10965),
.A2(n_1127),
.B(n_1128),
.Y(n_11235)
);

NAND2xp5_ASAP7_75t_L g11236 ( 
.A(n_11023),
.B(n_1128),
.Y(n_11236)
);

INVx1_ASAP7_75t_L g11237 ( 
.A(n_10954),
.Y(n_11237)
);

INVx8_ASAP7_75t_L g11238 ( 
.A(n_10843),
.Y(n_11238)
);

AND2x2_ASAP7_75t_L g11239 ( 
.A(n_10752),
.B(n_1128),
.Y(n_11239)
);

BUFx12f_ASAP7_75t_L g11240 ( 
.A(n_10903),
.Y(n_11240)
);

OAI21x1_ASAP7_75t_L g11241 ( 
.A1(n_10779),
.A2(n_1129),
.B(n_1130),
.Y(n_11241)
);

NAND2xp5_ASAP7_75t_L g11242 ( 
.A(n_10704),
.B(n_1129),
.Y(n_11242)
);

NAND3xp33_ASAP7_75t_L g11243 ( 
.A(n_10655),
.B(n_1129),
.C(n_1130),
.Y(n_11243)
);

NAND2xp5_ASAP7_75t_L g11244 ( 
.A(n_10735),
.B(n_1131),
.Y(n_11244)
);

AO21x2_ASAP7_75t_L g11245 ( 
.A1(n_10737),
.A2(n_1131),
.B(n_1132),
.Y(n_11245)
);

AO21x2_ASAP7_75t_L g11246 ( 
.A1(n_10747),
.A2(n_1131),
.B(n_1132),
.Y(n_11246)
);

BUFx3_ASAP7_75t_L g11247 ( 
.A(n_10904),
.Y(n_11247)
);

INVx1_ASAP7_75t_L g11248 ( 
.A(n_10978),
.Y(n_11248)
);

AOI22x1_ASAP7_75t_L g11249 ( 
.A1(n_10757),
.A2(n_1135),
.B1(n_1133),
.B2(n_1134),
.Y(n_11249)
);

AOI21x1_ASAP7_75t_L g11250 ( 
.A1(n_10920),
.A2(n_10921),
.B(n_11011),
.Y(n_11250)
);

AND2x4_ASAP7_75t_L g11251 ( 
.A(n_10654),
.B(n_1133),
.Y(n_11251)
);

AO21x2_ASAP7_75t_L g11252 ( 
.A1(n_10727),
.A2(n_1133),
.B(n_1134),
.Y(n_11252)
);

INVx1_ASAP7_75t_L g11253 ( 
.A(n_10885),
.Y(n_11253)
);

BUFx3_ASAP7_75t_L g11254 ( 
.A(n_11043),
.Y(n_11254)
);

OAI21xp5_ASAP7_75t_L g11255 ( 
.A1(n_10651),
.A2(n_1134),
.B(n_1135),
.Y(n_11255)
);

INVx1_ASAP7_75t_L g11256 ( 
.A(n_10888),
.Y(n_11256)
);

AOI22xp33_ASAP7_75t_L g11257 ( 
.A1(n_10751),
.A2(n_1137),
.B1(n_1135),
.B2(n_1136),
.Y(n_11257)
);

OA21x2_ASAP7_75t_L g11258 ( 
.A1(n_10949),
.A2(n_1136),
.B(n_1137),
.Y(n_11258)
);

NOR2xp33_ASAP7_75t_L g11259 ( 
.A(n_10731),
.B(n_1136),
.Y(n_11259)
);

OAI21x1_ASAP7_75t_L g11260 ( 
.A1(n_10791),
.A2(n_1138),
.B(n_1139),
.Y(n_11260)
);

NAND2xp5_ASAP7_75t_L g11261 ( 
.A(n_10775),
.B(n_1138),
.Y(n_11261)
);

INVx1_ASAP7_75t_L g11262 ( 
.A(n_10974),
.Y(n_11262)
);

HB1xp67_ASAP7_75t_L g11263 ( 
.A(n_10783),
.Y(n_11263)
);

HB1xp67_ASAP7_75t_L g11264 ( 
.A(n_10796),
.Y(n_11264)
);

INVx1_ASAP7_75t_L g11265 ( 
.A(n_10673),
.Y(n_11265)
);

BUFx2_ASAP7_75t_R g11266 ( 
.A(n_10992),
.Y(n_11266)
);

OAI22xp5_ASAP7_75t_L g11267 ( 
.A1(n_10927),
.A2(n_1141),
.B1(n_1139),
.B2(n_1140),
.Y(n_11267)
);

INVx3_ASAP7_75t_L g11268 ( 
.A(n_10756),
.Y(n_11268)
);

BUFx4f_ASAP7_75t_L g11269 ( 
.A(n_10903),
.Y(n_11269)
);

OAI21xp5_ASAP7_75t_L g11270 ( 
.A1(n_10830),
.A2(n_11060),
.B(n_10812),
.Y(n_11270)
);

OAI21x1_ASAP7_75t_L g11271 ( 
.A1(n_10792),
.A2(n_1139),
.B(n_1140),
.Y(n_11271)
);

NAND2x1_ASAP7_75t_L g11272 ( 
.A(n_10821),
.B(n_1140),
.Y(n_11272)
);

OAI21x1_ASAP7_75t_L g11273 ( 
.A1(n_10694),
.A2(n_10922),
.B(n_10815),
.Y(n_11273)
);

OA21x2_ASAP7_75t_L g11274 ( 
.A1(n_10805),
.A2(n_1141),
.B(n_1142),
.Y(n_11274)
);

AO21x2_ASAP7_75t_L g11275 ( 
.A1(n_10798),
.A2(n_1141),
.B(n_1142),
.Y(n_11275)
);

OAI21xp5_ASAP7_75t_L g11276 ( 
.A1(n_10675),
.A2(n_1142),
.B(n_1143),
.Y(n_11276)
);

BUFx3_ASAP7_75t_L g11277 ( 
.A(n_10982),
.Y(n_11277)
);

AO21x2_ASAP7_75t_L g11278 ( 
.A1(n_10801),
.A2(n_1143),
.B(n_1144),
.Y(n_11278)
);

NAND2x1p5_ASAP7_75t_L g11279 ( 
.A(n_10687),
.B(n_1145),
.Y(n_11279)
);

BUFx6f_ASAP7_75t_L g11280 ( 
.A(n_10940),
.Y(n_11280)
);

INVx2_ASAP7_75t_L g11281 ( 
.A(n_11057),
.Y(n_11281)
);

AOI21xp33_ASAP7_75t_L g11282 ( 
.A1(n_11082),
.A2(n_1145),
.B(n_1146),
.Y(n_11282)
);

CKINVDCx6p67_ASAP7_75t_R g11283 ( 
.A(n_10829),
.Y(n_11283)
);

NAND2x1p5_ASAP7_75t_L g11284 ( 
.A(n_10975),
.B(n_1145),
.Y(n_11284)
);

AOI22xp33_ASAP7_75t_L g11285 ( 
.A1(n_10837),
.A2(n_1148),
.B1(n_1146),
.B2(n_1147),
.Y(n_11285)
);

OR2x6_ASAP7_75t_L g11286 ( 
.A(n_10829),
.B(n_1146),
.Y(n_11286)
);

OA21x2_ASAP7_75t_L g11287 ( 
.A1(n_10789),
.A2(n_1147),
.B(n_1148),
.Y(n_11287)
);

INVx1_ASAP7_75t_L g11288 ( 
.A(n_10713),
.Y(n_11288)
);

OAI21xp5_ASAP7_75t_L g11289 ( 
.A1(n_10650),
.A2(n_1149),
.B(n_1150),
.Y(n_11289)
);

OAI21x1_ASAP7_75t_L g11290 ( 
.A1(n_10709),
.A2(n_1149),
.B(n_1150),
.Y(n_11290)
);

INVx2_ASAP7_75t_L g11291 ( 
.A(n_11057),
.Y(n_11291)
);

BUFx6f_ASAP7_75t_L g11292 ( 
.A(n_10721),
.Y(n_11292)
);

OR3x4_ASAP7_75t_SL g11293 ( 
.A(n_10705),
.B(n_1149),
.C(n_1150),
.Y(n_11293)
);

AO21x2_ASAP7_75t_L g11294 ( 
.A1(n_10818),
.A2(n_1152),
.B(n_1153),
.Y(n_11294)
);

NAND2x1p5_ASAP7_75t_L g11295 ( 
.A(n_10976),
.B(n_1152),
.Y(n_11295)
);

INVx2_ASAP7_75t_L g11296 ( 
.A(n_10836),
.Y(n_11296)
);

OAI21xp5_ASAP7_75t_L g11297 ( 
.A1(n_10777),
.A2(n_1152),
.B(n_1153),
.Y(n_11297)
);

OAI21x1_ASAP7_75t_L g11298 ( 
.A1(n_10718),
.A2(n_1154),
.B(n_1155),
.Y(n_11298)
);

O2A1O1Ixp33_ASAP7_75t_L g11299 ( 
.A1(n_10966),
.A2(n_1156),
.B(n_1154),
.C(n_1155),
.Y(n_11299)
);

NAND2xp5_ASAP7_75t_L g11300 ( 
.A(n_10841),
.B(n_1154),
.Y(n_11300)
);

INVx3_ASAP7_75t_L g11301 ( 
.A(n_10953),
.Y(n_11301)
);

NAND3xp33_ASAP7_75t_L g11302 ( 
.A(n_10884),
.B(n_1155),
.C(n_1156),
.Y(n_11302)
);

NAND2xp5_ASAP7_75t_L g11303 ( 
.A(n_10844),
.B(n_1157),
.Y(n_11303)
);

AOI21x1_ASAP7_75t_L g11304 ( 
.A1(n_11005),
.A2(n_1157),
.B(n_1158),
.Y(n_11304)
);

OAI22xp5_ASAP7_75t_L g11305 ( 
.A1(n_10703),
.A2(n_1161),
.B1(n_1159),
.B2(n_1160),
.Y(n_11305)
);

OAI21x1_ASAP7_75t_L g11306 ( 
.A1(n_10726),
.A2(n_1159),
.B(n_1160),
.Y(n_11306)
);

CKINVDCx20_ASAP7_75t_R g11307 ( 
.A(n_10896),
.Y(n_11307)
);

BUFx4f_ASAP7_75t_L g11308 ( 
.A(n_10681),
.Y(n_11308)
);

INVx4_ASAP7_75t_L g11309 ( 
.A(n_10814),
.Y(n_11309)
);

AO21x2_ASAP7_75t_L g11310 ( 
.A1(n_10822),
.A2(n_1159),
.B(n_1160),
.Y(n_11310)
);

CKINVDCx6p67_ASAP7_75t_R g11311 ( 
.A(n_10808),
.Y(n_11311)
);

CKINVDCx5p33_ASAP7_75t_R g11312 ( 
.A(n_11041),
.Y(n_11312)
);

CKINVDCx5p33_ASAP7_75t_R g11313 ( 
.A(n_10874),
.Y(n_11313)
);

OAI21x1_ASAP7_75t_L g11314 ( 
.A1(n_10728),
.A2(n_1162),
.B(n_1163),
.Y(n_11314)
);

INVx2_ASAP7_75t_L g11315 ( 
.A(n_10730),
.Y(n_11315)
);

OAI21x1_ASAP7_75t_L g11316 ( 
.A1(n_10910),
.A2(n_1162),
.B(n_1163),
.Y(n_11316)
);

AO21x2_ASAP7_75t_L g11317 ( 
.A1(n_10823),
.A2(n_1164),
.B(n_1165),
.Y(n_11317)
);

INVx2_ASAP7_75t_L g11318 ( 
.A(n_10664),
.Y(n_11318)
);

BUFx2_ASAP7_75t_L g11319 ( 
.A(n_10953),
.Y(n_11319)
);

BUFx6f_ASAP7_75t_L g11320 ( 
.A(n_10984),
.Y(n_11320)
);

INVx2_ASAP7_75t_L g11321 ( 
.A(n_10664),
.Y(n_11321)
);

BUFx8_ASAP7_75t_L g11322 ( 
.A(n_10989),
.Y(n_11322)
);

INVx2_ASAP7_75t_L g11323 ( 
.A(n_11074),
.Y(n_11323)
);

INVx1_ASAP7_75t_SL g11324 ( 
.A(n_10991),
.Y(n_11324)
);

OAI21x1_ASAP7_75t_L g11325 ( 
.A1(n_10707),
.A2(n_1164),
.B(n_1165),
.Y(n_11325)
);

INVx3_ASAP7_75t_SL g11326 ( 
.A(n_11067),
.Y(n_11326)
);

AND2x4_ASAP7_75t_L g11327 ( 
.A(n_11014),
.B(n_1164),
.Y(n_11327)
);

BUFx2_ASAP7_75t_L g11328 ( 
.A(n_10953),
.Y(n_11328)
);

INVx5_ASAP7_75t_L g11329 ( 
.A(n_11014),
.Y(n_11329)
);

OAI21x1_ASAP7_75t_L g11330 ( 
.A1(n_11078),
.A2(n_1167),
.B(n_1168),
.Y(n_11330)
);

NAND2xp5_ASAP7_75t_L g11331 ( 
.A(n_10969),
.B(n_1167),
.Y(n_11331)
);

AO31x2_ASAP7_75t_L g11332 ( 
.A1(n_10659),
.A2(n_1169),
.A3(n_1167),
.B(n_1168),
.Y(n_11332)
);

NAND2xp5_ASAP7_75t_L g11333 ( 
.A(n_10994),
.B(n_1168),
.Y(n_11333)
);

AND2x4_ASAP7_75t_L g11334 ( 
.A(n_11004),
.B(n_1170),
.Y(n_11334)
);

BUFx3_ASAP7_75t_L g11335 ( 
.A(n_10895),
.Y(n_11335)
);

OAI21x1_ASAP7_75t_L g11336 ( 
.A1(n_10740),
.A2(n_10686),
.B(n_10680),
.Y(n_11336)
);

CKINVDCx16_ASAP7_75t_R g11337 ( 
.A(n_10897),
.Y(n_11337)
);

OAI21x1_ASAP7_75t_L g11338 ( 
.A1(n_10690),
.A2(n_10666),
.B(n_11077),
.Y(n_11338)
);

BUFx2_ASAP7_75t_L g11339 ( 
.A(n_11081),
.Y(n_11339)
);

OAI21x1_ASAP7_75t_L g11340 ( 
.A1(n_10743),
.A2(n_1170),
.B(n_1171),
.Y(n_11340)
);

AOI21xp5_ASAP7_75t_L g11341 ( 
.A1(n_10935),
.A2(n_1170),
.B(n_1171),
.Y(n_11341)
);

BUFx3_ASAP7_75t_L g11342 ( 
.A(n_11037),
.Y(n_11342)
);

NAND2xp5_ASAP7_75t_L g11343 ( 
.A(n_10793),
.B(n_1171),
.Y(n_11343)
);

OA21x2_ASAP7_75t_L g11344 ( 
.A1(n_11010),
.A2(n_1172),
.B(n_1173),
.Y(n_11344)
);

BUFx12f_ASAP7_75t_L g11345 ( 
.A(n_11070),
.Y(n_11345)
);

OA21x2_ASAP7_75t_L g11346 ( 
.A1(n_10788),
.A2(n_1172),
.B(n_1173),
.Y(n_11346)
);

BUFx6f_ASAP7_75t_L g11347 ( 
.A(n_10880),
.Y(n_11347)
);

CKINVDCx20_ASAP7_75t_R g11348 ( 
.A(n_11024),
.Y(n_11348)
);

BUFx2_ASAP7_75t_L g11349 ( 
.A(n_11009),
.Y(n_11349)
);

INVx1_ASAP7_75t_L g11350 ( 
.A(n_11002),
.Y(n_11350)
);

INVx3_ASAP7_75t_L g11351 ( 
.A(n_11028),
.Y(n_11351)
);

BUFx3_ASAP7_75t_L g11352 ( 
.A(n_10915),
.Y(n_11352)
);

INVx1_ASAP7_75t_L g11353 ( 
.A(n_11002),
.Y(n_11353)
);

INVx1_ASAP7_75t_L g11354 ( 
.A(n_11007),
.Y(n_11354)
);

OAI21x1_ASAP7_75t_L g11355 ( 
.A1(n_11000),
.A2(n_1172),
.B(n_1174),
.Y(n_11355)
);

NAND3xp33_ASAP7_75t_L g11356 ( 
.A(n_10833),
.B(n_1174),
.C(n_1175),
.Y(n_11356)
);

NAND2xp5_ASAP7_75t_L g11357 ( 
.A(n_10898),
.B(n_1174),
.Y(n_11357)
);

AND2x2_ASAP7_75t_L g11358 ( 
.A(n_10932),
.B(n_1175),
.Y(n_11358)
);

INVx2_ASAP7_75t_L g11359 ( 
.A(n_10875),
.Y(n_11359)
);

OAI21x1_ASAP7_75t_L g11360 ( 
.A1(n_10700),
.A2(n_1175),
.B(n_1176),
.Y(n_11360)
);

OAI21x1_ASAP7_75t_L g11361 ( 
.A1(n_10883),
.A2(n_1176),
.B(n_1177),
.Y(n_11361)
);

INVx6_ASAP7_75t_L g11362 ( 
.A(n_10668),
.Y(n_11362)
);

OA21x2_ASAP7_75t_L g11363 ( 
.A1(n_10901),
.A2(n_1176),
.B(n_1177),
.Y(n_11363)
);

AO21x1_ASAP7_75t_L g11364 ( 
.A1(n_10817),
.A2(n_1178),
.B(n_1179),
.Y(n_11364)
);

OAI21x1_ASAP7_75t_L g11365 ( 
.A1(n_10899),
.A2(n_1178),
.B(n_1179),
.Y(n_11365)
);

BUFx2_ASAP7_75t_L g11366 ( 
.A(n_10855),
.Y(n_11366)
);

BUFx12f_ASAP7_75t_L g11367 ( 
.A(n_10955),
.Y(n_11367)
);

INVx3_ASAP7_75t_L g11368 ( 
.A(n_10908),
.Y(n_11368)
);

INVx2_ASAP7_75t_L g11369 ( 
.A(n_10911),
.Y(n_11369)
);

INVx3_ASAP7_75t_L g11370 ( 
.A(n_10933),
.Y(n_11370)
);

INVx1_ASAP7_75t_L g11371 ( 
.A(n_11007),
.Y(n_11371)
);

INVx1_ASAP7_75t_L g11372 ( 
.A(n_11063),
.Y(n_11372)
);

INVx8_ASAP7_75t_L g11373 ( 
.A(n_10712),
.Y(n_11373)
);

INVx1_ASAP7_75t_L g11374 ( 
.A(n_11063),
.Y(n_11374)
);

OAI21xp5_ASAP7_75t_L g11375 ( 
.A1(n_10867),
.A2(n_1180),
.B(n_1181),
.Y(n_11375)
);

OAI21x1_ASAP7_75t_L g11376 ( 
.A1(n_10939),
.A2(n_1180),
.B(n_1181),
.Y(n_11376)
);

OAI21x1_ASAP7_75t_L g11377 ( 
.A1(n_10950),
.A2(n_1180),
.B(n_1181),
.Y(n_11377)
);

OAI21x1_ASAP7_75t_L g11378 ( 
.A1(n_10988),
.A2(n_1182),
.B(n_1183),
.Y(n_11378)
);

INVx1_ASAP7_75t_L g11379 ( 
.A(n_10763),
.Y(n_11379)
);

OAI21x1_ASAP7_75t_L g11380 ( 
.A1(n_11040),
.A2(n_1182),
.B(n_1183),
.Y(n_11380)
);

OA21x2_ASAP7_75t_L g11381 ( 
.A1(n_10956),
.A2(n_1182),
.B(n_1183),
.Y(n_11381)
);

OAI21x1_ASAP7_75t_L g11382 ( 
.A1(n_11051),
.A2(n_1184),
.B(n_1185),
.Y(n_11382)
);

NAND2xp5_ASAP7_75t_L g11383 ( 
.A(n_10958),
.B(n_1184),
.Y(n_11383)
);

NAND2xp5_ASAP7_75t_L g11384 ( 
.A(n_10995),
.B(n_1184),
.Y(n_11384)
);

OAI21x1_ASAP7_75t_L g11385 ( 
.A1(n_10865),
.A2(n_1185),
.B(n_1186),
.Y(n_11385)
);

BUFx3_ASAP7_75t_L g11386 ( 
.A(n_10943),
.Y(n_11386)
);

INVx1_ASAP7_75t_L g11387 ( 
.A(n_10763),
.Y(n_11387)
);

BUFx6f_ASAP7_75t_L g11388 ( 
.A(n_11016),
.Y(n_11388)
);

HB1xp67_ASAP7_75t_L g11389 ( 
.A(n_11025),
.Y(n_11389)
);

OAI21xp5_ASAP7_75t_L g11390 ( 
.A1(n_10715),
.A2(n_1185),
.B(n_1186),
.Y(n_11390)
);

OAI21x1_ASAP7_75t_L g11391 ( 
.A1(n_10866),
.A2(n_1187),
.B(n_1188),
.Y(n_11391)
);

BUFx2_ASAP7_75t_L g11392 ( 
.A(n_11027),
.Y(n_11392)
);

BUFx2_ASAP7_75t_R g11393 ( 
.A(n_11029),
.Y(n_11393)
);

OA21x2_ASAP7_75t_L g11394 ( 
.A1(n_10881),
.A2(n_1187),
.B(n_1188),
.Y(n_11394)
);

OAI21x1_ASAP7_75t_L g11395 ( 
.A1(n_10869),
.A2(n_1187),
.B(n_1188),
.Y(n_11395)
);

NAND2xp5_ASAP7_75t_L g11396 ( 
.A(n_10853),
.B(n_1189),
.Y(n_11396)
);

AO21x2_ASAP7_75t_L g11397 ( 
.A1(n_10669),
.A2(n_1189),
.B(n_1190),
.Y(n_11397)
);

BUFx6f_ASAP7_75t_L g11398 ( 
.A(n_10774),
.Y(n_11398)
);

INVx6_ASAP7_75t_L g11399 ( 
.A(n_10807),
.Y(n_11399)
);

NOR2x1_ASAP7_75t_R g11400 ( 
.A(n_10998),
.B(n_11066),
.Y(n_11400)
);

OAI21x1_ASAP7_75t_L g11401 ( 
.A1(n_10952),
.A2(n_10912),
.B(n_10803),
.Y(n_11401)
);

BUFx2_ASAP7_75t_R g11402 ( 
.A(n_10971),
.Y(n_11402)
);

OAI21x1_ASAP7_75t_L g11403 ( 
.A1(n_10804),
.A2(n_1190),
.B(n_1191),
.Y(n_11403)
);

INVx1_ASAP7_75t_L g11404 ( 
.A(n_10813),
.Y(n_11404)
);

INVx2_ASAP7_75t_L g11405 ( 
.A(n_10813),
.Y(n_11405)
);

INVx1_ASAP7_75t_L g11406 ( 
.A(n_10973),
.Y(n_11406)
);

AND2x4_ASAP7_75t_L g11407 ( 
.A(n_11064),
.B(n_1190),
.Y(n_11407)
);

NAND2x1p5_ASAP7_75t_L g11408 ( 
.A(n_10890),
.B(n_1191),
.Y(n_11408)
);

INVx1_ASAP7_75t_L g11409 ( 
.A(n_10973),
.Y(n_11409)
);

INVx2_ASAP7_75t_L g11410 ( 
.A(n_10819),
.Y(n_11410)
);

NAND2xp5_ASAP7_75t_L g11411 ( 
.A(n_11053),
.B(n_1192),
.Y(n_11411)
);

OAI21x1_ASAP7_75t_L g11412 ( 
.A1(n_10961),
.A2(n_11021),
.B(n_11019),
.Y(n_11412)
);

NOR2xp33_ASAP7_75t_SL g11413 ( 
.A(n_10981),
.B(n_1192),
.Y(n_11413)
);

OA21x2_ASAP7_75t_L g11414 ( 
.A1(n_10670),
.A2(n_1193),
.B(n_1194),
.Y(n_11414)
);

INVx1_ASAP7_75t_L g11415 ( 
.A(n_10872),
.Y(n_11415)
);

HB1xp67_ASAP7_75t_L g11416 ( 
.A(n_10872),
.Y(n_11416)
);

AND2x4_ASAP7_75t_L g11417 ( 
.A(n_10964),
.B(n_1193),
.Y(n_11417)
);

NOR2xp33_ASAP7_75t_L g11418 ( 
.A(n_10739),
.B(n_1193),
.Y(n_11418)
);

NAND2x1p5_ASAP7_75t_L g11419 ( 
.A(n_11042),
.B(n_1195),
.Y(n_11419)
);

INVx1_ASAP7_75t_L g11420 ( 
.A(n_11056),
.Y(n_11420)
);

NAND2x1p5_ASAP7_75t_L g11421 ( 
.A(n_11069),
.B(n_1196),
.Y(n_11421)
);

INVx2_ASAP7_75t_L g11422 ( 
.A(n_11073),
.Y(n_11422)
);

BUFx2_ASAP7_75t_R g11423 ( 
.A(n_10946),
.Y(n_11423)
);

NOR2xp33_ASAP7_75t_L g11424 ( 
.A(n_10889),
.B(n_1196),
.Y(n_11424)
);

NAND2xp5_ASAP7_75t_L g11425 ( 
.A(n_10699),
.B(n_10692),
.Y(n_11425)
);

OA21x2_ASAP7_75t_L g11426 ( 
.A1(n_10907),
.A2(n_1197),
.B(n_1198),
.Y(n_11426)
);

BUFx2_ASAP7_75t_L g11427 ( 
.A(n_11072),
.Y(n_11427)
);

OA21x2_ASAP7_75t_L g11428 ( 
.A1(n_10977),
.A2(n_1197),
.B(n_1198),
.Y(n_11428)
);

OAI21x1_ASAP7_75t_L g11429 ( 
.A1(n_11033),
.A2(n_1197),
.B(n_1199),
.Y(n_11429)
);

OAI21x1_ASAP7_75t_L g11430 ( 
.A1(n_10993),
.A2(n_1199),
.B(n_1200),
.Y(n_11430)
);

OR2x6_ASAP7_75t_L g11431 ( 
.A(n_11008),
.B(n_1200),
.Y(n_11431)
);

INVx4_ASAP7_75t_L g11432 ( 
.A(n_11006),
.Y(n_11432)
);

OAI21xp5_ASAP7_75t_L g11433 ( 
.A1(n_10930),
.A2(n_1201),
.B(n_1202),
.Y(n_11433)
);

BUFx2_ASAP7_75t_SL g11434 ( 
.A(n_11062),
.Y(n_11434)
);

INVx1_ASAP7_75t_L g11435 ( 
.A(n_11026),
.Y(n_11435)
);

AOI22xp33_ASAP7_75t_L g11436 ( 
.A1(n_10802),
.A2(n_1203),
.B1(n_1201),
.B2(n_1202),
.Y(n_11436)
);

INVx1_ASAP7_75t_L g11437 ( 
.A(n_10925),
.Y(n_11437)
);

OAI21x1_ASAP7_75t_L g11438 ( 
.A1(n_10999),
.A2(n_1203),
.B(n_1204),
.Y(n_11438)
);

CKINVDCx11_ASAP7_75t_R g11439 ( 
.A(n_10778),
.Y(n_11439)
);

BUFx3_ASAP7_75t_L g11440 ( 
.A(n_11055),
.Y(n_11440)
);

OA21x2_ASAP7_75t_L g11441 ( 
.A1(n_11012),
.A2(n_10849),
.B(n_11075),
.Y(n_11441)
);

AOI22xp33_ASAP7_75t_L g11442 ( 
.A1(n_10662),
.A2(n_1206),
.B1(n_1204),
.B2(n_1205),
.Y(n_11442)
);

OAI21xp5_ASAP7_75t_L g11443 ( 
.A1(n_10742),
.A2(n_1205),
.B(n_1206),
.Y(n_11443)
);

INVx1_ASAP7_75t_SL g11444 ( 
.A(n_10876),
.Y(n_11444)
);

AND2x4_ASAP7_75t_L g11445 ( 
.A(n_10648),
.B(n_1205),
.Y(n_11445)
);

OAI21x1_ASAP7_75t_L g11446 ( 
.A1(n_11301),
.A2(n_10909),
.B(n_10882),
.Y(n_11446)
);

AND2x4_ASAP7_75t_L g11447 ( 
.A(n_11094),
.B(n_11072),
.Y(n_11447)
);

OAI21x1_ASAP7_75t_L g11448 ( 
.A1(n_11176),
.A2(n_10780),
.B(n_10886),
.Y(n_11448)
);

OAI21x1_ASAP7_75t_L g11449 ( 
.A1(n_11087),
.A2(n_10857),
.B(n_10838),
.Y(n_11449)
);

OAI21x1_ASAP7_75t_L g11450 ( 
.A1(n_11158),
.A2(n_10944),
.B(n_10738),
.Y(n_11450)
);

OAI21x1_ASAP7_75t_L g11451 ( 
.A1(n_11250),
.A2(n_10733),
.B(n_10834),
.Y(n_11451)
);

AND2x4_ASAP7_75t_L g11452 ( 
.A(n_11101),
.B(n_10753),
.Y(n_11452)
);

AND2x2_ASAP7_75t_L g11453 ( 
.A(n_11186),
.B(n_11083),
.Y(n_11453)
);

OAI21x1_ASAP7_75t_L g11454 ( 
.A1(n_11265),
.A2(n_11079),
.B(n_10685),
.Y(n_11454)
);

OAI21x1_ASAP7_75t_L g11455 ( 
.A1(n_11288),
.A2(n_10873),
.B(n_10765),
.Y(n_11455)
);

OAI21x1_ASAP7_75t_L g11456 ( 
.A1(n_11318),
.A2(n_10684),
.B(n_10859),
.Y(n_11456)
);

NAND2xp5_ASAP7_75t_L g11457 ( 
.A(n_11427),
.B(n_10809),
.Y(n_11457)
);

NAND2x1p5_ASAP7_75t_L g11458 ( 
.A(n_11329),
.B(n_11030),
.Y(n_11458)
);

OA21x2_ASAP7_75t_L g11459 ( 
.A1(n_11319),
.A2(n_10871),
.B(n_10996),
.Y(n_11459)
);

AO21x2_ASAP7_75t_L g11460 ( 
.A1(n_11350),
.A2(n_10835),
.B(n_10970),
.Y(n_11460)
);

INVxp67_ASAP7_75t_SL g11461 ( 
.A(n_11263),
.Y(n_11461)
);

OAI21x1_ASAP7_75t_L g11462 ( 
.A1(n_11321),
.A2(n_10945),
.B(n_10937),
.Y(n_11462)
);

OAI21x1_ASAP7_75t_L g11463 ( 
.A1(n_11353),
.A2(n_10947),
.B(n_10983),
.Y(n_11463)
);

NOR2xp33_ASAP7_75t_R g11464 ( 
.A(n_11190),
.B(n_11093),
.Y(n_11464)
);

AO31x2_ASAP7_75t_L g11465 ( 
.A1(n_11366),
.A2(n_10810),
.A3(n_10936),
.B(n_10848),
.Y(n_11465)
);

HB1xp67_ASAP7_75t_L g11466 ( 
.A(n_11168),
.Y(n_11466)
);

AO21x2_ASAP7_75t_L g11467 ( 
.A1(n_11354),
.A2(n_10918),
.B(n_10879),
.Y(n_11467)
);

OAI21x1_ASAP7_75t_L g11468 ( 
.A1(n_11371),
.A2(n_11020),
.B(n_10736),
.Y(n_11468)
);

NAND3xp33_ASAP7_75t_L g11469 ( 
.A(n_11270),
.B(n_10693),
.C(n_10854),
.Y(n_11469)
);

INVx2_ASAP7_75t_L g11470 ( 
.A(n_11440),
.Y(n_11470)
);

INVx2_ASAP7_75t_L g11471 ( 
.A(n_11368),
.Y(n_11471)
);

OAI21x1_ASAP7_75t_L g11472 ( 
.A1(n_11372),
.A2(n_11374),
.B(n_11291),
.Y(n_11472)
);

INVx1_ASAP7_75t_L g11473 ( 
.A(n_11113),
.Y(n_11473)
);

AOI21xp5_ASAP7_75t_L g11474 ( 
.A1(n_11341),
.A2(n_11235),
.B(n_11299),
.Y(n_11474)
);

AO21x2_ASAP7_75t_L g11475 ( 
.A1(n_11264),
.A2(n_10725),
.B(n_10868),
.Y(n_11475)
);

AOI21xp5_ASAP7_75t_L g11476 ( 
.A1(n_11444),
.A2(n_10683),
.B(n_10863),
.Y(n_11476)
);

INVx1_ASAP7_75t_L g11477 ( 
.A(n_11416),
.Y(n_11477)
);

INVx2_ASAP7_75t_L g11478 ( 
.A(n_11370),
.Y(n_11478)
);

INVx3_ASAP7_75t_L g11479 ( 
.A(n_11106),
.Y(n_11479)
);

AND2x2_ASAP7_75t_L g11480 ( 
.A(n_11102),
.B(n_11104),
.Y(n_11480)
);

OA21x2_ASAP7_75t_L g11481 ( 
.A1(n_11328),
.A2(n_10928),
.B(n_11061),
.Y(n_11481)
);

NOR2xp33_ASAP7_75t_L g11482 ( 
.A(n_11326),
.B(n_10924),
.Y(n_11482)
);

AOI22xp33_ASAP7_75t_L g11483 ( 
.A1(n_11437),
.A2(n_11434),
.B1(n_11439),
.B2(n_11302),
.Y(n_11483)
);

OAI21x1_ASAP7_75t_L g11484 ( 
.A1(n_11281),
.A2(n_10902),
.B(n_10860),
.Y(n_11484)
);

NAND2x1p5_ASAP7_75t_L g11485 ( 
.A(n_11329),
.B(n_10951),
.Y(n_11485)
);

INVx2_ASAP7_75t_L g11486 ( 
.A(n_11111),
.Y(n_11486)
);

INVx2_ASAP7_75t_L g11487 ( 
.A(n_11359),
.Y(n_11487)
);

OAI21x1_ASAP7_75t_SL g11488 ( 
.A1(n_11205),
.A2(n_10759),
.B(n_10816),
.Y(n_11488)
);

NAND3xp33_ASAP7_75t_L g11489 ( 
.A(n_11171),
.B(n_11084),
.C(n_10732),
.Y(n_11489)
);

INVx1_ASAP7_75t_L g11490 ( 
.A(n_11121),
.Y(n_11490)
);

AO31x2_ASAP7_75t_L g11491 ( 
.A1(n_11405),
.A2(n_10723),
.A3(n_10905),
.B(n_10806),
.Y(n_11491)
);

OAI21x1_ASAP7_75t_L g11492 ( 
.A1(n_11404),
.A2(n_10934),
.B(n_10926),
.Y(n_11492)
);

CKINVDCx5p33_ASAP7_75t_R g11493 ( 
.A(n_11107),
.Y(n_11493)
);

OAI21xp5_ASAP7_75t_L g11494 ( 
.A1(n_11336),
.A2(n_10894),
.B(n_10825),
.Y(n_11494)
);

INVx2_ASAP7_75t_L g11495 ( 
.A(n_11369),
.Y(n_11495)
);

OAI21x1_ASAP7_75t_SL g11496 ( 
.A1(n_11196),
.A2(n_10828),
.B(n_10770),
.Y(n_11496)
);

OAI21x1_ASAP7_75t_L g11497 ( 
.A1(n_11406),
.A2(n_11409),
.B(n_11415),
.Y(n_11497)
);

NAND2xp5_ASAP7_75t_L g11498 ( 
.A(n_11389),
.B(n_11050),
.Y(n_11498)
);

HB1xp67_ASAP7_75t_L g11499 ( 
.A(n_11175),
.Y(n_11499)
);

INVx2_ASAP7_75t_L g11500 ( 
.A(n_11422),
.Y(n_11500)
);

INVx1_ASAP7_75t_L g11501 ( 
.A(n_11132),
.Y(n_11501)
);

NAND2xp5_ASAP7_75t_L g11502 ( 
.A(n_11392),
.B(n_10716),
.Y(n_11502)
);

OAI21x1_ASAP7_75t_L g11503 ( 
.A1(n_11379),
.A2(n_10862),
.B(n_11039),
.Y(n_11503)
);

OAI21x1_ASAP7_75t_L g11504 ( 
.A1(n_11387),
.A2(n_11068),
.B(n_10661),
.Y(n_11504)
);

INVx6_ASAP7_75t_L g11505 ( 
.A(n_11322),
.Y(n_11505)
);

BUFx8_ASAP7_75t_L g11506 ( 
.A(n_11118),
.Y(n_11506)
);

OAI21x1_ASAP7_75t_L g11507 ( 
.A1(n_11098),
.A2(n_10972),
.B(n_11036),
.Y(n_11507)
);

INVx1_ASAP7_75t_L g11508 ( 
.A(n_11135),
.Y(n_11508)
);

AOI21xp33_ASAP7_75t_SL g11509 ( 
.A1(n_11120),
.A2(n_11052),
.B(n_11054),
.Y(n_11509)
);

INVx1_ASAP7_75t_L g11510 ( 
.A(n_11167),
.Y(n_11510)
);

OA21x2_ASAP7_75t_L g11511 ( 
.A1(n_11339),
.A2(n_11034),
.B(n_10967),
.Y(n_11511)
);

OAI21x1_ASAP7_75t_L g11512 ( 
.A1(n_11096),
.A2(n_10925),
.B(n_10957),
.Y(n_11512)
);

INVx2_ASAP7_75t_L g11513 ( 
.A(n_11410),
.Y(n_11513)
);

NAND2xp5_ASAP7_75t_L g11514 ( 
.A(n_11088),
.B(n_10891),
.Y(n_11514)
);

OAI21x1_ASAP7_75t_L g11515 ( 
.A1(n_11097),
.A2(n_11047),
.B(n_10957),
.Y(n_11515)
);

OR2x2_ASAP7_75t_L g11516 ( 
.A(n_11092),
.B(n_10786),
.Y(n_11516)
);

BUFx3_ASAP7_75t_L g11517 ( 
.A(n_11194),
.Y(n_11517)
);

INVx1_ASAP7_75t_L g11518 ( 
.A(n_11179),
.Y(n_11518)
);

OAI21x1_ASAP7_75t_L g11519 ( 
.A1(n_11112),
.A2(n_11109),
.B(n_11105),
.Y(n_11519)
);

AO21x2_ASAP7_75t_L g11520 ( 
.A1(n_11130),
.A2(n_11244),
.B(n_11242),
.Y(n_11520)
);

INVx2_ASAP7_75t_L g11521 ( 
.A(n_11089),
.Y(n_11521)
);

AND2x4_ASAP7_75t_L g11522 ( 
.A(n_11156),
.B(n_10786),
.Y(n_11522)
);

OAI21x1_ASAP7_75t_L g11523 ( 
.A1(n_11099),
.A2(n_11047),
.B(n_11022),
.Y(n_11523)
);

OAI21x1_ASAP7_75t_L g11524 ( 
.A1(n_11139),
.A2(n_11110),
.B(n_11189),
.Y(n_11524)
);

INVx1_ASAP7_75t_L g11525 ( 
.A(n_11197),
.Y(n_11525)
);

OAI21x1_ASAP7_75t_L g11526 ( 
.A1(n_11203),
.A2(n_10959),
.B(n_1206),
.Y(n_11526)
);

INVx3_ASAP7_75t_L g11527 ( 
.A(n_11220),
.Y(n_11527)
);

OAI21x1_ASAP7_75t_L g11528 ( 
.A1(n_11221),
.A2(n_11237),
.B(n_11224),
.Y(n_11528)
);

OAI21x1_ASAP7_75t_L g11529 ( 
.A1(n_11248),
.A2(n_1207),
.B(n_1208),
.Y(n_11529)
);

NAND2xp5_ASAP7_75t_L g11530 ( 
.A(n_11349),
.B(n_1207),
.Y(n_11530)
);

BUFx3_ASAP7_75t_L g11531 ( 
.A(n_11254),
.Y(n_11531)
);

NAND2xp5_ASAP7_75t_L g11532 ( 
.A(n_11095),
.B(n_1207),
.Y(n_11532)
);

INVx2_ASAP7_75t_L g11533 ( 
.A(n_11115),
.Y(n_11533)
);

INVx4_ASAP7_75t_L g11534 ( 
.A(n_11136),
.Y(n_11534)
);

OA21x2_ASAP7_75t_L g11535 ( 
.A1(n_11253),
.A2(n_1208),
.B(n_1209),
.Y(n_11535)
);

OAI21x1_ASAP7_75t_L g11536 ( 
.A1(n_11296),
.A2(n_1208),
.B(n_1209),
.Y(n_11536)
);

NAND2xp5_ASAP7_75t_L g11537 ( 
.A(n_11420),
.B(n_1209),
.Y(n_11537)
);

BUFx3_ASAP7_75t_L g11538 ( 
.A(n_11103),
.Y(n_11538)
);

HB1xp67_ASAP7_75t_L g11539 ( 
.A(n_11435),
.Y(n_11539)
);

OAI21x1_ASAP7_75t_L g11540 ( 
.A1(n_11141),
.A2(n_1210),
.B(n_1211),
.Y(n_11540)
);

NAND2xp5_ASAP7_75t_L g11541 ( 
.A(n_11147),
.B(n_1211),
.Y(n_11541)
);

INVx1_ASAP7_75t_L g11542 ( 
.A(n_11172),
.Y(n_11542)
);

AND2x2_ASAP7_75t_L g11543 ( 
.A(n_11215),
.B(n_1211),
.Y(n_11543)
);

NAND2xp5_ASAP7_75t_L g11544 ( 
.A(n_11165),
.B(n_1212),
.Y(n_11544)
);

BUFx2_ASAP7_75t_L g11545 ( 
.A(n_11086),
.Y(n_11545)
);

AND2x2_ASAP7_75t_L g11546 ( 
.A(n_11309),
.B(n_1212),
.Y(n_11546)
);

OAI21x1_ASAP7_75t_L g11547 ( 
.A1(n_11273),
.A2(n_1212),
.B(n_1213),
.Y(n_11547)
);

OAI21x1_ASAP7_75t_L g11548 ( 
.A1(n_11401),
.A2(n_1213),
.B(n_1214),
.Y(n_11548)
);

BUFx3_ASAP7_75t_L g11549 ( 
.A(n_11240),
.Y(n_11549)
);

A2O1A1Ixp33_ASAP7_75t_L g11550 ( 
.A1(n_11269),
.A2(n_1215),
.B(n_1213),
.C(n_1214),
.Y(n_11550)
);

OAI21x1_ASAP7_75t_SL g11551 ( 
.A1(n_11133),
.A2(n_1214),
.B(n_1215),
.Y(n_11551)
);

OA21x2_ASAP7_75t_L g11552 ( 
.A1(n_11256),
.A2(n_1215),
.B(n_1216),
.Y(n_11552)
);

INVx2_ASAP7_75t_L g11553 ( 
.A(n_11164),
.Y(n_11553)
);

INVx1_ASAP7_75t_L g11554 ( 
.A(n_11181),
.Y(n_11554)
);

CKINVDCx11_ASAP7_75t_R g11555 ( 
.A(n_11293),
.Y(n_11555)
);

NAND2xp5_ASAP7_75t_L g11556 ( 
.A(n_11149),
.B(n_1216),
.Y(n_11556)
);

OAI21xp5_ASAP7_75t_L g11557 ( 
.A1(n_11356),
.A2(n_1217),
.B(n_1218),
.Y(n_11557)
);

OAI21x1_ASAP7_75t_L g11558 ( 
.A1(n_11268),
.A2(n_11262),
.B(n_11202),
.Y(n_11558)
);

OR2x2_ASAP7_75t_L g11559 ( 
.A(n_11324),
.B(n_1217),
.Y(n_11559)
);

HB1xp67_ASAP7_75t_L g11560 ( 
.A(n_11170),
.Y(n_11560)
);

OAI21x1_ASAP7_75t_L g11561 ( 
.A1(n_11183),
.A2(n_1218),
.B(n_1219),
.Y(n_11561)
);

OR2x2_ASAP7_75t_L g11562 ( 
.A(n_11315),
.B(n_1219),
.Y(n_11562)
);

INVx1_ASAP7_75t_L g11563 ( 
.A(n_11204),
.Y(n_11563)
);

INVx1_ASAP7_75t_L g11564 ( 
.A(n_11214),
.Y(n_11564)
);

AOI21xp5_ASAP7_75t_L g11565 ( 
.A1(n_11425),
.A2(n_1220),
.B(n_1221),
.Y(n_11565)
);

INVx2_ASAP7_75t_L g11566 ( 
.A(n_11234),
.Y(n_11566)
);

INVx1_ASAP7_75t_L g11567 ( 
.A(n_11261),
.Y(n_11567)
);

OAI21x1_ASAP7_75t_L g11568 ( 
.A1(n_11323),
.A2(n_1220),
.B(n_1221),
.Y(n_11568)
);

AND2x2_ASAP7_75t_L g11569 ( 
.A(n_11162),
.B(n_1220),
.Y(n_11569)
);

CKINVDCx5p33_ASAP7_75t_R g11570 ( 
.A(n_11312),
.Y(n_11570)
);

HB1xp67_ASAP7_75t_L g11571 ( 
.A(n_11217),
.Y(n_11571)
);

AND2x4_ASAP7_75t_L g11572 ( 
.A(n_11146),
.B(n_1222),
.Y(n_11572)
);

AND2x4_ASAP7_75t_L g11573 ( 
.A(n_11247),
.B(n_1223),
.Y(n_11573)
);

INVxp67_ASAP7_75t_L g11574 ( 
.A(n_11266),
.Y(n_11574)
);

INVxp67_ASAP7_75t_SL g11575 ( 
.A(n_11198),
.Y(n_11575)
);

OAI21xp5_ASAP7_75t_L g11576 ( 
.A1(n_11127),
.A2(n_1223),
.B(n_1224),
.Y(n_11576)
);

OAI21x1_ASAP7_75t_L g11577 ( 
.A1(n_11304),
.A2(n_11151),
.B(n_11150),
.Y(n_11577)
);

NAND2xp5_ASAP7_75t_SL g11578 ( 
.A(n_11162),
.B(n_1223),
.Y(n_11578)
);

NAND2xp5_ASAP7_75t_L g11579 ( 
.A(n_11199),
.B(n_1224),
.Y(n_11579)
);

INVx1_ASAP7_75t_L g11580 ( 
.A(n_11129),
.Y(n_11580)
);

AO21x2_ASAP7_75t_L g11581 ( 
.A1(n_11182),
.A2(n_1224),
.B(n_1225),
.Y(n_11581)
);

OA21x2_ASAP7_75t_L g11582 ( 
.A1(n_11236),
.A2(n_1226),
.B(n_1227),
.Y(n_11582)
);

INVx1_ASAP7_75t_L g11583 ( 
.A(n_11201),
.Y(n_11583)
);

OAI21x1_ASAP7_75t_L g11584 ( 
.A1(n_11145),
.A2(n_1226),
.B(n_1227),
.Y(n_11584)
);

INVx2_ASAP7_75t_L g11585 ( 
.A(n_11388),
.Y(n_11585)
);

AO21x2_ASAP7_75t_L g11586 ( 
.A1(n_11143),
.A2(n_1226),
.B(n_1227),
.Y(n_11586)
);

AO21x2_ASAP7_75t_L g11587 ( 
.A1(n_11282),
.A2(n_1228),
.B(n_1229),
.Y(n_11587)
);

OAI21x1_ASAP7_75t_L g11588 ( 
.A1(n_11134),
.A2(n_1228),
.B(n_1229),
.Y(n_11588)
);

INVx2_ASAP7_75t_SL g11589 ( 
.A(n_11163),
.Y(n_11589)
);

INVx2_ASAP7_75t_L g11590 ( 
.A(n_11258),
.Y(n_11590)
);

INVx2_ASAP7_75t_L g11591 ( 
.A(n_11352),
.Y(n_11591)
);

AO31x2_ASAP7_75t_L g11592 ( 
.A1(n_11123),
.A2(n_11218),
.A3(n_11364),
.B(n_11432),
.Y(n_11592)
);

INVx3_ASAP7_75t_L g11593 ( 
.A(n_11345),
.Y(n_11593)
);

INVx1_ASAP7_75t_L g11594 ( 
.A(n_11148),
.Y(n_11594)
);

INVx1_ASAP7_75t_L g11595 ( 
.A(n_11148),
.Y(n_11595)
);

A2O1A1Ixp33_ASAP7_75t_L g11596 ( 
.A1(n_11373),
.A2(n_1232),
.B(n_1230),
.C(n_1231),
.Y(n_11596)
);

AOI21xp5_ASAP7_75t_L g11597 ( 
.A1(n_11267),
.A2(n_2450),
.B(n_2449),
.Y(n_11597)
);

AO21x2_ASAP7_75t_L g11598 ( 
.A1(n_11206),
.A2(n_1231),
.B(n_1232),
.Y(n_11598)
);

NOR2xp33_ASAP7_75t_SL g11599 ( 
.A(n_11138),
.B(n_1233),
.Y(n_11599)
);

A2O1A1Ixp33_ASAP7_75t_L g11600 ( 
.A1(n_11418),
.A2(n_1235),
.B(n_1233),
.C(n_1234),
.Y(n_11600)
);

INVx2_ASAP7_75t_L g11601 ( 
.A(n_11386),
.Y(n_11601)
);

NAND2x1p5_ASAP7_75t_L g11602 ( 
.A(n_11142),
.B(n_1234),
.Y(n_11602)
);

AND2x2_ASAP7_75t_L g11603 ( 
.A(n_11162),
.B(n_1234),
.Y(n_11603)
);

NAND2xp5_ASAP7_75t_L g11604 ( 
.A(n_11274),
.B(n_1235),
.Y(n_11604)
);

NOR2xp33_ASAP7_75t_L g11605 ( 
.A(n_11090),
.B(n_1236),
.Y(n_11605)
);

BUFx12f_ASAP7_75t_L g11606 ( 
.A(n_11157),
.Y(n_11606)
);

INVx1_ASAP7_75t_L g11607 ( 
.A(n_11114),
.Y(n_11607)
);

BUFx2_ASAP7_75t_L g11608 ( 
.A(n_11230),
.Y(n_11608)
);

OAI21x1_ASAP7_75t_L g11609 ( 
.A1(n_11154),
.A2(n_11122),
.B(n_11117),
.Y(n_11609)
);

BUFx3_ASAP7_75t_L g11610 ( 
.A(n_11124),
.Y(n_11610)
);

AND2x2_ASAP7_75t_L g11611 ( 
.A(n_11311),
.B(n_1236),
.Y(n_11611)
);

AND2x2_ASAP7_75t_L g11612 ( 
.A(n_11292),
.B(n_1236),
.Y(n_11612)
);

NOR2xp33_ASAP7_75t_L g11613 ( 
.A(n_11108),
.B(n_2438),
.Y(n_11613)
);

INVx1_ASAP7_75t_L g11614 ( 
.A(n_11287),
.Y(n_11614)
);

AND2x4_ASAP7_75t_L g11615 ( 
.A(n_11187),
.B(n_1237),
.Y(n_11615)
);

OAI21x1_ASAP7_75t_L g11616 ( 
.A1(n_11128),
.A2(n_1237),
.B(n_1238),
.Y(n_11616)
);

INVxp67_ASAP7_75t_SL g11617 ( 
.A(n_11342),
.Y(n_11617)
);

OAI21x1_ASAP7_75t_L g11618 ( 
.A1(n_11169),
.A2(n_1238),
.B(n_1239),
.Y(n_11618)
);

INVx2_ASAP7_75t_L g11619 ( 
.A(n_11347),
.Y(n_11619)
);

AOI21x1_ASAP7_75t_L g11620 ( 
.A1(n_11119),
.A2(n_1238),
.B(n_1239),
.Y(n_11620)
);

NOR2xp33_ASAP7_75t_L g11621 ( 
.A(n_11313),
.B(n_2440),
.Y(n_11621)
);

AOI21x1_ASAP7_75t_L g11622 ( 
.A1(n_11188),
.A2(n_1239),
.B(n_1240),
.Y(n_11622)
);

OAI21x1_ASAP7_75t_L g11623 ( 
.A1(n_11178),
.A2(n_1240),
.B(n_1241),
.Y(n_11623)
);

OAI21x1_ASAP7_75t_L g11624 ( 
.A1(n_11338),
.A2(n_1240),
.B(n_1241),
.Y(n_11624)
);

CKINVDCx14_ASAP7_75t_R g11625 ( 
.A(n_11283),
.Y(n_11625)
);

AND2x2_ASAP7_75t_L g11626 ( 
.A(n_11192),
.B(n_1242),
.Y(n_11626)
);

INVx2_ASAP7_75t_L g11627 ( 
.A(n_11320),
.Y(n_11627)
);

AND2x2_ASAP7_75t_L g11628 ( 
.A(n_11277),
.B(n_1243),
.Y(n_11628)
);

AOI22xp33_ASAP7_75t_L g11629 ( 
.A1(n_11208),
.A2(n_1245),
.B1(n_1243),
.B2(n_1244),
.Y(n_11629)
);

NAND2x1p5_ASAP7_75t_L g11630 ( 
.A(n_11308),
.B(n_11272),
.Y(n_11630)
);

BUFx3_ASAP7_75t_L g11631 ( 
.A(n_11140),
.Y(n_11631)
);

CKINVDCx20_ASAP7_75t_R g11632 ( 
.A(n_11307),
.Y(n_11632)
);

AO31x2_ASAP7_75t_L g11633 ( 
.A1(n_11259),
.A2(n_11125),
.A3(n_11126),
.B(n_11424),
.Y(n_11633)
);

OAI21x1_ASAP7_75t_L g11634 ( 
.A1(n_11412),
.A2(n_1244),
.B(n_1245),
.Y(n_11634)
);

OAI21xp5_ASAP7_75t_L g11635 ( 
.A1(n_11131),
.A2(n_1244),
.B(n_1245),
.Y(n_11635)
);

BUFx3_ASAP7_75t_L g11636 ( 
.A(n_11362),
.Y(n_11636)
);

INVx2_ASAP7_75t_L g11637 ( 
.A(n_11091),
.Y(n_11637)
);

OAI21x1_ASAP7_75t_L g11638 ( 
.A1(n_11209),
.A2(n_1246),
.B(n_1247),
.Y(n_11638)
);

AOI21xp5_ASAP7_75t_L g11639 ( 
.A1(n_11396),
.A2(n_11233),
.B(n_11433),
.Y(n_11639)
);

AOI21xp5_ASAP7_75t_L g11640 ( 
.A1(n_11255),
.A2(n_11297),
.B(n_11276),
.Y(n_11640)
);

INVx2_ASAP7_75t_SL g11641 ( 
.A(n_11238),
.Y(n_11641)
);

AOI21xp33_ASAP7_75t_SL g11642 ( 
.A1(n_11337),
.A2(n_1246),
.B(n_1247),
.Y(n_11642)
);

BUFx12f_ASAP7_75t_L g11643 ( 
.A(n_11367),
.Y(n_11643)
);

INVx2_ASAP7_75t_L g11644 ( 
.A(n_11344),
.Y(n_11644)
);

INVx2_ASAP7_75t_L g11645 ( 
.A(n_11351),
.Y(n_11645)
);

INVx5_ASAP7_75t_L g11646 ( 
.A(n_11286),
.Y(n_11646)
);

INVx1_ASAP7_75t_L g11647 ( 
.A(n_11346),
.Y(n_11647)
);

OAI21x1_ASAP7_75t_L g11648 ( 
.A1(n_11219),
.A2(n_1247),
.B(n_1248),
.Y(n_11648)
);

BUFx6f_ASAP7_75t_L g11649 ( 
.A(n_11200),
.Y(n_11649)
);

OA21x2_ASAP7_75t_L g11650 ( 
.A1(n_11303),
.A2(n_1248),
.B(n_1249),
.Y(n_11650)
);

INVx1_ASAP7_75t_L g11651 ( 
.A(n_11363),
.Y(n_11651)
);

INVx1_ASAP7_75t_L g11652 ( 
.A(n_11381),
.Y(n_11652)
);

AO31x2_ASAP7_75t_L g11653 ( 
.A1(n_11153),
.A2(n_1250),
.A3(n_1248),
.B(n_1249),
.Y(n_11653)
);

OAI21x1_ASAP7_75t_L g11654 ( 
.A1(n_11279),
.A2(n_1250),
.B(n_1251),
.Y(n_11654)
);

OA21x2_ASAP7_75t_L g11655 ( 
.A1(n_11411),
.A2(n_1250),
.B(n_1251),
.Y(n_11655)
);

INVx1_ASAP7_75t_L g11656 ( 
.A(n_11394),
.Y(n_11656)
);

HB1xp67_ASAP7_75t_L g11657 ( 
.A(n_11100),
.Y(n_11657)
);

INVx2_ASAP7_75t_L g11658 ( 
.A(n_11166),
.Y(n_11658)
);

AO21x1_ASAP7_75t_L g11659 ( 
.A1(n_11327),
.A2(n_1251),
.B(n_1252),
.Y(n_11659)
);

INVx1_ASAP7_75t_L g11660 ( 
.A(n_11100),
.Y(n_11660)
);

NOR2xp33_ASAP7_75t_SL g11661 ( 
.A(n_11393),
.B(n_1252),
.Y(n_11661)
);

INVx2_ASAP7_75t_L g11662 ( 
.A(n_11284),
.Y(n_11662)
);

AOI21xp5_ASAP7_75t_L g11663 ( 
.A1(n_11443),
.A2(n_2439),
.B(n_2438),
.Y(n_11663)
);

AO31x2_ASAP7_75t_L g11664 ( 
.A1(n_11331),
.A2(n_1254),
.A3(n_1252),
.B(n_1253),
.Y(n_11664)
);

OAI21x1_ASAP7_75t_L g11665 ( 
.A1(n_11152),
.A2(n_1253),
.B(n_1254),
.Y(n_11665)
);

OAI21x1_ASAP7_75t_L g11666 ( 
.A1(n_11295),
.A2(n_1253),
.B(n_1255),
.Y(n_11666)
);

OAI21x1_ASAP7_75t_L g11667 ( 
.A1(n_11161),
.A2(n_1255),
.B(n_1257),
.Y(n_11667)
);

INVx1_ASAP7_75t_L g11668 ( 
.A(n_11275),
.Y(n_11668)
);

OAI21x1_ASAP7_75t_L g11669 ( 
.A1(n_11300),
.A2(n_11185),
.B(n_11180),
.Y(n_11669)
);

OR2x6_ASAP7_75t_L g11670 ( 
.A(n_11116),
.B(n_1255),
.Y(n_11670)
);

INVx2_ASAP7_75t_L g11671 ( 
.A(n_11174),
.Y(n_11671)
);

OR2x6_ASAP7_75t_L g11672 ( 
.A(n_11137),
.B(n_1257),
.Y(n_11672)
);

OAI21x1_ASAP7_75t_L g11673 ( 
.A1(n_11316),
.A2(n_1257),
.B(n_1258),
.Y(n_11673)
);

BUFx6f_ASAP7_75t_L g11674 ( 
.A(n_11231),
.Y(n_11674)
);

INVx3_ASAP7_75t_L g11675 ( 
.A(n_11195),
.Y(n_11675)
);

HB1xp67_ASAP7_75t_L g11676 ( 
.A(n_11294),
.Y(n_11676)
);

INVx4_ASAP7_75t_SL g11677 ( 
.A(n_11211),
.Y(n_11677)
);

NAND2xp5_ASAP7_75t_L g11678 ( 
.A(n_11225),
.B(n_1258),
.Y(n_11678)
);

NAND2xp5_ASAP7_75t_L g11679 ( 
.A(n_11232),
.B(n_11245),
.Y(n_11679)
);

INVxp67_ASAP7_75t_L g11680 ( 
.A(n_11310),
.Y(n_11680)
);

INVx1_ASAP7_75t_SL g11681 ( 
.A(n_11210),
.Y(n_11681)
);

HB1xp67_ASAP7_75t_L g11682 ( 
.A(n_11317),
.Y(n_11682)
);

OA21x2_ASAP7_75t_L g11683 ( 
.A1(n_11343),
.A2(n_1258),
.B(n_1259),
.Y(n_11683)
);

NAND2xp5_ASAP7_75t_L g11684 ( 
.A(n_11252),
.B(n_1259),
.Y(n_11684)
);

BUFx6f_ASAP7_75t_L g11685 ( 
.A(n_11251),
.Y(n_11685)
);

AND2x2_ASAP7_75t_L g11686 ( 
.A(n_11193),
.B(n_1260),
.Y(n_11686)
);

INVx1_ASAP7_75t_L g11687 ( 
.A(n_11246),
.Y(n_11687)
);

OA21x2_ASAP7_75t_L g11688 ( 
.A1(n_11357),
.A2(n_1260),
.B(n_1261),
.Y(n_11688)
);

NAND2xp5_ASAP7_75t_L g11689 ( 
.A(n_11278),
.B(n_1260),
.Y(n_11689)
);

INVx3_ASAP7_75t_L g11690 ( 
.A(n_11280),
.Y(n_11690)
);

INVx1_ASAP7_75t_L g11691 ( 
.A(n_11332),
.Y(n_11691)
);

INVx6_ASAP7_75t_L g11692 ( 
.A(n_11335),
.Y(n_11692)
);

OAI21x1_ASAP7_75t_L g11693 ( 
.A1(n_11383),
.A2(n_1261),
.B(n_1262),
.Y(n_11693)
);

INVx3_ASAP7_75t_L g11694 ( 
.A(n_11398),
.Y(n_11694)
);

OAI21x1_ASAP7_75t_L g11695 ( 
.A1(n_11384),
.A2(n_1262),
.B(n_1263),
.Y(n_11695)
);

OR2x2_ASAP7_75t_L g11696 ( 
.A(n_11332),
.B(n_1262),
.Y(n_11696)
);

OAI21xp5_ASAP7_75t_L g11697 ( 
.A1(n_11243),
.A2(n_1263),
.B(n_1264),
.Y(n_11697)
);

OA21x2_ASAP7_75t_L g11698 ( 
.A1(n_11223),
.A2(n_1263),
.B(n_1264),
.Y(n_11698)
);

AOI21x1_ASAP7_75t_L g11699 ( 
.A1(n_11213),
.A2(n_1264),
.B(n_1265),
.Y(n_11699)
);

OA21x2_ASAP7_75t_L g11700 ( 
.A1(n_11333),
.A2(n_1265),
.B(n_1266),
.Y(n_11700)
);

OA21x2_ASAP7_75t_L g11701 ( 
.A1(n_11358),
.A2(n_1266),
.B(n_1267),
.Y(n_11701)
);

INVx1_ASAP7_75t_L g11702 ( 
.A(n_11414),
.Y(n_11702)
);

AOI21xp5_ASAP7_75t_L g11703 ( 
.A1(n_11400),
.A2(n_1268),
.B(n_1269),
.Y(n_11703)
);

INVx1_ASAP7_75t_L g11704 ( 
.A(n_11226),
.Y(n_11704)
);

INVx2_ASAP7_75t_L g11705 ( 
.A(n_11407),
.Y(n_11705)
);

BUFx6f_ASAP7_75t_L g11706 ( 
.A(n_11334),
.Y(n_11706)
);

AO31x2_ASAP7_75t_L g11707 ( 
.A1(n_11305),
.A2(n_1272),
.A3(n_1270),
.B(n_1271),
.Y(n_11707)
);

AND2x4_ASAP7_75t_L g11708 ( 
.A(n_11085),
.B(n_1270),
.Y(n_11708)
);

INVx6_ASAP7_75t_L g11709 ( 
.A(n_11239),
.Y(n_11709)
);

NOR2x1_ASAP7_75t_SL g11710 ( 
.A(n_11431),
.B(n_1270),
.Y(n_11710)
);

INVx1_ASAP7_75t_L g11711 ( 
.A(n_11227),
.Y(n_11711)
);

OA21x2_ASAP7_75t_L g11712 ( 
.A1(n_11228),
.A2(n_1271),
.B(n_1272),
.Y(n_11712)
);

NOR2x1_ASAP7_75t_SL g11713 ( 
.A(n_11397),
.B(n_1271),
.Y(n_11713)
);

AND2x2_ASAP7_75t_L g11714 ( 
.A(n_11399),
.B(n_1272),
.Y(n_11714)
);

NOR2x1_ASAP7_75t_SL g11715 ( 
.A(n_11173),
.B(n_1273),
.Y(n_11715)
);

NAND2xp5_ASAP7_75t_SL g11716 ( 
.A(n_11348),
.B(n_1273),
.Y(n_11716)
);

OAI21x1_ASAP7_75t_L g11717 ( 
.A1(n_11144),
.A2(n_1273),
.B(n_1275),
.Y(n_11717)
);

OAI21x1_ASAP7_75t_L g11718 ( 
.A1(n_11212),
.A2(n_1275),
.B(n_1276),
.Y(n_11718)
);

AO21x2_ASAP7_75t_L g11719 ( 
.A1(n_11177),
.A2(n_1276),
.B(n_1277),
.Y(n_11719)
);

INVx1_ASAP7_75t_L g11720 ( 
.A(n_11241),
.Y(n_11720)
);

OAI21x1_ASAP7_75t_L g11721 ( 
.A1(n_11260),
.A2(n_11271),
.B(n_11216),
.Y(n_11721)
);

OAI21x1_ASAP7_75t_L g11722 ( 
.A1(n_11207),
.A2(n_1277),
.B(n_1278),
.Y(n_11722)
);

OR2x6_ASAP7_75t_L g11723 ( 
.A(n_11155),
.B(n_1278),
.Y(n_11723)
);

OAI21xp5_ASAP7_75t_L g11724 ( 
.A1(n_11375),
.A2(n_1278),
.B(n_1279),
.Y(n_11724)
);

OAI21x1_ASAP7_75t_L g11725 ( 
.A1(n_11159),
.A2(n_1279),
.B(n_1280),
.Y(n_11725)
);

AND2x2_ASAP7_75t_L g11726 ( 
.A(n_11191),
.B(n_1279),
.Y(n_11726)
);

INVx1_ASAP7_75t_L g11727 ( 
.A(n_11085),
.Y(n_11727)
);

OAI21x1_ASAP7_75t_L g11728 ( 
.A1(n_11222),
.A2(n_1280),
.B(n_1281),
.Y(n_11728)
);

INVx2_ASAP7_75t_L g11729 ( 
.A(n_11421),
.Y(n_11729)
);

INVx2_ASAP7_75t_L g11730 ( 
.A(n_11360),
.Y(n_11730)
);

OAI21x1_ASAP7_75t_L g11731 ( 
.A1(n_11184),
.A2(n_1281),
.B(n_1282),
.Y(n_11731)
);

INVx1_ASAP7_75t_L g11732 ( 
.A(n_11325),
.Y(n_11732)
);

NAND2xp5_ASAP7_75t_L g11733 ( 
.A(n_11441),
.B(n_1281),
.Y(n_11733)
);

HB1xp67_ASAP7_75t_L g11734 ( 
.A(n_11417),
.Y(n_11734)
);

INVx1_ASAP7_75t_L g11735 ( 
.A(n_11330),
.Y(n_11735)
);

AOI21xp5_ASAP7_75t_L g11736 ( 
.A1(n_11413),
.A2(n_2452),
.B(n_2451),
.Y(n_11736)
);

OA21x2_ASAP7_75t_L g11737 ( 
.A1(n_11290),
.A2(n_1282),
.B(n_1284),
.Y(n_11737)
);

OR2x6_ASAP7_75t_L g11738 ( 
.A(n_11160),
.B(n_1282),
.Y(n_11738)
);

BUFx2_ASAP7_75t_R g11739 ( 
.A(n_11402),
.Y(n_11739)
);

INVxp67_ASAP7_75t_SL g11740 ( 
.A(n_11408),
.Y(n_11740)
);

INVxp67_ASAP7_75t_L g11741 ( 
.A(n_11211),
.Y(n_11741)
);

OAI21x1_ASAP7_75t_L g11742 ( 
.A1(n_11298),
.A2(n_1284),
.B(n_1285),
.Y(n_11742)
);

AOI21xp5_ASAP7_75t_L g11743 ( 
.A1(n_11289),
.A2(n_1286),
.B(n_1287),
.Y(n_11743)
);

AOI22xp5_ASAP7_75t_L g11744 ( 
.A1(n_11445),
.A2(n_1288),
.B1(n_1286),
.B2(n_1287),
.Y(n_11744)
);

BUFx3_ASAP7_75t_L g11745 ( 
.A(n_11419),
.Y(n_11745)
);

OAI21xp5_ASAP7_75t_L g11746 ( 
.A1(n_11390),
.A2(n_1286),
.B(n_1288),
.Y(n_11746)
);

AND2x4_ASAP7_75t_L g11747 ( 
.A(n_11355),
.B(n_1288),
.Y(n_11747)
);

INVx6_ASAP7_75t_L g11748 ( 
.A(n_11423),
.Y(n_11748)
);

OA21x2_ASAP7_75t_L g11749 ( 
.A1(n_11306),
.A2(n_1289),
.B(n_1290),
.Y(n_11749)
);

INVx1_ASAP7_75t_L g11750 ( 
.A(n_11314),
.Y(n_11750)
);

AND2x4_ASAP7_75t_L g11751 ( 
.A(n_11361),
.B(n_1290),
.Y(n_11751)
);

A2O1A1Ixp33_ASAP7_75t_L g11752 ( 
.A1(n_11429),
.A2(n_11438),
.B(n_11430),
.C(n_11436),
.Y(n_11752)
);

INVx1_ASAP7_75t_L g11753 ( 
.A(n_11403),
.Y(n_11753)
);

OAI21xp5_ASAP7_75t_L g11754 ( 
.A1(n_11426),
.A2(n_1290),
.B(n_1291),
.Y(n_11754)
);

OAI21x1_ASAP7_75t_L g11755 ( 
.A1(n_11340),
.A2(n_1291),
.B(n_1292),
.Y(n_11755)
);

AO31x2_ASAP7_75t_L g11756 ( 
.A1(n_11428),
.A2(n_1293),
.A3(n_1291),
.B(n_1292),
.Y(n_11756)
);

OAI21x1_ASAP7_75t_L g11757 ( 
.A1(n_11380),
.A2(n_1293),
.B(n_1294),
.Y(n_11757)
);

INVx2_ASAP7_75t_L g11758 ( 
.A(n_11382),
.Y(n_11758)
);

BUFx2_ASAP7_75t_L g11759 ( 
.A(n_11365),
.Y(n_11759)
);

INVx1_ASAP7_75t_L g11760 ( 
.A(n_11376),
.Y(n_11760)
);

INVx2_ASAP7_75t_L g11761 ( 
.A(n_11377),
.Y(n_11761)
);

OAI21x1_ASAP7_75t_SL g11762 ( 
.A1(n_11229),
.A2(n_1293),
.B(n_1294),
.Y(n_11762)
);

AND2x2_ASAP7_75t_L g11763 ( 
.A(n_11378),
.B(n_1295),
.Y(n_11763)
);

NOR2xp33_ASAP7_75t_L g11764 ( 
.A(n_11257),
.B(n_2446),
.Y(n_11764)
);

OAI21x1_ASAP7_75t_L g11765 ( 
.A1(n_11385),
.A2(n_1295),
.B(n_1296),
.Y(n_11765)
);

OAI21x1_ASAP7_75t_L g11766 ( 
.A1(n_11391),
.A2(n_1295),
.B(n_1296),
.Y(n_11766)
);

AO21x2_ASAP7_75t_L g11767 ( 
.A1(n_11395),
.A2(n_11249),
.B(n_11285),
.Y(n_11767)
);

OAI21x1_ASAP7_75t_L g11768 ( 
.A1(n_11442),
.A2(n_1296),
.B(n_1297),
.Y(n_11768)
);

NOR2xp33_ASAP7_75t_L g11769 ( 
.A(n_11326),
.B(n_2449),
.Y(n_11769)
);

NAND2xp5_ASAP7_75t_L g11770 ( 
.A(n_11427),
.B(n_1297),
.Y(n_11770)
);

AOI21xp5_ASAP7_75t_L g11771 ( 
.A1(n_11427),
.A2(n_2451),
.B(n_2450),
.Y(n_11771)
);

AO31x2_ASAP7_75t_L g11772 ( 
.A1(n_11427),
.A2(n_1299),
.A3(n_1297),
.B(n_1298),
.Y(n_11772)
);

AOI21xp5_ASAP7_75t_L g11773 ( 
.A1(n_11427),
.A2(n_2452),
.B(n_1298),
.Y(n_11773)
);

NAND2x1p5_ASAP7_75t_L g11774 ( 
.A(n_11329),
.B(n_1298),
.Y(n_11774)
);

INVx3_ASAP7_75t_L g11775 ( 
.A(n_11106),
.Y(n_11775)
);

NAND2xp5_ASAP7_75t_L g11776 ( 
.A(n_11427),
.B(n_1299),
.Y(n_11776)
);

AO31x2_ASAP7_75t_L g11777 ( 
.A1(n_11427),
.A2(n_1301),
.A3(n_1299),
.B(n_1300),
.Y(n_11777)
);

OR2x2_ASAP7_75t_L g11778 ( 
.A(n_11113),
.B(n_1300),
.Y(n_11778)
);

OAI21x1_ASAP7_75t_L g11779 ( 
.A1(n_11301),
.A2(n_1300),
.B(n_1301),
.Y(n_11779)
);

NOR2x1_ASAP7_75t_SL g11780 ( 
.A(n_11329),
.B(n_1302),
.Y(n_11780)
);

AOI21x1_ASAP7_75t_L g11781 ( 
.A1(n_11319),
.A2(n_1302),
.B(n_1303),
.Y(n_11781)
);

INVx1_ASAP7_75t_L g11782 ( 
.A(n_11087),
.Y(n_11782)
);

INVx1_ASAP7_75t_L g11783 ( 
.A(n_11087),
.Y(n_11783)
);

CKINVDCx5p33_ASAP7_75t_R g11784 ( 
.A(n_11093),
.Y(n_11784)
);

OAI21x1_ASAP7_75t_L g11785 ( 
.A1(n_11301),
.A2(n_1302),
.B(n_1303),
.Y(n_11785)
);

NAND2xp5_ASAP7_75t_SL g11786 ( 
.A(n_11319),
.B(n_1304),
.Y(n_11786)
);

INVx4_ASAP7_75t_SL g11787 ( 
.A(n_11240),
.Y(n_11787)
);

OA21x2_ASAP7_75t_L g11788 ( 
.A1(n_11319),
.A2(n_1304),
.B(n_1305),
.Y(n_11788)
);

OA21x2_ASAP7_75t_L g11789 ( 
.A1(n_11319),
.A2(n_1304),
.B(n_1305),
.Y(n_11789)
);

OAI21x1_ASAP7_75t_L g11790 ( 
.A1(n_11301),
.A2(n_1306),
.B(n_1307),
.Y(n_11790)
);

AO21x2_ASAP7_75t_L g11791 ( 
.A1(n_11265),
.A2(n_1306),
.B(n_1308),
.Y(n_11791)
);

NAND2x1p5_ASAP7_75t_L g11792 ( 
.A(n_11329),
.B(n_1308),
.Y(n_11792)
);

AOI21xp5_ASAP7_75t_L g11793 ( 
.A1(n_11427),
.A2(n_2447),
.B(n_2445),
.Y(n_11793)
);

INVx1_ASAP7_75t_SL g11794 ( 
.A(n_11086),
.Y(n_11794)
);

AOI21x1_ASAP7_75t_L g11795 ( 
.A1(n_11319),
.A2(n_1309),
.B(n_1310),
.Y(n_11795)
);

NAND2xp5_ASAP7_75t_L g11796 ( 
.A(n_11427),
.B(n_1309),
.Y(n_11796)
);

BUFx2_ASAP7_75t_L g11797 ( 
.A(n_11086),
.Y(n_11797)
);

AOI22x1_ASAP7_75t_L g11798 ( 
.A1(n_11427),
.A2(n_1311),
.B1(n_1309),
.B2(n_1310),
.Y(n_11798)
);

NAND2xp5_ASAP7_75t_L g11799 ( 
.A(n_11427),
.B(n_1310),
.Y(n_11799)
);

INVx2_ASAP7_75t_L g11800 ( 
.A(n_11168),
.Y(n_11800)
);

AOI21x1_ASAP7_75t_L g11801 ( 
.A1(n_11319),
.A2(n_1311),
.B(n_1312),
.Y(n_11801)
);

INVx2_ASAP7_75t_L g11802 ( 
.A(n_11168),
.Y(n_11802)
);

BUFx2_ASAP7_75t_L g11803 ( 
.A(n_11086),
.Y(n_11803)
);

OR2x6_ASAP7_75t_L g11804 ( 
.A(n_11124),
.B(n_1312),
.Y(n_11804)
);

OA21x2_ASAP7_75t_L g11805 ( 
.A1(n_11319),
.A2(n_1313),
.B(n_1314),
.Y(n_11805)
);

OAI21x1_ASAP7_75t_L g11806 ( 
.A1(n_11301),
.A2(n_1313),
.B(n_1314),
.Y(n_11806)
);

INVx2_ASAP7_75t_L g11807 ( 
.A(n_11168),
.Y(n_11807)
);

INVx3_ASAP7_75t_L g11808 ( 
.A(n_11106),
.Y(n_11808)
);

NOR2x1_ASAP7_75t_SL g11809 ( 
.A(n_11329),
.B(n_1315),
.Y(n_11809)
);

HB1xp67_ASAP7_75t_L g11810 ( 
.A(n_11168),
.Y(n_11810)
);

BUFx2_ASAP7_75t_L g11811 ( 
.A(n_11086),
.Y(n_11811)
);

INVx1_ASAP7_75t_L g11812 ( 
.A(n_11087),
.Y(n_11812)
);

BUFx6f_ASAP7_75t_L g11813 ( 
.A(n_11106),
.Y(n_11813)
);

NAND2xp5_ASAP7_75t_L g11814 ( 
.A(n_11427),
.B(n_1315),
.Y(n_11814)
);

OAI21x1_ASAP7_75t_L g11815 ( 
.A1(n_11301),
.A2(n_1315),
.B(n_1316),
.Y(n_11815)
);

NOR2xp33_ASAP7_75t_L g11816 ( 
.A(n_11326),
.B(n_1316),
.Y(n_11816)
);

AOI21xp5_ASAP7_75t_L g11817 ( 
.A1(n_11427),
.A2(n_2437),
.B(n_2436),
.Y(n_11817)
);

INVx2_ASAP7_75t_L g11818 ( 
.A(n_11168),
.Y(n_11818)
);

BUFx3_ASAP7_75t_L g11819 ( 
.A(n_11632),
.Y(n_11819)
);

AND2x2_ASAP7_75t_L g11820 ( 
.A(n_11545),
.B(n_1317),
.Y(n_11820)
);

NOR2xp67_ASAP7_75t_L g11821 ( 
.A(n_11574),
.B(n_1317),
.Y(n_11821)
);

NAND2xp5_ASAP7_75t_L g11822 ( 
.A(n_11614),
.B(n_1318),
.Y(n_11822)
);

AND2x2_ASAP7_75t_L g11823 ( 
.A(n_11797),
.B(n_11803),
.Y(n_11823)
);

AND2x2_ASAP7_75t_L g11824 ( 
.A(n_11811),
.B(n_1318),
.Y(n_11824)
);

HB1xp67_ASAP7_75t_L g11825 ( 
.A(n_11607),
.Y(n_11825)
);

AND2x4_ASAP7_75t_L g11826 ( 
.A(n_11617),
.B(n_1318),
.Y(n_11826)
);

AOI21x1_ASAP7_75t_SL g11827 ( 
.A1(n_11457),
.A2(n_1319),
.B(n_1320),
.Y(n_11827)
);

OAI22xp5_ASAP7_75t_L g11828 ( 
.A1(n_11794),
.A2(n_1321),
.B1(n_1319),
.B2(n_1320),
.Y(n_11828)
);

OR2x2_ASAP7_75t_L g11829 ( 
.A(n_11567),
.B(n_1320),
.Y(n_11829)
);

INVx2_ASAP7_75t_L g11830 ( 
.A(n_11669),
.Y(n_11830)
);

AOI21xp5_ASAP7_75t_SL g11831 ( 
.A1(n_11780),
.A2(n_1321),
.B(n_1322),
.Y(n_11831)
);

AND2x2_ASAP7_75t_L g11832 ( 
.A(n_11480),
.B(n_1321),
.Y(n_11832)
);

OA21x2_ASAP7_75t_L g11833 ( 
.A1(n_11800),
.A2(n_11807),
.B(n_11802),
.Y(n_11833)
);

A2O1A1Ixp33_ASAP7_75t_L g11834 ( 
.A1(n_11476),
.A2(n_1324),
.B(n_1322),
.C(n_1323),
.Y(n_11834)
);

NAND2xp5_ASAP7_75t_L g11835 ( 
.A(n_11647),
.B(n_1322),
.Y(n_11835)
);

INVx2_ASAP7_75t_L g11836 ( 
.A(n_11528),
.Y(n_11836)
);

NAND2xp5_ASAP7_75t_L g11837 ( 
.A(n_11651),
.B(n_1323),
.Y(n_11837)
);

AND2x2_ASAP7_75t_L g11838 ( 
.A(n_11486),
.B(n_1323),
.Y(n_11838)
);

INVx2_ASAP7_75t_L g11839 ( 
.A(n_11472),
.Y(n_11839)
);

AOI21x1_ASAP7_75t_SL g11840 ( 
.A1(n_11733),
.A2(n_1324),
.B(n_1325),
.Y(n_11840)
);

INVx2_ASAP7_75t_L g11841 ( 
.A(n_11577),
.Y(n_11841)
);

INVx2_ASAP7_75t_SL g11842 ( 
.A(n_11505),
.Y(n_11842)
);

OAI22xp5_ASAP7_75t_SL g11843 ( 
.A1(n_11625),
.A2(n_1326),
.B1(n_1324),
.B2(n_1325),
.Y(n_11843)
);

INVx2_ASAP7_75t_SL g11844 ( 
.A(n_11506),
.Y(n_11844)
);

AND2x2_ASAP7_75t_L g11845 ( 
.A(n_11453),
.B(n_1325),
.Y(n_11845)
);

AND2x2_ASAP7_75t_L g11846 ( 
.A(n_11479),
.B(n_1326),
.Y(n_11846)
);

AND2x4_ASAP7_75t_L g11847 ( 
.A(n_11775),
.B(n_1327),
.Y(n_11847)
);

INVx1_ASAP7_75t_L g11848 ( 
.A(n_11657),
.Y(n_11848)
);

AND2x2_ASAP7_75t_L g11849 ( 
.A(n_11808),
.B(n_1327),
.Y(n_11849)
);

INVx1_ASAP7_75t_SL g11850 ( 
.A(n_11739),
.Y(n_11850)
);

AOI21x1_ASAP7_75t_SL g11851 ( 
.A1(n_11502),
.A2(n_1328),
.B(n_1329),
.Y(n_11851)
);

INVx1_ASAP7_75t_L g11852 ( 
.A(n_11660),
.Y(n_11852)
);

INVx1_ASAP7_75t_L g11853 ( 
.A(n_11490),
.Y(n_11853)
);

AND2x2_ASAP7_75t_L g11854 ( 
.A(n_11645),
.B(n_1328),
.Y(n_11854)
);

AND2x4_ASAP7_75t_L g11855 ( 
.A(n_11787),
.B(n_1328),
.Y(n_11855)
);

INVx1_ASAP7_75t_L g11856 ( 
.A(n_11501),
.Y(n_11856)
);

INVx1_ASAP7_75t_L g11857 ( 
.A(n_11508),
.Y(n_11857)
);

AND2x4_ASAP7_75t_L g11858 ( 
.A(n_11591),
.B(n_1329),
.Y(n_11858)
);

INVx1_ASAP7_75t_L g11859 ( 
.A(n_11510),
.Y(n_11859)
);

OA21x2_ASAP7_75t_L g11860 ( 
.A1(n_11818),
.A2(n_1330),
.B(n_1331),
.Y(n_11860)
);

BUFx3_ASAP7_75t_L g11861 ( 
.A(n_11784),
.Y(n_11861)
);

NAND2xp5_ASAP7_75t_L g11862 ( 
.A(n_11652),
.B(n_1330),
.Y(n_11862)
);

AO21x1_ASAP7_75t_L g11863 ( 
.A1(n_11461),
.A2(n_1330),
.B(n_1331),
.Y(n_11863)
);

HB1xp67_ASAP7_75t_L g11864 ( 
.A(n_11759),
.Y(n_11864)
);

AOI21x1_ASAP7_75t_SL g11865 ( 
.A1(n_11537),
.A2(n_1332),
.B(n_1333),
.Y(n_11865)
);

AND2x2_ASAP7_75t_L g11866 ( 
.A(n_11499),
.B(n_1332),
.Y(n_11866)
);

OAI31xp33_ASAP7_75t_SL g11867 ( 
.A1(n_11575),
.A2(n_1334),
.A3(n_1332),
.B(n_1333),
.Y(n_11867)
);

NAND2xp5_ASAP7_75t_L g11868 ( 
.A(n_11656),
.B(n_1333),
.Y(n_11868)
);

INVx1_ASAP7_75t_SL g11869 ( 
.A(n_11464),
.Y(n_11869)
);

OR2x2_ASAP7_75t_L g11870 ( 
.A(n_11473),
.B(n_11520),
.Y(n_11870)
);

OA21x2_ASAP7_75t_L g11871 ( 
.A1(n_11524),
.A2(n_1334),
.B(n_1335),
.Y(n_11871)
);

OAI22xp5_ASAP7_75t_L g11872 ( 
.A1(n_11483),
.A2(n_1337),
.B1(n_1335),
.B2(n_1336),
.Y(n_11872)
);

NOR2xp67_ASAP7_75t_L g11873 ( 
.A(n_11646),
.B(n_1335),
.Y(n_11873)
);

BUFx2_ASAP7_75t_L g11874 ( 
.A(n_11643),
.Y(n_11874)
);

AND2x2_ASAP7_75t_L g11875 ( 
.A(n_11522),
.B(n_1336),
.Y(n_11875)
);

HB1xp67_ASAP7_75t_L g11876 ( 
.A(n_11454),
.Y(n_11876)
);

BUFx3_ASAP7_75t_L g11877 ( 
.A(n_11493),
.Y(n_11877)
);

OR2x2_ASAP7_75t_L g11878 ( 
.A(n_11516),
.B(n_1337),
.Y(n_11878)
);

AND2x4_ASAP7_75t_L g11879 ( 
.A(n_11601),
.B(n_1337),
.Y(n_11879)
);

AOI21xp5_ASAP7_75t_SL g11880 ( 
.A1(n_11809),
.A2(n_1338),
.B(n_1339),
.Y(n_11880)
);

OR2x2_ASAP7_75t_L g11881 ( 
.A(n_11514),
.B(n_1338),
.Y(n_11881)
);

BUFx3_ASAP7_75t_L g11882 ( 
.A(n_11606),
.Y(n_11882)
);

NAND2xp5_ASAP7_75t_L g11883 ( 
.A(n_11542),
.B(n_1339),
.Y(n_11883)
);

OA21x2_ASAP7_75t_L g11884 ( 
.A1(n_11558),
.A2(n_1339),
.B(n_1340),
.Y(n_11884)
);

INVxp67_ASAP7_75t_L g11885 ( 
.A(n_11661),
.Y(n_11885)
);

OAI22xp5_ASAP7_75t_L g11886 ( 
.A1(n_11469),
.A2(n_11498),
.B1(n_11776),
.B2(n_11770),
.Y(n_11886)
);

OAI22xp5_ASAP7_75t_L g11887 ( 
.A1(n_11796),
.A2(n_1342),
.B1(n_1340),
.B2(n_1341),
.Y(n_11887)
);

AOI21xp5_ASAP7_75t_SL g11888 ( 
.A1(n_11708),
.A2(n_1340),
.B(n_1341),
.Y(n_11888)
);

NAND2xp5_ASAP7_75t_L g11889 ( 
.A(n_11554),
.B(n_1342),
.Y(n_11889)
);

INVx2_ASAP7_75t_L g11890 ( 
.A(n_11772),
.Y(n_11890)
);

AND2x4_ASAP7_75t_L g11891 ( 
.A(n_11452),
.B(n_1342),
.Y(n_11891)
);

OA21x2_ASAP7_75t_L g11892 ( 
.A1(n_11519),
.A2(n_1343),
.B(n_1344),
.Y(n_11892)
);

OR2x2_ASAP7_75t_L g11893 ( 
.A(n_11532),
.B(n_1343),
.Y(n_11893)
);

O2A1O1Ixp33_ASAP7_75t_L g11894 ( 
.A1(n_11509),
.A2(n_1345),
.B(n_1346),
.C(n_1344),
.Y(n_11894)
);

CKINVDCx5p33_ASAP7_75t_R g11895 ( 
.A(n_11570),
.Y(n_11895)
);

INVx1_ASAP7_75t_L g11896 ( 
.A(n_11518),
.Y(n_11896)
);

AOI22xp5_ASAP7_75t_L g11897 ( 
.A1(n_11460),
.A2(n_1345),
.B1(n_1343),
.B2(n_1344),
.Y(n_11897)
);

AND2x2_ASAP7_75t_L g11898 ( 
.A(n_11627),
.B(n_11675),
.Y(n_11898)
);

AND2x4_ASAP7_75t_L g11899 ( 
.A(n_11527),
.B(n_1346),
.Y(n_11899)
);

AOI21xp5_ASAP7_75t_SL g11900 ( 
.A1(n_11788),
.A2(n_1346),
.B(n_1347),
.Y(n_11900)
);

CKINVDCx5p33_ASAP7_75t_R g11901 ( 
.A(n_11517),
.Y(n_11901)
);

OR2x2_ASAP7_75t_L g11902 ( 
.A(n_11778),
.B(n_11477),
.Y(n_11902)
);

NOR2xp67_ASAP7_75t_L g11903 ( 
.A(n_11646),
.B(n_1347),
.Y(n_11903)
);

O2A1O1Ixp33_ASAP7_75t_L g11904 ( 
.A1(n_11676),
.A2(n_1349),
.B(n_1350),
.C(n_1348),
.Y(n_11904)
);

OA21x2_ASAP7_75t_L g11905 ( 
.A1(n_11727),
.A2(n_1347),
.B(n_1348),
.Y(n_11905)
);

CKINVDCx5p33_ASAP7_75t_R g11906 ( 
.A(n_11538),
.Y(n_11906)
);

AND2x2_ASAP7_75t_L g11907 ( 
.A(n_11471),
.B(n_1348),
.Y(n_11907)
);

NAND2xp5_ASAP7_75t_L g11908 ( 
.A(n_11799),
.B(n_1349),
.Y(n_11908)
);

NAND2xp5_ASAP7_75t_L g11909 ( 
.A(n_11814),
.B(n_1349),
.Y(n_11909)
);

AOI21xp5_ASAP7_75t_L g11910 ( 
.A1(n_11679),
.A2(n_1350),
.B(n_1351),
.Y(n_11910)
);

AOI21xp5_ASAP7_75t_L g11911 ( 
.A1(n_11475),
.A2(n_11639),
.B(n_11771),
.Y(n_11911)
);

AOI21x1_ASAP7_75t_SL g11912 ( 
.A1(n_11569),
.A2(n_1350),
.B(n_1351),
.Y(n_11912)
);

O2A1O1Ixp33_ASAP7_75t_L g11913 ( 
.A1(n_11682),
.A2(n_1354),
.B(n_1355),
.C(n_1352),
.Y(n_11913)
);

OAI22xp5_ASAP7_75t_L g11914 ( 
.A1(n_11458),
.A2(n_1354),
.B1(n_1351),
.B2(n_1352),
.Y(n_11914)
);

INVx2_ASAP7_75t_L g11915 ( 
.A(n_11772),
.Y(n_11915)
);

AOI21xp5_ASAP7_75t_SL g11916 ( 
.A1(n_11789),
.A2(n_1352),
.B(n_1354),
.Y(n_11916)
);

OAI22xp5_ASAP7_75t_SL g11917 ( 
.A1(n_11630),
.A2(n_1357),
.B1(n_1355),
.B2(n_1356),
.Y(n_11917)
);

BUFx3_ASAP7_75t_L g11918 ( 
.A(n_11608),
.Y(n_11918)
);

CKINVDCx5p33_ASAP7_75t_R g11919 ( 
.A(n_11555),
.Y(n_11919)
);

O2A1O1Ixp33_ASAP7_75t_L g11920 ( 
.A1(n_11560),
.A2(n_1359),
.B(n_1360),
.C(n_1358),
.Y(n_11920)
);

OAI22xp5_ASAP7_75t_L g11921 ( 
.A1(n_11485),
.A2(n_1359),
.B1(n_1356),
.B2(n_1358),
.Y(n_11921)
);

OAI22xp5_ASAP7_75t_L g11922 ( 
.A1(n_11744),
.A2(n_1359),
.B1(n_1356),
.B2(n_1358),
.Y(n_11922)
);

AND2x2_ASAP7_75t_L g11923 ( 
.A(n_11478),
.B(n_1360),
.Y(n_11923)
);

OA21x2_ASAP7_75t_L g11924 ( 
.A1(n_11466),
.A2(n_1360),
.B(n_1361),
.Y(n_11924)
);

NOR2xp33_ASAP7_75t_SL g11925 ( 
.A(n_11534),
.B(n_1361),
.Y(n_11925)
);

AOI21xp5_ASAP7_75t_L g11926 ( 
.A1(n_11773),
.A2(n_1361),
.B(n_1362),
.Y(n_11926)
);

NAND2xp5_ASAP7_75t_L g11927 ( 
.A(n_11563),
.B(n_1363),
.Y(n_11927)
);

OA22x2_ASAP7_75t_L g11928 ( 
.A1(n_11741),
.A2(n_1365),
.B1(n_1363),
.B2(n_1364),
.Y(n_11928)
);

A2O1A1Ixp33_ASAP7_75t_L g11929 ( 
.A1(n_11565),
.A2(n_1366),
.B(n_1364),
.C(n_1365),
.Y(n_11929)
);

AOI21x1_ASAP7_75t_SL g11930 ( 
.A1(n_11603),
.A2(n_1364),
.B(n_1366),
.Y(n_11930)
);

HB1xp67_ASAP7_75t_L g11931 ( 
.A(n_11539),
.Y(n_11931)
);

AOI21xp5_ASAP7_75t_L g11932 ( 
.A1(n_11793),
.A2(n_1366),
.B(n_1367),
.Y(n_11932)
);

INVx1_ASAP7_75t_L g11933 ( 
.A(n_11525),
.Y(n_11933)
);

INVx1_ASAP7_75t_L g11934 ( 
.A(n_11564),
.Y(n_11934)
);

INVx1_ASAP7_75t_L g11935 ( 
.A(n_11594),
.Y(n_11935)
);

A2O1A1Ixp33_ASAP7_75t_L g11936 ( 
.A1(n_11640),
.A2(n_11494),
.B(n_11449),
.C(n_11474),
.Y(n_11936)
);

CKINVDCx11_ASAP7_75t_R g11937 ( 
.A(n_11804),
.Y(n_11937)
);

NAND2xp5_ASAP7_75t_L g11938 ( 
.A(n_11644),
.B(n_1367),
.Y(n_11938)
);

OAI22xp5_ASAP7_75t_L g11939 ( 
.A1(n_11511),
.A2(n_1370),
.B1(n_1368),
.B2(n_1369),
.Y(n_11939)
);

OA21x2_ASAP7_75t_L g11940 ( 
.A1(n_11810),
.A2(n_1368),
.B(n_1369),
.Y(n_11940)
);

OAI22xp5_ASAP7_75t_L g11941 ( 
.A1(n_11709),
.A2(n_11481),
.B1(n_11748),
.B2(n_11482),
.Y(n_11941)
);

AOI21xp5_ASAP7_75t_L g11942 ( 
.A1(n_11817),
.A2(n_1368),
.B(n_1369),
.Y(n_11942)
);

HB1xp67_ASAP7_75t_L g11943 ( 
.A(n_11700),
.Y(n_11943)
);

AOI21x1_ASAP7_75t_SL g11944 ( 
.A1(n_11615),
.A2(n_1370),
.B(n_1371),
.Y(n_11944)
);

OA21x2_ASAP7_75t_L g11945 ( 
.A1(n_11680),
.A2(n_1370),
.B(n_1371),
.Y(n_11945)
);

BUFx6f_ASAP7_75t_L g11946 ( 
.A(n_11549),
.Y(n_11946)
);

AND2x4_ASAP7_75t_L g11947 ( 
.A(n_11447),
.B(n_1371),
.Y(n_11947)
);

NAND2xp5_ASAP7_75t_L g11948 ( 
.A(n_11571),
.B(n_1372),
.Y(n_11948)
);

BUFx3_ASAP7_75t_L g11949 ( 
.A(n_11636),
.Y(n_11949)
);

HB1xp67_ASAP7_75t_L g11950 ( 
.A(n_11758),
.Y(n_11950)
);

AND2x2_ASAP7_75t_L g11951 ( 
.A(n_11694),
.B(n_1372),
.Y(n_11951)
);

AOI21xp5_ASAP7_75t_SL g11952 ( 
.A1(n_11805),
.A2(n_11710),
.B(n_11552),
.Y(n_11952)
);

AOI21xp5_ASAP7_75t_SL g11953 ( 
.A1(n_11535),
.A2(n_11578),
.B(n_11786),
.Y(n_11953)
);

NAND2xp5_ASAP7_75t_L g11954 ( 
.A(n_11732),
.B(n_1373),
.Y(n_11954)
);

NAND2xp5_ASAP7_75t_L g11955 ( 
.A(n_11735),
.B(n_1373),
.Y(n_11955)
);

NAND2xp5_ASAP7_75t_L g11956 ( 
.A(n_11750),
.B(n_1373),
.Y(n_11956)
);

OA21x2_ASAP7_75t_L g11957 ( 
.A1(n_11497),
.A2(n_1374),
.B(n_1375),
.Y(n_11957)
);

OR2x2_ASAP7_75t_L g11958 ( 
.A(n_11782),
.B(n_1374),
.Y(n_11958)
);

A2O1A1Ixp33_ASAP7_75t_SL g11959 ( 
.A1(n_11769),
.A2(n_1377),
.B(n_1375),
.C(n_1376),
.Y(n_11959)
);

OR2x2_ASAP7_75t_L g11960 ( 
.A(n_11783),
.B(n_1375),
.Y(n_11960)
);

A2O1A1Ixp33_ASAP7_75t_L g11961 ( 
.A1(n_11451),
.A2(n_1378),
.B(n_1376),
.C(n_1377),
.Y(n_11961)
);

OR2x2_ASAP7_75t_L g11962 ( 
.A(n_11812),
.B(n_1377),
.Y(n_11962)
);

O2A1O1Ixp33_ASAP7_75t_L g11963 ( 
.A1(n_11642),
.A2(n_1380),
.B(n_1381),
.C(n_1379),
.Y(n_11963)
);

OAI22xp5_ASAP7_75t_L g11964 ( 
.A1(n_11734),
.A2(n_1380),
.B1(n_1378),
.B2(n_1379),
.Y(n_11964)
);

AOI21x1_ASAP7_75t_SL g11965 ( 
.A1(n_11546),
.A2(n_1381),
.B(n_1382),
.Y(n_11965)
);

AND2x2_ASAP7_75t_L g11966 ( 
.A(n_11813),
.B(n_1381),
.Y(n_11966)
);

O2A1O1Ixp33_ASAP7_75t_L g11967 ( 
.A1(n_11600),
.A2(n_1384),
.B(n_1385),
.C(n_1383),
.Y(n_11967)
);

OAI211xp5_ASAP7_75t_L g11968 ( 
.A1(n_11703),
.A2(n_11754),
.B(n_11576),
.C(n_11597),
.Y(n_11968)
);

NOR2x1_ASAP7_75t_SL g11969 ( 
.A(n_11586),
.B(n_1382),
.Y(n_11969)
);

NAND2xp5_ASAP7_75t_L g11970 ( 
.A(n_11753),
.B(n_1384),
.Y(n_11970)
);

OAI22xp5_ASAP7_75t_L g11971 ( 
.A1(n_11692),
.A2(n_11470),
.B1(n_11681),
.B2(n_11489),
.Y(n_11971)
);

AND2x2_ASAP7_75t_L g11972 ( 
.A(n_11813),
.B(n_1384),
.Y(n_11972)
);

OA21x2_ASAP7_75t_L g11973 ( 
.A1(n_11637),
.A2(n_1385),
.B(n_1386),
.Y(n_11973)
);

AOI21x1_ASAP7_75t_SL g11974 ( 
.A1(n_11626),
.A2(n_1385),
.B(n_1386),
.Y(n_11974)
);

O2A1O1Ixp33_ASAP7_75t_L g11975 ( 
.A1(n_11716),
.A2(n_1389),
.B(n_1390),
.C(n_1388),
.Y(n_11975)
);

HB1xp67_ASAP7_75t_L g11976 ( 
.A(n_11761),
.Y(n_11976)
);

INVx2_ASAP7_75t_L g11977 ( 
.A(n_11777),
.Y(n_11977)
);

AOI21xp5_ASAP7_75t_L g11978 ( 
.A1(n_11544),
.A2(n_1387),
.B(n_1388),
.Y(n_11978)
);

NAND2xp5_ASAP7_75t_L g11979 ( 
.A(n_11760),
.B(n_1387),
.Y(n_11979)
);

OR2x2_ASAP7_75t_L g11980 ( 
.A(n_11595),
.B(n_1388),
.Y(n_11980)
);

BUFx6f_ASAP7_75t_L g11981 ( 
.A(n_11610),
.Y(n_11981)
);

O2A1O1Ixp33_ASAP7_75t_L g11982 ( 
.A1(n_11596),
.A2(n_1392),
.B(n_1393),
.C(n_1391),
.Y(n_11982)
);

AOI21xp5_ASAP7_75t_L g11983 ( 
.A1(n_11541),
.A2(n_1389),
.B(n_1391),
.Y(n_11983)
);

AND2x4_ASAP7_75t_L g11984 ( 
.A(n_11631),
.B(n_1389),
.Y(n_11984)
);

HB1xp67_ASAP7_75t_L g11985 ( 
.A(n_11730),
.Y(n_11985)
);

AOI21x1_ASAP7_75t_SL g11986 ( 
.A1(n_11611),
.A2(n_1391),
.B(n_1392),
.Y(n_11986)
);

O2A1O1Ixp5_ASAP7_75t_L g11987 ( 
.A1(n_11635),
.A2(n_1395),
.B(n_1393),
.C(n_1394),
.Y(n_11987)
);

NOR2xp67_ASAP7_75t_L g11988 ( 
.A(n_11593),
.B(n_1393),
.Y(n_11988)
);

AND2x2_ASAP7_75t_L g11989 ( 
.A(n_11658),
.B(n_1395),
.Y(n_11989)
);

OA21x2_ASAP7_75t_L g11990 ( 
.A1(n_11702),
.A2(n_1395),
.B(n_1396),
.Y(n_11990)
);

AOI21xp5_ASAP7_75t_SL g11991 ( 
.A1(n_11459),
.A2(n_1397),
.B(n_1398),
.Y(n_11991)
);

AOI31xp33_ASAP7_75t_L g11992 ( 
.A1(n_11602),
.A2(n_1406),
.A3(n_1414),
.B(n_1397),
.Y(n_11992)
);

HB1xp67_ASAP7_75t_L g11993 ( 
.A(n_11704),
.Y(n_11993)
);

NAND2xp5_ASAP7_75t_L g11994 ( 
.A(n_11711),
.B(n_1397),
.Y(n_11994)
);

OAI22xp5_ASAP7_75t_L g11995 ( 
.A1(n_11671),
.A2(n_1401),
.B1(n_1398),
.B2(n_1400),
.Y(n_11995)
);

CKINVDCx6p67_ASAP7_75t_R g11996 ( 
.A(n_11531),
.Y(n_11996)
);

AND2x2_ASAP7_75t_L g11997 ( 
.A(n_11720),
.B(n_1398),
.Y(n_11997)
);

AND2x2_ASAP7_75t_L g11998 ( 
.A(n_11740),
.B(n_1400),
.Y(n_11998)
);

O2A1O1Ixp33_ASAP7_75t_L g11999 ( 
.A1(n_11550),
.A2(n_1402),
.B(n_1403),
.C(n_1401),
.Y(n_11999)
);

O2A1O1Ixp33_ASAP7_75t_L g12000 ( 
.A1(n_11496),
.A2(n_11604),
.B(n_11687),
.C(n_11668),
.Y(n_12000)
);

NOR2xp67_ASAP7_75t_L g12001 ( 
.A(n_11583),
.B(n_1400),
.Y(n_12001)
);

AND2x4_ASAP7_75t_SL g12002 ( 
.A(n_11573),
.B(n_1401),
.Y(n_12002)
);

AOI21xp5_ASAP7_75t_SL g12003 ( 
.A1(n_11713),
.A2(n_1402),
.B(n_1403),
.Y(n_12003)
);

OAI22xp5_ASAP7_75t_L g12004 ( 
.A1(n_11629),
.A2(n_11663),
.B1(n_11743),
.B2(n_11559),
.Y(n_12004)
);

OAI22xp5_ASAP7_75t_L g12005 ( 
.A1(n_11723),
.A2(n_1406),
.B1(n_1404),
.B2(n_1405),
.Y(n_12005)
);

AND2x2_ASAP7_75t_L g12006 ( 
.A(n_11589),
.B(n_1404),
.Y(n_12006)
);

AND2x4_ASAP7_75t_L g12007 ( 
.A(n_11729),
.B(n_11641),
.Y(n_12007)
);

O2A1O1Ixp5_ASAP7_75t_L g12008 ( 
.A1(n_11659),
.A2(n_1407),
.B(n_1405),
.C(n_1406),
.Y(n_12008)
);

AND2x2_ASAP7_75t_L g12009 ( 
.A(n_11690),
.B(n_1405),
.Y(n_12009)
);

INVx1_ASAP7_75t_L g12010 ( 
.A(n_11777),
.Y(n_12010)
);

NAND2x1_ASAP7_75t_L g12011 ( 
.A(n_11487),
.B(n_1407),
.Y(n_12011)
);

OA21x2_ASAP7_75t_L g12012 ( 
.A1(n_11580),
.A2(n_1408),
.B(n_1409),
.Y(n_12012)
);

INVx2_ASAP7_75t_L g12013 ( 
.A(n_11590),
.Y(n_12013)
);

AND2x2_ASAP7_75t_L g12014 ( 
.A(n_11543),
.B(n_1408),
.Y(n_12014)
);

AND2x2_ASAP7_75t_L g12015 ( 
.A(n_11745),
.B(n_1409),
.Y(n_12015)
);

NOR2xp67_ASAP7_75t_L g12016 ( 
.A(n_11495),
.B(n_1409),
.Y(n_12016)
);

NAND2xp5_ASAP7_75t_L g12017 ( 
.A(n_11512),
.B(n_1410),
.Y(n_12017)
);

NAND2xp5_ASAP7_75t_L g12018 ( 
.A(n_11515),
.B(n_1410),
.Y(n_12018)
);

INVx2_ASAP7_75t_L g12019 ( 
.A(n_11609),
.Y(n_12019)
);

A2O1A1Ixp33_ASAP7_75t_L g12020 ( 
.A1(n_11455),
.A2(n_1412),
.B(n_1410),
.C(n_1411),
.Y(n_12020)
);

INVx4_ASAP7_75t_L g12021 ( 
.A(n_11649),
.Y(n_12021)
);

INVx1_ASAP7_75t_L g12022 ( 
.A(n_11791),
.Y(n_12022)
);

AOI21xp5_ASAP7_75t_L g12023 ( 
.A1(n_11556),
.A2(n_1411),
.B(n_1412),
.Y(n_12023)
);

AND2x2_ASAP7_75t_L g12024 ( 
.A(n_11649),
.B(n_1411),
.Y(n_12024)
);

O2A1O1Ixp33_ASAP7_75t_L g12025 ( 
.A1(n_11488),
.A2(n_1415),
.B(n_1416),
.C(n_1414),
.Y(n_12025)
);

OAI22xp5_ASAP7_75t_L g12026 ( 
.A1(n_11738),
.A2(n_1416),
.B1(n_1413),
.B2(n_1415),
.Y(n_12026)
);

AOI21xp5_ASAP7_75t_L g12027 ( 
.A1(n_11579),
.A2(n_1417),
.B(n_1418),
.Y(n_12027)
);

OAI22xp5_ASAP7_75t_L g12028 ( 
.A1(n_11530),
.A2(n_1419),
.B1(n_1417),
.B2(n_1418),
.Y(n_12028)
);

NAND2xp5_ASAP7_75t_L g12029 ( 
.A(n_11581),
.B(n_1418),
.Y(n_12029)
);

NOR2xp67_ASAP7_75t_L g12030 ( 
.A(n_11500),
.B(n_1419),
.Y(n_12030)
);

AOI221xp5_ASAP7_75t_L g12031 ( 
.A1(n_11691),
.A2(n_1421),
.B1(n_1419),
.B2(n_1420),
.C(n_1422),
.Y(n_12031)
);

BUFx3_ASAP7_75t_L g12032 ( 
.A(n_11674),
.Y(n_12032)
);

OR2x2_ASAP7_75t_L g12033 ( 
.A(n_11562),
.B(n_1421),
.Y(n_12033)
);

AND2x2_ASAP7_75t_L g12034 ( 
.A(n_11662),
.B(n_1421),
.Y(n_12034)
);

CKINVDCx11_ASAP7_75t_R g12035 ( 
.A(n_11677),
.Y(n_12035)
);

OAI22xp5_ASAP7_75t_L g12036 ( 
.A1(n_11816),
.A2(n_11670),
.B1(n_11798),
.B2(n_11689),
.Y(n_12036)
);

AND2x2_ASAP7_75t_L g12037 ( 
.A(n_11448),
.B(n_1422),
.Y(n_12037)
);

OAI22xp5_ASAP7_75t_L g12038 ( 
.A1(n_11678),
.A2(n_1424),
.B1(n_1422),
.B2(n_1423),
.Y(n_12038)
);

HB1xp67_ASAP7_75t_L g12039 ( 
.A(n_11523),
.Y(n_12039)
);

INVx1_ASAP7_75t_L g12040 ( 
.A(n_11696),
.Y(n_12040)
);

INVx1_ASAP7_75t_L g12041 ( 
.A(n_11664),
.Y(n_12041)
);

AND2x2_ASAP7_75t_L g12042 ( 
.A(n_11633),
.B(n_1423),
.Y(n_12042)
);

OA21x2_ASAP7_75t_L g12043 ( 
.A1(n_11513),
.A2(n_1423),
.B(n_1424),
.Y(n_12043)
);

AND2x2_ASAP7_75t_L g12044 ( 
.A(n_11633),
.B(n_1424),
.Y(n_12044)
);

OAI22xp5_ASAP7_75t_L g12045 ( 
.A1(n_11684),
.A2(n_1427),
.B1(n_1425),
.B2(n_1426),
.Y(n_12045)
);

O2A1O1Ixp5_ASAP7_75t_L g12046 ( 
.A1(n_11620),
.A2(n_1427),
.B(n_1425),
.C(n_1426),
.Y(n_12046)
);

INVx3_ASAP7_75t_L g12047 ( 
.A(n_11706),
.Y(n_12047)
);

OA21x2_ASAP7_75t_L g12048 ( 
.A1(n_11705),
.A2(n_1425),
.B(n_1427),
.Y(n_12048)
);

AND2x2_ASAP7_75t_L g12049 ( 
.A(n_11628),
.B(n_1428),
.Y(n_12049)
);

BUFx2_ASAP7_75t_L g12050 ( 
.A(n_11634),
.Y(n_12050)
);

AOI21xp5_ASAP7_75t_SL g12051 ( 
.A1(n_11572),
.A2(n_1428),
.B(n_1429),
.Y(n_12051)
);

INVxp67_ASAP7_75t_L g12052 ( 
.A(n_11599),
.Y(n_12052)
);

INVx1_ASAP7_75t_L g12053 ( 
.A(n_11664),
.Y(n_12053)
);

AND2x4_ASAP7_75t_L g12054 ( 
.A(n_11706),
.B(n_1428),
.Y(n_12054)
);

OA21x2_ASAP7_75t_L g12055 ( 
.A1(n_11521),
.A2(n_1429),
.B(n_1430),
.Y(n_12055)
);

OR2x2_ASAP7_75t_L g12056 ( 
.A(n_11491),
.B(n_11655),
.Y(n_12056)
);

INVx2_ASAP7_75t_L g12057 ( 
.A(n_11547),
.Y(n_12057)
);

INVx2_ASAP7_75t_L g12058 ( 
.A(n_11548),
.Y(n_12058)
);

OR2x2_ASAP7_75t_L g12059 ( 
.A(n_11491),
.B(n_1429),
.Y(n_12059)
);

OAI22xp5_ASAP7_75t_L g12060 ( 
.A1(n_11746),
.A2(n_1432),
.B1(n_1430),
.B2(n_1431),
.Y(n_12060)
);

INVx1_ASAP7_75t_L g12061 ( 
.A(n_11529),
.Y(n_12061)
);

AND2x4_ASAP7_75t_L g12062 ( 
.A(n_11585),
.B(n_11619),
.Y(n_12062)
);

OAI22xp5_ASAP7_75t_L g12063 ( 
.A1(n_11621),
.A2(n_11724),
.B1(n_11557),
.B2(n_11781),
.Y(n_12063)
);

CKINVDCx5p33_ASAP7_75t_R g12064 ( 
.A(n_11674),
.Y(n_12064)
);

INVx2_ASAP7_75t_L g12065 ( 
.A(n_11721),
.Y(n_12065)
);

AND2x2_ASAP7_75t_L g12066 ( 
.A(n_11446),
.B(n_11686),
.Y(n_12066)
);

AOI21x1_ASAP7_75t_SL g12067 ( 
.A1(n_11714),
.A2(n_1430),
.B(n_1431),
.Y(n_12067)
);

INVx1_ASAP7_75t_L g12068 ( 
.A(n_11582),
.Y(n_12068)
);

OAI22xp5_ASAP7_75t_L g12069 ( 
.A1(n_11795),
.A2(n_1433),
.B1(n_1431),
.B2(n_1432),
.Y(n_12069)
);

NAND2xp5_ASAP7_75t_L g12070 ( 
.A(n_11650),
.B(n_1433),
.Y(n_12070)
);

AND2x2_ASAP7_75t_L g12071 ( 
.A(n_11612),
.B(n_1434),
.Y(n_12071)
);

INVx1_ASAP7_75t_L g12072 ( 
.A(n_11683),
.Y(n_12072)
);

HB1xp67_ASAP7_75t_L g12073 ( 
.A(n_11507),
.Y(n_12073)
);

NAND2xp5_ASAP7_75t_L g12074 ( 
.A(n_11688),
.B(n_11467),
.Y(n_12074)
);

AOI21x1_ASAP7_75t_SL g12075 ( 
.A1(n_11763),
.A2(n_1434),
.B(n_1435),
.Y(n_12075)
);

A2O1A1Ixp33_ASAP7_75t_L g12076 ( 
.A1(n_11456),
.A2(n_1436),
.B(n_1434),
.C(n_1435),
.Y(n_12076)
);

AND2x2_ASAP7_75t_L g12077 ( 
.A(n_11450),
.B(n_1435),
.Y(n_12077)
);

NAND2xp5_ASAP7_75t_L g12078 ( 
.A(n_11701),
.B(n_1436),
.Y(n_12078)
);

NAND2xp5_ASAP7_75t_L g12079 ( 
.A(n_11592),
.B(n_1436),
.Y(n_12079)
);

AND2x2_ASAP7_75t_L g12080 ( 
.A(n_11685),
.B(n_1437),
.Y(n_12080)
);

INVx1_ASAP7_75t_L g12081 ( 
.A(n_11737),
.Y(n_12081)
);

INVx2_ASAP7_75t_L g12082 ( 
.A(n_11533),
.Y(n_12082)
);

AOI21xp5_ASAP7_75t_SL g12083 ( 
.A1(n_11715),
.A2(n_1437),
.B(n_1438),
.Y(n_12083)
);

HB1xp67_ASAP7_75t_L g12084 ( 
.A(n_11492),
.Y(n_12084)
);

CKINVDCx5p33_ASAP7_75t_R g12085 ( 
.A(n_11685),
.Y(n_12085)
);

NAND2xp5_ASAP7_75t_SL g12086 ( 
.A(n_11774),
.B(n_11792),
.Y(n_12086)
);

OAI22xp5_ASAP7_75t_L g12087 ( 
.A1(n_11801),
.A2(n_1440),
.B1(n_1438),
.B2(n_1439),
.Y(n_12087)
);

AND2x2_ASAP7_75t_L g12088 ( 
.A(n_11592),
.B(n_1438),
.Y(n_12088)
);

OAI22xp5_ASAP7_75t_L g12089 ( 
.A1(n_11697),
.A2(n_11736),
.B1(n_11752),
.B2(n_11764),
.Y(n_12089)
);

AND2x2_ASAP7_75t_L g12090 ( 
.A(n_11605),
.B(n_1439),
.Y(n_12090)
);

A2O1A1Ixp33_ASAP7_75t_L g12091 ( 
.A1(n_11468),
.A2(n_11463),
.B(n_11462),
.C(n_11484),
.Y(n_12091)
);

INVx1_ASAP7_75t_L g12092 ( 
.A(n_11749),
.Y(n_12092)
);

AND2x2_ASAP7_75t_L g12093 ( 
.A(n_11693),
.B(n_1439),
.Y(n_12093)
);

INVx3_ASAP7_75t_SL g12094 ( 
.A(n_11672),
.Y(n_12094)
);

CKINVDCx20_ASAP7_75t_R g12095 ( 
.A(n_11726),
.Y(n_12095)
);

AOI21xp5_ASAP7_75t_L g12096 ( 
.A1(n_11504),
.A2(n_11503),
.B(n_11698),
.Y(n_12096)
);

INVx2_ASAP7_75t_L g12097 ( 
.A(n_11553),
.Y(n_12097)
);

AND2x4_ASAP7_75t_L g12098 ( 
.A(n_11747),
.B(n_1440),
.Y(n_12098)
);

NAND2xp5_ASAP7_75t_L g12099 ( 
.A(n_11653),
.B(n_1441),
.Y(n_12099)
);

BUFx6f_ASAP7_75t_L g12100 ( 
.A(n_11667),
.Y(n_12100)
);

HB1xp67_ASAP7_75t_L g12101 ( 
.A(n_11695),
.Y(n_12101)
);

OAI22xp5_ASAP7_75t_L g12102 ( 
.A1(n_11613),
.A2(n_1443),
.B1(n_1441),
.B2(n_1442),
.Y(n_12102)
);

NAND2xp5_ASAP7_75t_L g12103 ( 
.A(n_11653),
.B(n_1442),
.Y(n_12103)
);

AND2x4_ASAP7_75t_L g12104 ( 
.A(n_11751),
.B(n_1443),
.Y(n_12104)
);

AOI21xp5_ASAP7_75t_L g12105 ( 
.A1(n_11767),
.A2(n_1443),
.B(n_1444),
.Y(n_12105)
);

AOI21x1_ASAP7_75t_SL g12106 ( 
.A1(n_11551),
.A2(n_1444),
.B(n_1445),
.Y(n_12106)
);

AND2x4_ASAP7_75t_L g12107 ( 
.A(n_11526),
.B(n_1444),
.Y(n_12107)
);

O2A1O1Ixp33_ASAP7_75t_L g12108 ( 
.A1(n_11762),
.A2(n_1447),
.B(n_1448),
.C(n_1446),
.Y(n_12108)
);

NAND2xp5_ASAP7_75t_L g12109 ( 
.A(n_11465),
.B(n_1445),
.Y(n_12109)
);

AOI21xp5_ASAP7_75t_SL g12110 ( 
.A1(n_11712),
.A2(n_11719),
.B(n_11598),
.Y(n_12110)
);

OR2x2_ASAP7_75t_L g12111 ( 
.A(n_11756),
.B(n_1446),
.Y(n_12111)
);

AOI21xp5_ASAP7_75t_L g12112 ( 
.A1(n_11587),
.A2(n_1446),
.B(n_1447),
.Y(n_12112)
);

AND2x2_ASAP7_75t_L g12113 ( 
.A(n_11779),
.B(n_1448),
.Y(n_12113)
);

O2A1O1Ixp33_ASAP7_75t_L g12114 ( 
.A1(n_11465),
.A2(n_1450),
.B(n_1451),
.C(n_1449),
.Y(n_12114)
);

OAI22xp5_ASAP7_75t_L g12115 ( 
.A1(n_11622),
.A2(n_1450),
.B1(n_1448),
.B2(n_1449),
.Y(n_12115)
);

AND2x4_ASAP7_75t_L g12116 ( 
.A(n_11654),
.B(n_1449),
.Y(n_12116)
);

CKINVDCx20_ASAP7_75t_R g12117 ( 
.A(n_11566),
.Y(n_12117)
);

AOI21x1_ASAP7_75t_SL g12118 ( 
.A1(n_11624),
.A2(n_1450),
.B(n_1451),
.Y(n_12118)
);

NAND2xp5_ASAP7_75t_L g12119 ( 
.A(n_11756),
.B(n_1451),
.Y(n_12119)
);

OAI22xp5_ASAP7_75t_L g12120 ( 
.A1(n_11699),
.A2(n_11707),
.B1(n_11718),
.B2(n_11717),
.Y(n_12120)
);

AND2x2_ASAP7_75t_L g12121 ( 
.A(n_11785),
.B(n_1452),
.Y(n_12121)
);

INVx2_ASAP7_75t_L g12122 ( 
.A(n_11568),
.Y(n_12122)
);

NAND2xp5_ASAP7_75t_L g12123 ( 
.A(n_11707),
.B(n_1452),
.Y(n_12123)
);

O2A1O1Ixp33_ASAP7_75t_L g12124 ( 
.A1(n_11722),
.A2(n_1455),
.B(n_1456),
.C(n_1454),
.Y(n_12124)
);

OA21x2_ASAP7_75t_L g12125 ( 
.A1(n_11815),
.A2(n_1453),
.B(n_1454),
.Y(n_12125)
);

AOI21xp5_ASAP7_75t_SL g12126 ( 
.A1(n_11790),
.A2(n_1453),
.B(n_1454),
.Y(n_12126)
);

OR2x2_ASAP7_75t_L g12127 ( 
.A(n_11540),
.B(n_11536),
.Y(n_12127)
);

AOI221xp5_ASAP7_75t_L g12128 ( 
.A1(n_11648),
.A2(n_1457),
.B1(n_1455),
.B2(n_1456),
.C(n_1458),
.Y(n_12128)
);

INVx1_ASAP7_75t_L g12129 ( 
.A(n_11561),
.Y(n_12129)
);

INVx1_ASAP7_75t_L g12130 ( 
.A(n_11618),
.Y(n_12130)
);

AOI21x1_ASAP7_75t_SL g12131 ( 
.A1(n_11806),
.A2(n_1456),
.B(n_1457),
.Y(n_12131)
);

NAND2xp5_ASAP7_75t_L g12132 ( 
.A(n_11623),
.B(n_1457),
.Y(n_12132)
);

BUFx2_ASAP7_75t_L g12133 ( 
.A(n_11584),
.Y(n_12133)
);

OAI22xp5_ASAP7_75t_L g12134 ( 
.A1(n_11666),
.A2(n_1460),
.B1(n_1458),
.B2(n_1459),
.Y(n_12134)
);

AOI21xp5_ASAP7_75t_SL g12135 ( 
.A1(n_11616),
.A2(n_1458),
.B(n_1459),
.Y(n_12135)
);

OA21x2_ASAP7_75t_L g12136 ( 
.A1(n_11638),
.A2(n_1459),
.B(n_1460),
.Y(n_12136)
);

AND2x2_ASAP7_75t_L g12137 ( 
.A(n_11588),
.B(n_1460),
.Y(n_12137)
);

NAND2xp5_ASAP7_75t_L g12138 ( 
.A(n_11665),
.B(n_1461),
.Y(n_12138)
);

BUFx3_ASAP7_75t_L g12139 ( 
.A(n_11768),
.Y(n_12139)
);

A2O1A1Ixp33_ASAP7_75t_SL g12140 ( 
.A1(n_11725),
.A2(n_1464),
.B(n_1462),
.C(n_1463),
.Y(n_12140)
);

NOR3xp33_ASAP7_75t_L g12141 ( 
.A(n_11673),
.B(n_1462),
.C(n_1463),
.Y(n_12141)
);

OAI22xp5_ASAP7_75t_L g12142 ( 
.A1(n_11728),
.A2(n_1464),
.B1(n_1462),
.B2(n_1463),
.Y(n_12142)
);

AND2x2_ASAP7_75t_L g12143 ( 
.A(n_11731),
.B(n_1465),
.Y(n_12143)
);

AOI21x1_ASAP7_75t_SL g12144 ( 
.A1(n_11765),
.A2(n_1465),
.B(n_1466),
.Y(n_12144)
);

INVx1_ASAP7_75t_L g12145 ( 
.A(n_11766),
.Y(n_12145)
);

AND2x4_ASAP7_75t_L g12146 ( 
.A(n_11757),
.B(n_1466),
.Y(n_12146)
);

INVx3_ASAP7_75t_L g12147 ( 
.A(n_11742),
.Y(n_12147)
);

A2O1A1Ixp33_ASAP7_75t_L g12148 ( 
.A1(n_11755),
.A2(n_1468),
.B(n_1466),
.C(n_1467),
.Y(n_12148)
);

A2O1A1Ixp33_ASAP7_75t_L g12149 ( 
.A1(n_11476),
.A2(n_1469),
.B(n_1467),
.C(n_1468),
.Y(n_12149)
);

NAND2xp5_ASAP7_75t_L g12150 ( 
.A(n_11614),
.B(n_1467),
.Y(n_12150)
);

INVx1_ASAP7_75t_L g12151 ( 
.A(n_11657),
.Y(n_12151)
);

INVx1_ASAP7_75t_SL g12152 ( 
.A(n_11632),
.Y(n_12152)
);

O2A1O1Ixp33_ASAP7_75t_L g12153 ( 
.A1(n_11509),
.A2(n_1470),
.B(n_1471),
.C(n_1469),
.Y(n_12153)
);

NAND2xp5_ASAP7_75t_L g12154 ( 
.A(n_11614),
.B(n_1468),
.Y(n_12154)
);

HB1xp67_ASAP7_75t_L g12155 ( 
.A(n_11607),
.Y(n_12155)
);

INVx2_ASAP7_75t_L g12156 ( 
.A(n_11669),
.Y(n_12156)
);

OAI211xp5_ASAP7_75t_L g12157 ( 
.A1(n_11509),
.A2(n_1473),
.B(n_1471),
.C(n_1472),
.Y(n_12157)
);

HB1xp67_ASAP7_75t_L g12158 ( 
.A(n_11607),
.Y(n_12158)
);

NAND2xp5_ASAP7_75t_L g12159 ( 
.A(n_11614),
.B(n_1473),
.Y(n_12159)
);

AND2x2_ASAP7_75t_L g12160 ( 
.A(n_11545),
.B(n_1473),
.Y(n_12160)
);

AOI21x1_ASAP7_75t_SL g12161 ( 
.A1(n_11457),
.A2(n_1474),
.B(n_1475),
.Y(n_12161)
);

OAI22xp5_ASAP7_75t_L g12162 ( 
.A1(n_11545),
.A2(n_1476),
.B1(n_1474),
.B2(n_1475),
.Y(n_12162)
);

INVx1_ASAP7_75t_L g12163 ( 
.A(n_11657),
.Y(n_12163)
);

INVx1_ASAP7_75t_L g12164 ( 
.A(n_11657),
.Y(n_12164)
);

OAI22xp5_ASAP7_75t_L g12165 ( 
.A1(n_11545),
.A2(n_1477),
.B1(n_1474),
.B2(n_1476),
.Y(n_12165)
);

O2A1O1Ixp33_ASAP7_75t_L g12166 ( 
.A1(n_11509),
.A2(n_1479),
.B(n_1480),
.C(n_1478),
.Y(n_12166)
);

INVx1_ASAP7_75t_L g12167 ( 
.A(n_11657),
.Y(n_12167)
);

OAI31xp33_ASAP7_75t_L g12168 ( 
.A1(n_11469),
.A2(n_1480),
.A3(n_1476),
.B(n_1479),
.Y(n_12168)
);

OAI22xp5_ASAP7_75t_L g12169 ( 
.A1(n_11545),
.A2(n_1482),
.B1(n_1480),
.B2(n_1481),
.Y(n_12169)
);

OA21x2_ASAP7_75t_L g12170 ( 
.A1(n_11545),
.A2(n_1482),
.B(n_1483),
.Y(n_12170)
);

INVx1_ASAP7_75t_L g12171 ( 
.A(n_11657),
.Y(n_12171)
);

AOI211xp5_ASAP7_75t_L g12172 ( 
.A1(n_11509),
.A2(n_1484),
.B(n_1482),
.C(n_1483),
.Y(n_12172)
);

OAI211xp5_ASAP7_75t_L g12173 ( 
.A1(n_11509),
.A2(n_1486),
.B(n_1484),
.C(n_1485),
.Y(n_12173)
);

OA21x2_ASAP7_75t_L g12174 ( 
.A1(n_11545),
.A2(n_1484),
.B(n_1485),
.Y(n_12174)
);

AND2x4_ASAP7_75t_L g12175 ( 
.A(n_11617),
.B(n_1485),
.Y(n_12175)
);

OA21x2_ASAP7_75t_L g12176 ( 
.A1(n_11545),
.A2(n_1486),
.B(n_1487),
.Y(n_12176)
);

INVxp33_ASAP7_75t_L g12177 ( 
.A(n_11464),
.Y(n_12177)
);

NAND2xp5_ASAP7_75t_L g12178 ( 
.A(n_11614),
.B(n_1486),
.Y(n_12178)
);

AND2x2_ASAP7_75t_SL g12179 ( 
.A(n_11545),
.B(n_1487),
.Y(n_12179)
);

INVx1_ASAP7_75t_L g12180 ( 
.A(n_11657),
.Y(n_12180)
);

OAI22xp5_ASAP7_75t_L g12181 ( 
.A1(n_11545),
.A2(n_1490),
.B1(n_1488),
.B2(n_1489),
.Y(n_12181)
);

OAI22xp5_ASAP7_75t_SL g12182 ( 
.A1(n_11625),
.A2(n_1490),
.B1(n_1488),
.B2(n_1489),
.Y(n_12182)
);

O2A1O1Ixp33_ASAP7_75t_L g12183 ( 
.A1(n_11509),
.A2(n_1491),
.B(n_1492),
.C(n_1490),
.Y(n_12183)
);

AOI21x1_ASAP7_75t_SL g12184 ( 
.A1(n_11457),
.A2(n_1489),
.B(n_1491),
.Y(n_12184)
);

INVx2_ASAP7_75t_L g12185 ( 
.A(n_11669),
.Y(n_12185)
);

AND2x2_ASAP7_75t_L g12186 ( 
.A(n_11545),
.B(n_1491),
.Y(n_12186)
);

NAND2xp5_ASAP7_75t_L g12187 ( 
.A(n_11614),
.B(n_1492),
.Y(n_12187)
);

OA21x2_ASAP7_75t_L g12188 ( 
.A1(n_11545),
.A2(n_1492),
.B(n_1493),
.Y(n_12188)
);

AOI21xp5_ASAP7_75t_L g12189 ( 
.A1(n_11476),
.A2(n_1493),
.B(n_1494),
.Y(n_12189)
);

AND2x4_ASAP7_75t_L g12190 ( 
.A(n_11617),
.B(n_1493),
.Y(n_12190)
);

O2A1O1Ixp5_ASAP7_75t_L g12191 ( 
.A1(n_11461),
.A2(n_1496),
.B(n_1494),
.C(n_1495),
.Y(n_12191)
);

OR2x2_ASAP7_75t_L g12192 ( 
.A(n_11567),
.B(n_1494),
.Y(n_12192)
);

OA21x2_ASAP7_75t_L g12193 ( 
.A1(n_11545),
.A2(n_1495),
.B(n_1496),
.Y(n_12193)
);

INVx1_ASAP7_75t_SL g12194 ( 
.A(n_11632),
.Y(n_12194)
);

OAI22xp5_ASAP7_75t_L g12195 ( 
.A1(n_11545),
.A2(n_1497),
.B1(n_1495),
.B2(n_1496),
.Y(n_12195)
);

AND2x2_ASAP7_75t_L g12196 ( 
.A(n_11545),
.B(n_1497),
.Y(n_12196)
);

INVx1_ASAP7_75t_L g12197 ( 
.A(n_11657),
.Y(n_12197)
);

AOI21xp5_ASAP7_75t_L g12198 ( 
.A1(n_11476),
.A2(n_1497),
.B(n_1498),
.Y(n_12198)
);

AND2x2_ASAP7_75t_L g12199 ( 
.A(n_11545),
.B(n_1498),
.Y(n_12199)
);

HB1xp67_ASAP7_75t_L g12200 ( 
.A(n_11607),
.Y(n_12200)
);

AND2x2_ASAP7_75t_L g12201 ( 
.A(n_11545),
.B(n_1498),
.Y(n_12201)
);

AOI21xp5_ASAP7_75t_L g12202 ( 
.A1(n_11476),
.A2(n_1499),
.B(n_1500),
.Y(n_12202)
);

HB1xp67_ASAP7_75t_L g12203 ( 
.A(n_11607),
.Y(n_12203)
);

BUFx12f_ASAP7_75t_L g12204 ( 
.A(n_11784),
.Y(n_12204)
);

NAND2xp5_ASAP7_75t_L g12205 ( 
.A(n_11614),
.B(n_1499),
.Y(n_12205)
);

A2O1A1Ixp33_ASAP7_75t_L g12206 ( 
.A1(n_11476),
.A2(n_1502),
.B(n_1500),
.C(n_1501),
.Y(n_12206)
);

INVx1_ASAP7_75t_L g12207 ( 
.A(n_11657),
.Y(n_12207)
);

AND2x2_ASAP7_75t_L g12208 ( 
.A(n_11545),
.B(n_1501),
.Y(n_12208)
);

INVx1_ASAP7_75t_L g12209 ( 
.A(n_11657),
.Y(n_12209)
);

BUFx3_ASAP7_75t_L g12210 ( 
.A(n_11632),
.Y(n_12210)
);

NAND2xp5_ASAP7_75t_L g12211 ( 
.A(n_11614),
.B(n_1502),
.Y(n_12211)
);

AND2x2_ASAP7_75t_L g12212 ( 
.A(n_11545),
.B(n_1502),
.Y(n_12212)
);

AND2x4_ASAP7_75t_L g12213 ( 
.A(n_11617),
.B(n_1503),
.Y(n_12213)
);

AND2x2_ASAP7_75t_L g12214 ( 
.A(n_11545),
.B(n_1504),
.Y(n_12214)
);

AND2x2_ASAP7_75t_L g12215 ( 
.A(n_11545),
.B(n_1504),
.Y(n_12215)
);

OA21x2_ASAP7_75t_L g12216 ( 
.A1(n_11545),
.A2(n_1504),
.B(n_1505),
.Y(n_12216)
);

AND2x2_ASAP7_75t_L g12217 ( 
.A(n_11545),
.B(n_1505),
.Y(n_12217)
);

BUFx6f_ASAP7_75t_L g12218 ( 
.A(n_11517),
.Y(n_12218)
);

NAND2xp5_ASAP7_75t_L g12219 ( 
.A(n_11614),
.B(n_1506),
.Y(n_12219)
);

OA21x2_ASAP7_75t_L g12220 ( 
.A1(n_11545),
.A2(n_1506),
.B(n_1507),
.Y(n_12220)
);

OAI22xp5_ASAP7_75t_L g12221 ( 
.A1(n_11545),
.A2(n_1508),
.B1(n_1506),
.B2(n_1507),
.Y(n_12221)
);

NAND2xp5_ASAP7_75t_L g12222 ( 
.A(n_11614),
.B(n_1508),
.Y(n_12222)
);

AOI21x1_ASAP7_75t_SL g12223 ( 
.A1(n_11457),
.A2(n_1508),
.B(n_1509),
.Y(n_12223)
);

AND2x4_ASAP7_75t_L g12224 ( 
.A(n_11617),
.B(n_1509),
.Y(n_12224)
);

BUFx2_ASAP7_75t_L g12225 ( 
.A(n_11632),
.Y(n_12225)
);

INVxp67_ASAP7_75t_SL g12226 ( 
.A(n_11575),
.Y(n_12226)
);

OR2x6_ASAP7_75t_L g12227 ( 
.A(n_12042),
.B(n_1510),
.Y(n_12227)
);

INVx1_ASAP7_75t_L g12228 ( 
.A(n_11848),
.Y(n_12228)
);

INVx1_ASAP7_75t_L g12229 ( 
.A(n_12151),
.Y(n_12229)
);

INVx3_ASAP7_75t_L g12230 ( 
.A(n_12218),
.Y(n_12230)
);

OAI21xp5_ASAP7_75t_L g12231 ( 
.A1(n_11911),
.A2(n_12105),
.B(n_11991),
.Y(n_12231)
);

AND2x4_ASAP7_75t_L g12232 ( 
.A(n_11949),
.B(n_1510),
.Y(n_12232)
);

OAI21x1_ASAP7_75t_L g12233 ( 
.A1(n_12013),
.A2(n_1511),
.B(n_1512),
.Y(n_12233)
);

INVx2_ASAP7_75t_L g12234 ( 
.A(n_12225),
.Y(n_12234)
);

INVx2_ASAP7_75t_L g12235 ( 
.A(n_12117),
.Y(n_12235)
);

OAI21xp5_ASAP7_75t_L g12236 ( 
.A1(n_11936),
.A2(n_1513),
.B(n_1512),
.Y(n_12236)
);

INVx1_ASAP7_75t_L g12237 ( 
.A(n_12163),
.Y(n_12237)
);

OAI21x1_ASAP7_75t_SL g12238 ( 
.A1(n_11863),
.A2(n_1511),
.B(n_1513),
.Y(n_12238)
);

INVx1_ASAP7_75t_L g12239 ( 
.A(n_12164),
.Y(n_12239)
);

INVx2_ASAP7_75t_L g12240 ( 
.A(n_12100),
.Y(n_12240)
);

INVx1_ASAP7_75t_L g12241 ( 
.A(n_12167),
.Y(n_12241)
);

INVx3_ASAP7_75t_L g12242 ( 
.A(n_12218),
.Y(n_12242)
);

AND2x2_ASAP7_75t_L g12243 ( 
.A(n_11823),
.B(n_1513),
.Y(n_12243)
);

INVx1_ASAP7_75t_L g12244 ( 
.A(n_12171),
.Y(n_12244)
);

AO21x2_ASAP7_75t_L g12245 ( 
.A1(n_12074),
.A2(n_1514),
.B(n_1515),
.Y(n_12245)
);

INVx1_ASAP7_75t_L g12246 ( 
.A(n_12180),
.Y(n_12246)
);

INVx1_ASAP7_75t_L g12247 ( 
.A(n_12197),
.Y(n_12247)
);

INVx1_ASAP7_75t_L g12248 ( 
.A(n_12207),
.Y(n_12248)
);

INVx1_ASAP7_75t_L g12249 ( 
.A(n_12209),
.Y(n_12249)
);

INVx1_ASAP7_75t_L g12250 ( 
.A(n_11825),
.Y(n_12250)
);

OAI21x1_ASAP7_75t_L g12251 ( 
.A1(n_11839),
.A2(n_1514),
.B(n_1515),
.Y(n_12251)
);

INVx1_ASAP7_75t_L g12252 ( 
.A(n_12155),
.Y(n_12252)
);

INVx1_ASAP7_75t_L g12253 ( 
.A(n_12158),
.Y(n_12253)
);

BUFx2_ASAP7_75t_L g12254 ( 
.A(n_11918),
.Y(n_12254)
);

INVx2_ASAP7_75t_L g12255 ( 
.A(n_12100),
.Y(n_12255)
);

AND2x2_ASAP7_75t_L g12256 ( 
.A(n_12066),
.B(n_1514),
.Y(n_12256)
);

INVx1_ASAP7_75t_L g12257 ( 
.A(n_12200),
.Y(n_12257)
);

INVx2_ASAP7_75t_L g12258 ( 
.A(n_12095),
.Y(n_12258)
);

INVx2_ASAP7_75t_L g12259 ( 
.A(n_12127),
.Y(n_12259)
);

NOR2x1_ASAP7_75t_R g12260 ( 
.A(n_12035),
.B(n_2441),
.Y(n_12260)
);

AND2x2_ASAP7_75t_L g12261 ( 
.A(n_12226),
.B(n_1516),
.Y(n_12261)
);

INVx1_ASAP7_75t_L g12262 ( 
.A(n_12203),
.Y(n_12262)
);

AND2x2_ASAP7_75t_L g12263 ( 
.A(n_11898),
.B(n_1516),
.Y(n_12263)
);

INVx2_ASAP7_75t_L g12264 ( 
.A(n_11969),
.Y(n_12264)
);

INVx3_ASAP7_75t_L g12265 ( 
.A(n_11882),
.Y(n_12265)
);

HB1xp67_ASAP7_75t_L g12266 ( 
.A(n_11892),
.Y(n_12266)
);

INVx2_ASAP7_75t_L g12267 ( 
.A(n_12055),
.Y(n_12267)
);

OAI21x1_ASAP7_75t_L g12268 ( 
.A1(n_11870),
.A2(n_1517),
.B(n_1518),
.Y(n_12268)
);

INVx1_ASAP7_75t_L g12269 ( 
.A(n_11934),
.Y(n_12269)
);

OA21x2_ASAP7_75t_L g12270 ( 
.A1(n_12096),
.A2(n_1517),
.B(n_1518),
.Y(n_12270)
);

INVx1_ASAP7_75t_L g12271 ( 
.A(n_11852),
.Y(n_12271)
);

INVx1_ASAP7_75t_L g12272 ( 
.A(n_11935),
.Y(n_12272)
);

INVx1_ASAP7_75t_L g12273 ( 
.A(n_11980),
.Y(n_12273)
);

OR2x2_ASAP7_75t_L g12274 ( 
.A(n_11902),
.B(n_1518),
.Y(n_12274)
);

AND2x2_ASAP7_75t_L g12275 ( 
.A(n_11832),
.B(n_12007),
.Y(n_12275)
);

INVx3_ASAP7_75t_L g12276 ( 
.A(n_11946),
.Y(n_12276)
);

INVx1_ASAP7_75t_L g12277 ( 
.A(n_12012),
.Y(n_12277)
);

BUFx3_ASAP7_75t_L g12278 ( 
.A(n_12204),
.Y(n_12278)
);

INVx1_ASAP7_75t_L g12279 ( 
.A(n_12017),
.Y(n_12279)
);

INVxp67_ASAP7_75t_L g12280 ( 
.A(n_12044),
.Y(n_12280)
);

INVx2_ASAP7_75t_L g12281 ( 
.A(n_11884),
.Y(n_12281)
);

OAI21x1_ASAP7_75t_L g12282 ( 
.A1(n_11836),
.A2(n_1519),
.B(n_1520),
.Y(n_12282)
);

INVx1_ASAP7_75t_L g12283 ( 
.A(n_12018),
.Y(n_12283)
);

AND2x2_ASAP7_75t_L g12284 ( 
.A(n_11850),
.B(n_1519),
.Y(n_12284)
);

INVx1_ASAP7_75t_L g12285 ( 
.A(n_11853),
.Y(n_12285)
);

INVx2_ASAP7_75t_L g12286 ( 
.A(n_12048),
.Y(n_12286)
);

INVx2_ASAP7_75t_L g12287 ( 
.A(n_11957),
.Y(n_12287)
);

OAI21x1_ASAP7_75t_L g12288 ( 
.A1(n_11833),
.A2(n_1519),
.B(n_1520),
.Y(n_12288)
);

INVx1_ASAP7_75t_L g12289 ( 
.A(n_11856),
.Y(n_12289)
);

INVx1_ASAP7_75t_L g12290 ( 
.A(n_11857),
.Y(n_12290)
);

INVx2_ASAP7_75t_L g12291 ( 
.A(n_12043),
.Y(n_12291)
);

NAND2xp5_ASAP7_75t_L g12292 ( 
.A(n_11943),
.B(n_1520),
.Y(n_12292)
);

NAND2xp5_ASAP7_75t_L g12293 ( 
.A(n_11897),
.B(n_1521),
.Y(n_12293)
);

INVx1_ASAP7_75t_L g12294 ( 
.A(n_11859),
.Y(n_12294)
);

INVx1_ASAP7_75t_L g12295 ( 
.A(n_11896),
.Y(n_12295)
);

INVx1_ASAP7_75t_L g12296 ( 
.A(n_11933),
.Y(n_12296)
);

NAND2xp5_ASAP7_75t_L g12297 ( 
.A(n_12072),
.B(n_1521),
.Y(n_12297)
);

INVx2_ASAP7_75t_L g12298 ( 
.A(n_12147),
.Y(n_12298)
);

AND2x2_ASAP7_75t_L g12299 ( 
.A(n_11845),
.B(n_1522),
.Y(n_12299)
);

INVx1_ASAP7_75t_L g12300 ( 
.A(n_12119),
.Y(n_12300)
);

INVx2_ASAP7_75t_L g12301 ( 
.A(n_11871),
.Y(n_12301)
);

OR2x6_ASAP7_75t_L g12302 ( 
.A(n_11874),
.B(n_1522),
.Y(n_12302)
);

INVx1_ASAP7_75t_L g12303 ( 
.A(n_12111),
.Y(n_12303)
);

INVx2_ASAP7_75t_L g12304 ( 
.A(n_12032),
.Y(n_12304)
);

INVx1_ASAP7_75t_L g12305 ( 
.A(n_12099),
.Y(n_12305)
);

INVx2_ASAP7_75t_L g12306 ( 
.A(n_11947),
.Y(n_12306)
);

AND2x2_ASAP7_75t_L g12307 ( 
.A(n_11820),
.B(n_1523),
.Y(n_12307)
);

INVx1_ASAP7_75t_L g12308 ( 
.A(n_12103),
.Y(n_12308)
);

INVx2_ASAP7_75t_L g12309 ( 
.A(n_11973),
.Y(n_12309)
);

AOI21x1_ASAP7_75t_L g12310 ( 
.A1(n_11948),
.A2(n_1523),
.B(n_1524),
.Y(n_12310)
);

INVx2_ASAP7_75t_L g12311 ( 
.A(n_11875),
.Y(n_12311)
);

BUFx3_ASAP7_75t_L g12312 ( 
.A(n_11819),
.Y(n_12312)
);

AND2x2_ASAP7_75t_L g12313 ( 
.A(n_11824),
.B(n_1523),
.Y(n_12313)
);

BUFx8_ASAP7_75t_L g12314 ( 
.A(n_11946),
.Y(n_12314)
);

INVx3_ASAP7_75t_L g12315 ( 
.A(n_12210),
.Y(n_12315)
);

BUFx2_ASAP7_75t_L g12316 ( 
.A(n_11919),
.Y(n_12316)
);

INVx2_ASAP7_75t_L g12317 ( 
.A(n_12057),
.Y(n_12317)
);

AO21x2_ASAP7_75t_L g12318 ( 
.A1(n_12109),
.A2(n_1524),
.B(n_1525),
.Y(n_12318)
);

AND2x2_ASAP7_75t_L g12319 ( 
.A(n_12160),
.B(n_1524),
.Y(n_12319)
);

AND2x2_ASAP7_75t_L g12320 ( 
.A(n_12186),
.B(n_1526),
.Y(n_12320)
);

BUFx6f_ASAP7_75t_L g12321 ( 
.A(n_11861),
.Y(n_12321)
);

INVxp33_ASAP7_75t_L g12322 ( 
.A(n_11821),
.Y(n_12322)
);

AO21x2_ASAP7_75t_L g12323 ( 
.A1(n_12079),
.A2(n_1526),
.B(n_1527),
.Y(n_12323)
);

INVx2_ASAP7_75t_L g12324 ( 
.A(n_11891),
.Y(n_12324)
);

AOI22xp33_ASAP7_75t_L g12325 ( 
.A1(n_12089),
.A2(n_1528),
.B1(n_1526),
.B2(n_1527),
.Y(n_12325)
);

INVx2_ASAP7_75t_L g12326 ( 
.A(n_12122),
.Y(n_12326)
);

INVx1_ASAP7_75t_L g12327 ( 
.A(n_12081),
.Y(n_12327)
);

INVx2_ASAP7_75t_L g12328 ( 
.A(n_12058),
.Y(n_12328)
);

OR2x2_ASAP7_75t_L g12329 ( 
.A(n_11883),
.B(n_1529),
.Y(n_12329)
);

AND2x4_ASAP7_75t_SL g12330 ( 
.A(n_11996),
.B(n_11981),
.Y(n_12330)
);

AOI22xp33_ASAP7_75t_L g12331 ( 
.A1(n_12092),
.A2(n_1531),
.B1(n_1529),
.B2(n_1530),
.Y(n_12331)
);

INVx2_ASAP7_75t_L g12332 ( 
.A(n_11905),
.Y(n_12332)
);

INVx2_ASAP7_75t_L g12333 ( 
.A(n_12011),
.Y(n_12333)
);

INVx2_ASAP7_75t_L g12334 ( 
.A(n_11860),
.Y(n_12334)
);

HB1xp67_ASAP7_75t_L g12335 ( 
.A(n_12170),
.Y(n_12335)
);

INVx3_ASAP7_75t_L g12336 ( 
.A(n_11981),
.Y(n_12336)
);

AND2x2_ASAP7_75t_L g12337 ( 
.A(n_12196),
.B(n_1529),
.Y(n_12337)
);

INVx2_ASAP7_75t_SL g12338 ( 
.A(n_11844),
.Y(n_12338)
);

INVx2_ASAP7_75t_L g12339 ( 
.A(n_12077),
.Y(n_12339)
);

INVx1_ASAP7_75t_L g12340 ( 
.A(n_12123),
.Y(n_12340)
);

OA21x2_ASAP7_75t_L g12341 ( 
.A1(n_12068),
.A2(n_1530),
.B(n_1531),
.Y(n_12341)
);

INVx2_ASAP7_75t_L g12342 ( 
.A(n_11841),
.Y(n_12342)
);

INVx2_ASAP7_75t_L g12343 ( 
.A(n_12125),
.Y(n_12343)
);

INVx1_ASAP7_75t_L g12344 ( 
.A(n_12041),
.Y(n_12344)
);

OA21x2_ASAP7_75t_L g12345 ( 
.A1(n_12091),
.A2(n_1531),
.B(n_1532),
.Y(n_12345)
);

INVx1_ASAP7_75t_L g12346 ( 
.A(n_12053),
.Y(n_12346)
);

BUFx12f_ASAP7_75t_L g12347 ( 
.A(n_11937),
.Y(n_12347)
);

AO21x2_ASAP7_75t_L g12348 ( 
.A1(n_11941),
.A2(n_1532),
.B(n_1533),
.Y(n_12348)
);

INVx1_ASAP7_75t_L g12349 ( 
.A(n_11993),
.Y(n_12349)
);

INVxp67_ASAP7_75t_SL g12350 ( 
.A(n_11988),
.Y(n_12350)
);

AND2x4_ASAP7_75t_L g12351 ( 
.A(n_12047),
.B(n_1533),
.Y(n_12351)
);

INVx1_ASAP7_75t_L g12352 ( 
.A(n_11990),
.Y(n_12352)
);

AND2x2_ASAP7_75t_L g12353 ( 
.A(n_12199),
.B(n_1533),
.Y(n_12353)
);

INVx3_ASAP7_75t_L g12354 ( 
.A(n_11877),
.Y(n_12354)
);

INVx1_ASAP7_75t_L g12355 ( 
.A(n_12010),
.Y(n_12355)
);

INVx1_ASAP7_75t_L g12356 ( 
.A(n_12070),
.Y(n_12356)
);

INVxp67_ASAP7_75t_L g12357 ( 
.A(n_12088),
.Y(n_12357)
);

INVx2_ASAP7_75t_L g12358 ( 
.A(n_12136),
.Y(n_12358)
);

AND2x4_ASAP7_75t_L g12359 ( 
.A(n_11842),
.B(n_1534),
.Y(n_12359)
);

INVx1_ASAP7_75t_L g12360 ( 
.A(n_12040),
.Y(n_12360)
);

OR2x2_ASAP7_75t_L g12361 ( 
.A(n_11889),
.B(n_1534),
.Y(n_12361)
);

INVx1_ASAP7_75t_L g12362 ( 
.A(n_12145),
.Y(n_12362)
);

AND2x2_ASAP7_75t_L g12363 ( 
.A(n_12201),
.B(n_12208),
.Y(n_12363)
);

NAND2xp5_ASAP7_75t_SL g12364 ( 
.A(n_11971),
.B(n_1534),
.Y(n_12364)
);

INVx1_ASAP7_75t_L g12365 ( 
.A(n_11829),
.Y(n_12365)
);

AND2x2_ASAP7_75t_L g12366 ( 
.A(n_12212),
.B(n_1535),
.Y(n_12366)
);

INVx2_ASAP7_75t_L g12367 ( 
.A(n_12056),
.Y(n_12367)
);

INVx1_ASAP7_75t_L g12368 ( 
.A(n_12192),
.Y(n_12368)
);

INVx2_ASAP7_75t_L g12369 ( 
.A(n_12059),
.Y(n_12369)
);

INVxp67_ASAP7_75t_L g12370 ( 
.A(n_12179),
.Y(n_12370)
);

AND2x2_ASAP7_75t_L g12371 ( 
.A(n_12214),
.B(n_1535),
.Y(n_12371)
);

INVx1_ASAP7_75t_L g12372 ( 
.A(n_12130),
.Y(n_12372)
);

OR2x6_ASAP7_75t_L g12373 ( 
.A(n_12083),
.B(n_1535),
.Y(n_12373)
);

INVxp67_ASAP7_75t_SL g12374 ( 
.A(n_12174),
.Y(n_12374)
);

INVx1_ASAP7_75t_L g12375 ( 
.A(n_12078),
.Y(n_12375)
);

INVx1_ASAP7_75t_L g12376 ( 
.A(n_12022),
.Y(n_12376)
);

INVx1_ASAP7_75t_L g12377 ( 
.A(n_12101),
.Y(n_12377)
);

INVx2_ASAP7_75t_L g12378 ( 
.A(n_12037),
.Y(n_12378)
);

INVx2_ASAP7_75t_L g12379 ( 
.A(n_12019),
.Y(n_12379)
);

INVxp67_ASAP7_75t_L g12380 ( 
.A(n_12176),
.Y(n_12380)
);

OAI21x1_ASAP7_75t_L g12381 ( 
.A1(n_12000),
.A2(n_1537),
.B(n_1538),
.Y(n_12381)
);

NAND2x1p5_ASAP7_75t_L g12382 ( 
.A(n_11873),
.B(n_1537),
.Y(n_12382)
);

INVx2_ASAP7_75t_L g12383 ( 
.A(n_11924),
.Y(n_12383)
);

NAND2xp5_ASAP7_75t_L g12384 ( 
.A(n_11940),
.B(n_1537),
.Y(n_12384)
);

AND2x4_ASAP7_75t_L g12385 ( 
.A(n_12021),
.B(n_1538),
.Y(n_12385)
);

INVx1_ASAP7_75t_L g12386 ( 
.A(n_11958),
.Y(n_12386)
);

INVx1_ASAP7_75t_L g12387 ( 
.A(n_11960),
.Y(n_12387)
);

AND2x2_ASAP7_75t_L g12388 ( 
.A(n_12215),
.B(n_1538),
.Y(n_12388)
);

AND2x2_ASAP7_75t_L g12389 ( 
.A(n_12217),
.B(n_1539),
.Y(n_12389)
);

AO31x2_ASAP7_75t_L g12390 ( 
.A1(n_11886),
.A2(n_1541),
.A3(n_1539),
.B(n_1540),
.Y(n_12390)
);

INVx1_ASAP7_75t_L g12391 ( 
.A(n_11962),
.Y(n_12391)
);

INVx2_ASAP7_75t_L g12392 ( 
.A(n_12061),
.Y(n_12392)
);

INVx1_ASAP7_75t_L g12393 ( 
.A(n_11927),
.Y(n_12393)
);

INVx2_ASAP7_75t_L g12394 ( 
.A(n_12094),
.Y(n_12394)
);

INVx1_ASAP7_75t_L g12395 ( 
.A(n_12133),
.Y(n_12395)
);

INVx1_ASAP7_75t_L g12396 ( 
.A(n_11866),
.Y(n_12396)
);

AND2x4_ASAP7_75t_L g12397 ( 
.A(n_11826),
.B(n_1540),
.Y(n_12397)
);

INVx2_ASAP7_75t_L g12398 ( 
.A(n_12065),
.Y(n_12398)
);

HB1xp67_ASAP7_75t_L g12399 ( 
.A(n_12188),
.Y(n_12399)
);

INVx1_ASAP7_75t_L g12400 ( 
.A(n_11822),
.Y(n_12400)
);

INVx2_ASAP7_75t_L g12401 ( 
.A(n_12139),
.Y(n_12401)
);

AND2x2_ASAP7_75t_L g12402 ( 
.A(n_12039),
.B(n_1540),
.Y(n_12402)
);

INVx1_ASAP7_75t_L g12403 ( 
.A(n_11835),
.Y(n_12403)
);

INVx2_ASAP7_75t_L g12404 ( 
.A(n_11890),
.Y(n_12404)
);

INVx3_ASAP7_75t_L g12405 ( 
.A(n_11855),
.Y(n_12405)
);

NOR2xp33_ASAP7_75t_L g12406 ( 
.A(n_12177),
.B(n_1541),
.Y(n_12406)
);

INVx1_ASAP7_75t_L g12407 ( 
.A(n_11837),
.Y(n_12407)
);

INVx3_ASAP7_75t_L g12408 ( 
.A(n_11901),
.Y(n_12408)
);

INVx2_ASAP7_75t_L g12409 ( 
.A(n_11915),
.Y(n_12409)
);

BUFx6f_ASAP7_75t_L g12410 ( 
.A(n_11966),
.Y(n_12410)
);

NAND2xp5_ASAP7_75t_L g12411 ( 
.A(n_11910),
.B(n_1542),
.Y(n_12411)
);

INVx2_ASAP7_75t_L g12412 ( 
.A(n_11977),
.Y(n_12412)
);

INVx2_ASAP7_75t_L g12413 ( 
.A(n_12129),
.Y(n_12413)
);

INVx2_ASAP7_75t_L g12414 ( 
.A(n_12175),
.Y(n_12414)
);

AO21x2_ASAP7_75t_L g12415 ( 
.A1(n_12073),
.A2(n_11876),
.B(n_11938),
.Y(n_12415)
);

INVx1_ASAP7_75t_L g12416 ( 
.A(n_11862),
.Y(n_12416)
);

OA21x2_ASAP7_75t_L g12417 ( 
.A1(n_12050),
.A2(n_1542),
.B(n_1543),
.Y(n_12417)
);

HB1xp67_ASAP7_75t_L g12418 ( 
.A(n_12193),
.Y(n_12418)
);

AND2x2_ASAP7_75t_L g12419 ( 
.A(n_12216),
.B(n_1542),
.Y(n_12419)
);

OR2x2_ASAP7_75t_L g12420 ( 
.A(n_11868),
.B(n_1543),
.Y(n_12420)
);

INVx2_ASAP7_75t_L g12421 ( 
.A(n_12190),
.Y(n_12421)
);

BUFx3_ASAP7_75t_L g12422 ( 
.A(n_11906),
.Y(n_12422)
);

INVx1_ASAP7_75t_L g12423 ( 
.A(n_12150),
.Y(n_12423)
);

OAI21x1_ASAP7_75t_L g12424 ( 
.A1(n_11830),
.A2(n_1544),
.B(n_1545),
.Y(n_12424)
);

OA21x2_ASAP7_75t_L g12425 ( 
.A1(n_12154),
.A2(n_1544),
.B(n_1545),
.Y(n_12425)
);

AND2x2_ASAP7_75t_L g12426 ( 
.A(n_12220),
.B(n_1544),
.Y(n_12426)
);

INVx2_ASAP7_75t_L g12427 ( 
.A(n_12213),
.Y(n_12427)
);

INVx1_ASAP7_75t_L g12428 ( 
.A(n_12159),
.Y(n_12428)
);

INVx2_ASAP7_75t_L g12429 ( 
.A(n_12224),
.Y(n_12429)
);

INVx1_ASAP7_75t_L g12430 ( 
.A(n_12178),
.Y(n_12430)
);

INVx1_ASAP7_75t_L g12431 ( 
.A(n_12187),
.Y(n_12431)
);

INVx2_ASAP7_75t_L g12432 ( 
.A(n_12107),
.Y(n_12432)
);

BUFx6f_ASAP7_75t_L g12433 ( 
.A(n_11972),
.Y(n_12433)
);

INVx2_ASAP7_75t_L g12434 ( 
.A(n_11907),
.Y(n_12434)
);

INVx1_ASAP7_75t_L g12435 ( 
.A(n_12205),
.Y(n_12435)
);

INVx1_ASAP7_75t_L g12436 ( 
.A(n_12211),
.Y(n_12436)
);

AO21x2_ASAP7_75t_L g12437 ( 
.A1(n_12219),
.A2(n_12222),
.B(n_11864),
.Y(n_12437)
);

INVx2_ASAP7_75t_L g12438 ( 
.A(n_11923),
.Y(n_12438)
);

INVx4_ASAP7_75t_SL g12439 ( 
.A(n_11843),
.Y(n_12439)
);

NOR2xp33_ASAP7_75t_L g12440 ( 
.A(n_11869),
.B(n_1546),
.Y(n_12440)
);

INVx1_ASAP7_75t_L g12441 ( 
.A(n_11945),
.Y(n_12441)
);

AO21x2_ASAP7_75t_L g12442 ( 
.A1(n_12029),
.A2(n_1546),
.B(n_1547),
.Y(n_12442)
);

INVx1_ASAP7_75t_L g12443 ( 
.A(n_11878),
.Y(n_12443)
);

OA21x2_ASAP7_75t_L g12444 ( 
.A1(n_12156),
.A2(n_1546),
.B(n_1547),
.Y(n_12444)
);

BUFx3_ASAP7_75t_L g12445 ( 
.A(n_12002),
.Y(n_12445)
);

AND2x2_ASAP7_75t_L g12446 ( 
.A(n_11998),
.B(n_1548),
.Y(n_12446)
);

INVx2_ASAP7_75t_L g12447 ( 
.A(n_11838),
.Y(n_12447)
);

INVx2_ASAP7_75t_L g12448 ( 
.A(n_12062),
.Y(n_12448)
);

INVx2_ASAP7_75t_SL g12449 ( 
.A(n_12064),
.Y(n_12449)
);

OAI21x1_ASAP7_75t_L g12450 ( 
.A1(n_12185),
.A2(n_1548),
.B(n_1549),
.Y(n_12450)
);

INVx1_ASAP7_75t_L g12451 ( 
.A(n_11954),
.Y(n_12451)
);

HB1xp67_ASAP7_75t_L g12452 ( 
.A(n_12084),
.Y(n_12452)
);

BUFx2_ASAP7_75t_L g12453 ( 
.A(n_12085),
.Y(n_12453)
);

OAI21x1_ASAP7_75t_L g12454 ( 
.A1(n_11955),
.A2(n_1548),
.B(n_1549),
.Y(n_12454)
);

BUFx3_ASAP7_75t_L g12455 ( 
.A(n_11984),
.Y(n_12455)
);

INVx2_ASAP7_75t_L g12456 ( 
.A(n_12082),
.Y(n_12456)
);

AND2x2_ASAP7_75t_L g12457 ( 
.A(n_11846),
.B(n_1549),
.Y(n_12457)
);

BUFx2_ASAP7_75t_L g12458 ( 
.A(n_11956),
.Y(n_12458)
);

OR2x2_ASAP7_75t_L g12459 ( 
.A(n_11970),
.B(n_1550),
.Y(n_12459)
);

HB1xp67_ASAP7_75t_L g12460 ( 
.A(n_11881),
.Y(n_12460)
);

NAND2xp5_ASAP7_75t_SL g12461 ( 
.A(n_12152),
.B(n_1550),
.Y(n_12461)
);

INVx1_ASAP7_75t_L g12462 ( 
.A(n_11979),
.Y(n_12462)
);

INVx1_ASAP7_75t_L g12463 ( 
.A(n_11994),
.Y(n_12463)
);

BUFx2_ASAP7_75t_L g12464 ( 
.A(n_12194),
.Y(n_12464)
);

INVx3_ASAP7_75t_L g12465 ( 
.A(n_11847),
.Y(n_12465)
);

INVx2_ASAP7_75t_L g12466 ( 
.A(n_12097),
.Y(n_12466)
);

AND2x4_ASAP7_75t_L g12467 ( 
.A(n_11849),
.B(n_1550),
.Y(n_12467)
);

AND2x4_ASAP7_75t_SL g12468 ( 
.A(n_11899),
.B(n_1551),
.Y(n_12468)
);

AND2x2_ASAP7_75t_L g12469 ( 
.A(n_11931),
.B(n_1551),
.Y(n_12469)
);

NAND2xp5_ASAP7_75t_L g12470 ( 
.A(n_12076),
.B(n_1552),
.Y(n_12470)
);

OA21x2_ASAP7_75t_L g12471 ( 
.A1(n_11950),
.A2(n_1552),
.B(n_1553),
.Y(n_12471)
);

HB1xp67_ASAP7_75t_L g12472 ( 
.A(n_11997),
.Y(n_12472)
);

AND2x4_ASAP7_75t_L g12473 ( 
.A(n_11854),
.B(n_1554),
.Y(n_12473)
);

OAI21x1_ASAP7_75t_L g12474 ( 
.A1(n_11976),
.A2(n_1554),
.B(n_1556),
.Y(n_12474)
);

INVx1_ASAP7_75t_L g12475 ( 
.A(n_12033),
.Y(n_12475)
);

INVx1_ASAP7_75t_L g12476 ( 
.A(n_11893),
.Y(n_12476)
);

INVx1_ASAP7_75t_L g12477 ( 
.A(n_11908),
.Y(n_12477)
);

INVx1_ASAP7_75t_L g12478 ( 
.A(n_11909),
.Y(n_12478)
);

NAND2xp5_ASAP7_75t_L g12479 ( 
.A(n_12020),
.B(n_1554),
.Y(n_12479)
);

INVx2_ASAP7_75t_L g12480 ( 
.A(n_11858),
.Y(n_12480)
);

INVx1_ASAP7_75t_L g12481 ( 
.A(n_12138),
.Y(n_12481)
);

INVx1_ASAP7_75t_L g12482 ( 
.A(n_12132),
.Y(n_12482)
);

INVx1_ASAP7_75t_L g12483 ( 
.A(n_11985),
.Y(n_12483)
);

HB1xp67_ASAP7_75t_L g12484 ( 
.A(n_12120),
.Y(n_12484)
);

AO21x2_ASAP7_75t_L g12485 ( 
.A1(n_11952),
.A2(n_11939),
.B(n_12001),
.Y(n_12485)
);

OAI21x1_ASAP7_75t_L g12486 ( 
.A1(n_12110),
.A2(n_1556),
.B(n_1557),
.Y(n_12486)
);

HB1xp67_ASAP7_75t_L g12487 ( 
.A(n_12014),
.Y(n_12487)
);

INVx3_ASAP7_75t_L g12488 ( 
.A(n_12104),
.Y(n_12488)
);

INVx1_ASAP7_75t_L g12489 ( 
.A(n_11989),
.Y(n_12489)
);

CKINVDCx5p33_ASAP7_75t_R g12490 ( 
.A(n_11895),
.Y(n_12490)
);

NAND2xp5_ASAP7_75t_L g12491 ( 
.A(n_11978),
.B(n_1557),
.Y(n_12491)
);

INVx2_ASAP7_75t_SL g12492 ( 
.A(n_12015),
.Y(n_12492)
);

INVx2_ASAP7_75t_L g12493 ( 
.A(n_11879),
.Y(n_12493)
);

OA21x2_ASAP7_75t_L g12494 ( 
.A1(n_11885),
.A2(n_1557),
.B(n_1558),
.Y(n_12494)
);

AO21x2_ASAP7_75t_L g12495 ( 
.A1(n_11903),
.A2(n_1558),
.B(n_1559),
.Y(n_12495)
);

HB1xp67_ASAP7_75t_L g12496 ( 
.A(n_12038),
.Y(n_12496)
);

NAND2xp5_ASAP7_75t_L g12497 ( 
.A(n_11983),
.B(n_1559),
.Y(n_12497)
);

INVx1_ASAP7_75t_L g12498 ( 
.A(n_12034),
.Y(n_12498)
);

INVx2_ASAP7_75t_L g12499 ( 
.A(n_12054),
.Y(n_12499)
);

HB1xp67_ASAP7_75t_L g12500 ( 
.A(n_12045),
.Y(n_12500)
);

HB1xp67_ASAP7_75t_L g12501 ( 
.A(n_11872),
.Y(n_12501)
);

BUFx3_ASAP7_75t_L g12502 ( 
.A(n_12049),
.Y(n_12502)
);

INVx1_ASAP7_75t_L g12503 ( 
.A(n_12093),
.Y(n_12503)
);

INVx2_ASAP7_75t_L g12504 ( 
.A(n_12146),
.Y(n_12504)
);

INVx1_ASAP7_75t_L g12505 ( 
.A(n_11904),
.Y(n_12505)
);

OR2x2_ASAP7_75t_L g12506 ( 
.A(n_11887),
.B(n_12028),
.Y(n_12506)
);

INVx3_ASAP7_75t_L g12507 ( 
.A(n_12098),
.Y(n_12507)
);

AOI22xp33_ASAP7_75t_L g12508 ( 
.A1(n_11928),
.A2(n_1562),
.B1(n_1560),
.B2(n_1561),
.Y(n_12508)
);

INVxp67_ASAP7_75t_L g12509 ( 
.A(n_11925),
.Y(n_12509)
);

INVx2_ASAP7_75t_L g12510 ( 
.A(n_12116),
.Y(n_12510)
);

OA21x2_ASAP7_75t_L g12511 ( 
.A1(n_12052),
.A2(n_1560),
.B(n_1562),
.Y(n_12511)
);

AO21x2_ASAP7_75t_L g12512 ( 
.A1(n_12114),
.A2(n_1560),
.B(n_1563),
.Y(n_12512)
);

HB1xp67_ASAP7_75t_L g12513 ( 
.A(n_12036),
.Y(n_12513)
);

AND2x2_ASAP7_75t_SL g12514 ( 
.A(n_11867),
.B(n_1563),
.Y(n_12514)
);

INVx2_ASAP7_75t_L g12515 ( 
.A(n_12071),
.Y(n_12515)
);

AO21x1_ASAP7_75t_SL g12516 ( 
.A1(n_11953),
.A2(n_1563),
.B(n_1564),
.Y(n_12516)
);

INVx1_ASAP7_75t_L g12517 ( 
.A(n_11913),
.Y(n_12517)
);

INVx1_ASAP7_75t_L g12518 ( 
.A(n_11920),
.Y(n_12518)
);

AND2x2_ASAP7_75t_L g12519 ( 
.A(n_12006),
.B(n_1564),
.Y(n_12519)
);

OAI21xp5_ASAP7_75t_L g12520 ( 
.A1(n_12191),
.A2(n_1567),
.B(n_1566),
.Y(n_12520)
);

OAI21x1_ASAP7_75t_L g12521 ( 
.A1(n_12086),
.A2(n_1565),
.B(n_1566),
.Y(n_12521)
);

INVx2_ASAP7_75t_L g12522 ( 
.A(n_12080),
.Y(n_12522)
);

INVx2_ASAP7_75t_L g12523 ( 
.A(n_11951),
.Y(n_12523)
);

INVx2_ASAP7_75t_L g12524 ( 
.A(n_12113),
.Y(n_12524)
);

OAI21x1_ASAP7_75t_L g12525 ( 
.A1(n_11827),
.A2(n_1565),
.B(n_1567),
.Y(n_12525)
);

INVx1_ASAP7_75t_L g12526 ( 
.A(n_12137),
.Y(n_12526)
);

INVx1_ASAP7_75t_L g12527 ( 
.A(n_12143),
.Y(n_12527)
);

INVx1_ASAP7_75t_L g12528 ( 
.A(n_12046),
.Y(n_12528)
);

BUFx6f_ASAP7_75t_L g12529 ( 
.A(n_12024),
.Y(n_12529)
);

INVx2_ASAP7_75t_L g12530 ( 
.A(n_12121),
.Y(n_12530)
);

INVx3_ASAP7_75t_L g12531 ( 
.A(n_12009),
.Y(n_12531)
);

INVx2_ASAP7_75t_L g12532 ( 
.A(n_11900),
.Y(n_12532)
);

HB1xp67_ASAP7_75t_L g12533 ( 
.A(n_12162),
.Y(n_12533)
);

INVx2_ASAP7_75t_L g12534 ( 
.A(n_11916),
.Y(n_12534)
);

OAI22xp5_ASAP7_75t_L g12535 ( 
.A1(n_12172),
.A2(n_1568),
.B1(n_1565),
.B2(n_1567),
.Y(n_12535)
);

INVx3_ASAP7_75t_L g12536 ( 
.A(n_12090),
.Y(n_12536)
);

INVx2_ASAP7_75t_L g12537 ( 
.A(n_11888),
.Y(n_12537)
);

AND2x2_ASAP7_75t_L g12538 ( 
.A(n_12165),
.B(n_1569),
.Y(n_12538)
);

INVxp67_ASAP7_75t_SL g12539 ( 
.A(n_11894),
.Y(n_12539)
);

INVx1_ASAP7_75t_L g12540 ( 
.A(n_12115),
.Y(n_12540)
);

INVx2_ASAP7_75t_L g12541 ( 
.A(n_11987),
.Y(n_12541)
);

AND2x2_ASAP7_75t_L g12542 ( 
.A(n_12169),
.B(n_1569),
.Y(n_12542)
);

AND2x2_ASAP7_75t_L g12543 ( 
.A(n_12181),
.B(n_1570),
.Y(n_12543)
);

INVx2_ASAP7_75t_L g12544 ( 
.A(n_12003),
.Y(n_12544)
);

INVx1_ASAP7_75t_L g12545 ( 
.A(n_12142),
.Y(n_12545)
);

OAI21xp5_ASAP7_75t_L g12546 ( 
.A1(n_12189),
.A2(n_1572),
.B(n_1571),
.Y(n_12546)
);

OAI22xp33_ASAP7_75t_L g12547 ( 
.A1(n_11992),
.A2(n_1580),
.B1(n_1588),
.B2(n_1570),
.Y(n_12547)
);

INVx2_ASAP7_75t_L g12548 ( 
.A(n_12008),
.Y(n_12548)
);

INVx1_ASAP7_75t_L g12549 ( 
.A(n_11961),
.Y(n_12549)
);

INVx2_ASAP7_75t_L g12550 ( 
.A(n_12051),
.Y(n_12550)
);

INVx2_ASAP7_75t_L g12551 ( 
.A(n_12126),
.Y(n_12551)
);

INVxp67_ASAP7_75t_L g12552 ( 
.A(n_12063),
.Y(n_12552)
);

INVx2_ASAP7_75t_L g12553 ( 
.A(n_11914),
.Y(n_12553)
);

OR2x6_ASAP7_75t_L g12554 ( 
.A(n_11831),
.B(n_1570),
.Y(n_12554)
);

INVx2_ASAP7_75t_L g12555 ( 
.A(n_11921),
.Y(n_12555)
);

INVx3_ASAP7_75t_L g12556 ( 
.A(n_11880),
.Y(n_12556)
);

INVx1_ASAP7_75t_L g12557 ( 
.A(n_11964),
.Y(n_12557)
);

AND2x4_ASAP7_75t_L g12558 ( 
.A(n_12141),
.B(n_1571),
.Y(n_12558)
);

INVx2_ASAP7_75t_L g12559 ( 
.A(n_12135),
.Y(n_12559)
);

NAND2xp5_ASAP7_75t_L g12560 ( 
.A(n_12023),
.B(n_1573),
.Y(n_12560)
);

INVx2_ASAP7_75t_L g12561 ( 
.A(n_11917),
.Y(n_12561)
);

NOR2xp33_ASAP7_75t_L g12562 ( 
.A(n_11968),
.B(n_1573),
.Y(n_12562)
);

INVx1_ASAP7_75t_L g12563 ( 
.A(n_11995),
.Y(n_12563)
);

AND2x2_ASAP7_75t_L g12564 ( 
.A(n_12195),
.B(n_1575),
.Y(n_12564)
);

INVx2_ASAP7_75t_L g12565 ( 
.A(n_12004),
.Y(n_12565)
);

INVx1_ASAP7_75t_L g12566 ( 
.A(n_12025),
.Y(n_12566)
);

INVx1_ASAP7_75t_L g12567 ( 
.A(n_12112),
.Y(n_12567)
);

INVx1_ASAP7_75t_L g12568 ( 
.A(n_12124),
.Y(n_12568)
);

OR2x2_ASAP7_75t_L g12569 ( 
.A(n_12027),
.B(n_1575),
.Y(n_12569)
);

INVx2_ASAP7_75t_SL g12570 ( 
.A(n_11828),
.Y(n_12570)
);

AND2x2_ASAP7_75t_L g12571 ( 
.A(n_12221),
.B(n_11929),
.Y(n_12571)
);

HB1xp67_ASAP7_75t_L g12572 ( 
.A(n_12069),
.Y(n_12572)
);

INVx2_ASAP7_75t_L g12573 ( 
.A(n_12087),
.Y(n_12573)
);

INVx1_ASAP7_75t_L g12574 ( 
.A(n_12134),
.Y(n_12574)
);

INVx3_ASAP7_75t_L g12575 ( 
.A(n_11840),
.Y(n_12575)
);

OAI21x1_ASAP7_75t_L g12576 ( 
.A1(n_12161),
.A2(n_1576),
.B(n_1577),
.Y(n_12576)
);

INVx2_ASAP7_75t_L g12577 ( 
.A(n_12005),
.Y(n_12577)
);

OR2x2_ASAP7_75t_L g12578 ( 
.A(n_11922),
.B(n_1576),
.Y(n_12578)
);

INVx1_ASAP7_75t_L g12579 ( 
.A(n_12148),
.Y(n_12579)
);

BUFx3_ASAP7_75t_L g12580 ( 
.A(n_12182),
.Y(n_12580)
);

INVx1_ASAP7_75t_L g12581 ( 
.A(n_12108),
.Y(n_12581)
);

INVx2_ASAP7_75t_L g12582 ( 
.A(n_12026),
.Y(n_12582)
);

OAI21xp5_ASAP7_75t_L g12583 ( 
.A1(n_12198),
.A2(n_1578),
.B(n_1577),
.Y(n_12583)
);

AND2x2_ASAP7_75t_L g12584 ( 
.A(n_12202),
.B(n_1576),
.Y(n_12584)
);

INVx1_ASAP7_75t_L g12585 ( 
.A(n_12153),
.Y(n_12585)
);

NAND2xp5_ASAP7_75t_L g12586 ( 
.A(n_12166),
.B(n_1578),
.Y(n_12586)
);

NOR2xp33_ASAP7_75t_L g12587 ( 
.A(n_12157),
.B(n_1578),
.Y(n_12587)
);

INVx1_ASAP7_75t_L g12588 ( 
.A(n_12183),
.Y(n_12588)
);

INVx2_ASAP7_75t_L g12589 ( 
.A(n_12102),
.Y(n_12589)
);

INVx2_ASAP7_75t_L g12590 ( 
.A(n_12060),
.Y(n_12590)
);

AO21x1_ASAP7_75t_SL g12591 ( 
.A1(n_11944),
.A2(n_1579),
.B(n_1580),
.Y(n_12591)
);

AOI21xp33_ASAP7_75t_L g12592 ( 
.A1(n_11959),
.A2(n_2438),
.B(n_2437),
.Y(n_12592)
);

INVx1_ASAP7_75t_L g12593 ( 
.A(n_12016),
.Y(n_12593)
);

AND2x2_ASAP7_75t_L g12594 ( 
.A(n_12030),
.B(n_1579),
.Y(n_12594)
);

INVx1_ASAP7_75t_L g12595 ( 
.A(n_11834),
.Y(n_12595)
);

AOI22xp5_ASAP7_75t_L g12596 ( 
.A1(n_12173),
.A2(n_11926),
.B1(n_11942),
.B2(n_11932),
.Y(n_12596)
);

INVx2_ASAP7_75t_L g12597 ( 
.A(n_12184),
.Y(n_12597)
);

OR2x2_ASAP7_75t_L g12598 ( 
.A(n_12149),
.B(n_1581),
.Y(n_12598)
);

CKINVDCx20_ASAP7_75t_R g12599 ( 
.A(n_11974),
.Y(n_12599)
);

INVx1_ASAP7_75t_L g12600 ( 
.A(n_12206),
.Y(n_12600)
);

INVx1_ASAP7_75t_L g12601 ( 
.A(n_12128),
.Y(n_12601)
);

OAI21x1_ASAP7_75t_L g12602 ( 
.A1(n_12223),
.A2(n_1581),
.B(n_1582),
.Y(n_12602)
);

INVx1_ASAP7_75t_L g12603 ( 
.A(n_11975),
.Y(n_12603)
);

AO21x2_ASAP7_75t_L g12604 ( 
.A1(n_11963),
.A2(n_12140),
.B(n_11967),
.Y(n_12604)
);

INVx2_ASAP7_75t_L g12605 ( 
.A(n_11851),
.Y(n_12605)
);

INVx1_ASAP7_75t_L g12606 ( 
.A(n_12031),
.Y(n_12606)
);

INVx1_ASAP7_75t_L g12607 ( 
.A(n_11982),
.Y(n_12607)
);

NAND2xp5_ASAP7_75t_SL g12608 ( 
.A(n_12168),
.B(n_1581),
.Y(n_12608)
);

INVx3_ASAP7_75t_L g12609 ( 
.A(n_11965),
.Y(n_12609)
);

BUFx2_ASAP7_75t_L g12610 ( 
.A(n_11865),
.Y(n_12610)
);

INVx1_ASAP7_75t_L g12611 ( 
.A(n_11999),
.Y(n_12611)
);

BUFx2_ASAP7_75t_SL g12612 ( 
.A(n_11986),
.Y(n_12612)
);

INVx2_ASAP7_75t_L g12613 ( 
.A(n_12075),
.Y(n_12613)
);

INVx1_ASAP7_75t_L g12614 ( 
.A(n_12118),
.Y(n_12614)
);

INVx2_ASAP7_75t_L g12615 ( 
.A(n_11912),
.Y(n_12615)
);

AO21x2_ASAP7_75t_L g12616 ( 
.A1(n_11930),
.A2(n_1582),
.B(n_1583),
.Y(n_12616)
);

INVx2_ASAP7_75t_L g12617 ( 
.A(n_12067),
.Y(n_12617)
);

AND2x2_ASAP7_75t_L g12618 ( 
.A(n_12106),
.B(n_1583),
.Y(n_12618)
);

HB1xp67_ASAP7_75t_L g12619 ( 
.A(n_12144),
.Y(n_12619)
);

OAI21x1_ASAP7_75t_L g12620 ( 
.A1(n_12131),
.A2(n_1583),
.B(n_1584),
.Y(n_12620)
);

INVx2_ASAP7_75t_L g12621 ( 
.A(n_12225),
.Y(n_12621)
);

AND2x2_ASAP7_75t_L g12622 ( 
.A(n_11823),
.B(n_1585),
.Y(n_12622)
);

INVx1_ASAP7_75t_L g12623 ( 
.A(n_11848),
.Y(n_12623)
);

OAI21x1_ASAP7_75t_L g12624 ( 
.A1(n_12013),
.A2(n_1585),
.B(n_1586),
.Y(n_12624)
);

NAND2xp5_ASAP7_75t_L g12625 ( 
.A(n_12226),
.B(n_1585),
.Y(n_12625)
);

CKINVDCx16_ASAP7_75t_R g12626 ( 
.A(n_12204),
.Y(n_12626)
);

NAND2xp5_ASAP7_75t_L g12627 ( 
.A(n_12226),
.B(n_1586),
.Y(n_12627)
);

INVx2_ASAP7_75t_L g12628 ( 
.A(n_12225),
.Y(n_12628)
);

INVx3_ASAP7_75t_L g12629 ( 
.A(n_12218),
.Y(n_12629)
);

NAND2xp5_ASAP7_75t_L g12630 ( 
.A(n_12226),
.B(n_1586),
.Y(n_12630)
);

INVx1_ASAP7_75t_L g12631 ( 
.A(n_11848),
.Y(n_12631)
);

INVx1_ASAP7_75t_L g12632 ( 
.A(n_11848),
.Y(n_12632)
);

INVx1_ASAP7_75t_L g12633 ( 
.A(n_11848),
.Y(n_12633)
);

INVx2_ASAP7_75t_L g12634 ( 
.A(n_12225),
.Y(n_12634)
);

OR2x2_ASAP7_75t_SL g12635 ( 
.A(n_12170),
.B(n_1587),
.Y(n_12635)
);

INVx5_ASAP7_75t_L g12636 ( 
.A(n_12204),
.Y(n_12636)
);

INVx1_ASAP7_75t_L g12637 ( 
.A(n_11848),
.Y(n_12637)
);

AO21x2_ASAP7_75t_L g12638 ( 
.A1(n_12074),
.A2(n_1587),
.B(n_1588),
.Y(n_12638)
);

OR2x2_ASAP7_75t_L g12639 ( 
.A(n_12226),
.B(n_1587),
.Y(n_12639)
);

AOI21x1_ASAP7_75t_L g12640 ( 
.A1(n_12042),
.A2(n_1589),
.B(n_1590),
.Y(n_12640)
);

INVx1_ASAP7_75t_L g12641 ( 
.A(n_11848),
.Y(n_12641)
);

INVx2_ASAP7_75t_L g12642 ( 
.A(n_12225),
.Y(n_12642)
);

AND2x2_ASAP7_75t_L g12643 ( 
.A(n_11823),
.B(n_1589),
.Y(n_12643)
);

INVx1_ASAP7_75t_L g12644 ( 
.A(n_11848),
.Y(n_12644)
);

AOI21xp5_ASAP7_75t_L g12645 ( 
.A1(n_11911),
.A2(n_2452),
.B(n_2451),
.Y(n_12645)
);

INVx2_ASAP7_75t_L g12646 ( 
.A(n_12225),
.Y(n_12646)
);

BUFx2_ASAP7_75t_L g12647 ( 
.A(n_11918),
.Y(n_12647)
);

HB1xp67_ASAP7_75t_L g12648 ( 
.A(n_11892),
.Y(n_12648)
);

NAND2x1p5_ASAP7_75t_L g12649 ( 
.A(n_11873),
.B(n_1589),
.Y(n_12649)
);

OAI21x1_ASAP7_75t_L g12650 ( 
.A1(n_12013),
.A2(n_1590),
.B(n_1591),
.Y(n_12650)
);

AND2x2_ASAP7_75t_L g12651 ( 
.A(n_11823),
.B(n_1590),
.Y(n_12651)
);

INVx2_ASAP7_75t_L g12652 ( 
.A(n_12225),
.Y(n_12652)
);

AO21x2_ASAP7_75t_L g12653 ( 
.A1(n_12074),
.A2(n_1591),
.B(n_1592),
.Y(n_12653)
);

INVx1_ASAP7_75t_L g12654 ( 
.A(n_11848),
.Y(n_12654)
);

INVxp67_ASAP7_75t_L g12655 ( 
.A(n_11823),
.Y(n_12655)
);

AO21x2_ASAP7_75t_L g12656 ( 
.A1(n_12074),
.A2(n_1592),
.B(n_1593),
.Y(n_12656)
);

NOR2xp67_ASAP7_75t_L g12657 ( 
.A(n_12347),
.B(n_2433),
.Y(n_12657)
);

INVxp67_ASAP7_75t_L g12658 ( 
.A(n_12260),
.Y(n_12658)
);

NOR2xp33_ASAP7_75t_SL g12659 ( 
.A(n_12316),
.B(n_1593),
.Y(n_12659)
);

BUFx3_ASAP7_75t_L g12660 ( 
.A(n_12314),
.Y(n_12660)
);

NAND2x1_ASAP7_75t_L g12661 ( 
.A(n_12275),
.B(n_1592),
.Y(n_12661)
);

NOR2xp33_ASAP7_75t_L g12662 ( 
.A(n_12626),
.B(n_1593),
.Y(n_12662)
);

NAND2xp5_ASAP7_75t_L g12663 ( 
.A(n_12374),
.B(n_1594),
.Y(n_12663)
);

NAND2xp5_ASAP7_75t_L g12664 ( 
.A(n_12335),
.B(n_1594),
.Y(n_12664)
);

BUFx2_ASAP7_75t_L g12665 ( 
.A(n_12453),
.Y(n_12665)
);

A2O1A1Ixp33_ASAP7_75t_L g12666 ( 
.A1(n_12231),
.A2(n_1596),
.B(n_1597),
.C(n_1595),
.Y(n_12666)
);

NOR2x1_ASAP7_75t_SL g12667 ( 
.A(n_12516),
.B(n_12591),
.Y(n_12667)
);

INVx1_ASAP7_75t_L g12668 ( 
.A(n_12487),
.Y(n_12668)
);

OAI22xp5_ASAP7_75t_L g12669 ( 
.A1(n_12655),
.A2(n_1596),
.B1(n_1594),
.B2(n_1595),
.Y(n_12669)
);

INVx2_ASAP7_75t_L g12670 ( 
.A(n_12312),
.Y(n_12670)
);

NOR2xp33_ASAP7_75t_L g12671 ( 
.A(n_12636),
.B(n_1595),
.Y(n_12671)
);

AND2x2_ASAP7_75t_L g12672 ( 
.A(n_12464),
.B(n_1596),
.Y(n_12672)
);

AND2x2_ASAP7_75t_L g12673 ( 
.A(n_12258),
.B(n_1597),
.Y(n_12673)
);

AOI221xp5_ASAP7_75t_L g12674 ( 
.A1(n_12484),
.A2(n_1599),
.B1(n_1597),
.B2(n_1598),
.C(n_1600),
.Y(n_12674)
);

AND2x2_ASAP7_75t_L g12675 ( 
.A(n_12363),
.B(n_1598),
.Y(n_12675)
);

AO32x2_ASAP7_75t_L g12676 ( 
.A1(n_12492),
.A2(n_1601),
.A3(n_1599),
.B1(n_1600),
.B2(n_1602),
.Y(n_12676)
);

AND2x2_ASAP7_75t_L g12677 ( 
.A(n_12254),
.B(n_1600),
.Y(n_12677)
);

AOI221xp5_ASAP7_75t_L g12678 ( 
.A1(n_12380),
.A2(n_1603),
.B1(n_1601),
.B2(n_1602),
.C(n_1604),
.Y(n_12678)
);

AND2x2_ASAP7_75t_L g12679 ( 
.A(n_12647),
.B(n_1601),
.Y(n_12679)
);

AND2x2_ASAP7_75t_L g12680 ( 
.A(n_12394),
.B(n_1603),
.Y(n_12680)
);

AND2x2_ASAP7_75t_L g12681 ( 
.A(n_12256),
.B(n_1603),
.Y(n_12681)
);

INVx2_ASAP7_75t_L g12682 ( 
.A(n_12502),
.Y(n_12682)
);

AND2x2_ASAP7_75t_L g12683 ( 
.A(n_12405),
.B(n_1604),
.Y(n_12683)
);

A2O1A1Ixp33_ASAP7_75t_L g12684 ( 
.A1(n_12645),
.A2(n_1606),
.B(n_1607),
.C(n_1605),
.Y(n_12684)
);

A2O1A1Ixp33_ASAP7_75t_L g12685 ( 
.A1(n_12236),
.A2(n_1606),
.B(n_1607),
.C(n_1605),
.Y(n_12685)
);

INVx3_ASAP7_75t_L g12686 ( 
.A(n_12278),
.Y(n_12686)
);

OAI22xp5_ASAP7_75t_SL g12687 ( 
.A1(n_12599),
.A2(n_12552),
.B1(n_12539),
.B2(n_12501),
.Y(n_12687)
);

OR2x2_ASAP7_75t_L g12688 ( 
.A(n_12472),
.B(n_1604),
.Y(n_12688)
);

NOR2x1_ASAP7_75t_SL g12689 ( 
.A(n_12264),
.B(n_12554),
.Y(n_12689)
);

NAND3xp33_ASAP7_75t_L g12690 ( 
.A(n_12562),
.B(n_1606),
.C(n_1608),
.Y(n_12690)
);

OAI21xp5_ASAP7_75t_L g12691 ( 
.A1(n_12514),
.A2(n_1608),
.B(n_1609),
.Y(n_12691)
);

INVx2_ASAP7_75t_SL g12692 ( 
.A(n_12330),
.Y(n_12692)
);

NOR2x1_ASAP7_75t_SL g12693 ( 
.A(n_12554),
.B(n_1608),
.Y(n_12693)
);

AOI22xp5_ASAP7_75t_L g12694 ( 
.A1(n_12485),
.A2(n_1611),
.B1(n_1609),
.B2(n_1610),
.Y(n_12694)
);

INVx3_ASAP7_75t_L g12695 ( 
.A(n_12321),
.Y(n_12695)
);

AND2x4_ASAP7_75t_L g12696 ( 
.A(n_12235),
.B(n_1609),
.Y(n_12696)
);

AND2x2_ASAP7_75t_L g12697 ( 
.A(n_12315),
.B(n_12338),
.Y(n_12697)
);

O2A1O1Ixp5_ASAP7_75t_L g12698 ( 
.A1(n_12565),
.A2(n_1612),
.B(n_1610),
.C(n_1611),
.Y(n_12698)
);

AO32x2_ASAP7_75t_L g12699 ( 
.A1(n_12570),
.A2(n_1612),
.A3(n_1610),
.B1(n_1611),
.B2(n_1613),
.Y(n_12699)
);

NOR2xp33_ASAP7_75t_SL g12700 ( 
.A(n_12490),
.B(n_12370),
.Y(n_12700)
);

OA21x2_ASAP7_75t_L g12701 ( 
.A1(n_12277),
.A2(n_1612),
.B(n_1613),
.Y(n_12701)
);

NAND4xp25_ASAP7_75t_L g12702 ( 
.A(n_12377),
.B(n_1615),
.C(n_1613),
.D(n_1614),
.Y(n_12702)
);

OAI22xp5_ASAP7_75t_L g12703 ( 
.A1(n_12513),
.A2(n_12533),
.B1(n_12500),
.B2(n_12496),
.Y(n_12703)
);

AND2x2_ASAP7_75t_L g12704 ( 
.A(n_12234),
.B(n_1614),
.Y(n_12704)
);

AND2x2_ASAP7_75t_L g12705 ( 
.A(n_12621),
.B(n_1614),
.Y(n_12705)
);

AOI211xp5_ASAP7_75t_L g12706 ( 
.A1(n_12399),
.A2(n_1617),
.B(n_1615),
.C(n_1616),
.Y(n_12706)
);

OAI211xp5_ASAP7_75t_L g12707 ( 
.A1(n_12619),
.A2(n_1618),
.B(n_1616),
.C(n_1617),
.Y(n_12707)
);

AND2x2_ASAP7_75t_L g12708 ( 
.A(n_12628),
.B(n_1616),
.Y(n_12708)
);

NOR2x1_ASAP7_75t_SL g12709 ( 
.A(n_12612),
.B(n_1617),
.Y(n_12709)
);

AND2x2_ASAP7_75t_L g12710 ( 
.A(n_12634),
.B(n_1618),
.Y(n_12710)
);

OA21x2_ASAP7_75t_L g12711 ( 
.A1(n_12352),
.A2(n_1618),
.B(n_1619),
.Y(n_12711)
);

AND2x4_ASAP7_75t_L g12712 ( 
.A(n_12455),
.B(n_1619),
.Y(n_12712)
);

INVx1_ASAP7_75t_L g12713 ( 
.A(n_12469),
.Y(n_12713)
);

OAI211xp5_ASAP7_75t_L g12714 ( 
.A1(n_12418),
.A2(n_1621),
.B(n_1619),
.C(n_1620),
.Y(n_12714)
);

NOR2x1_ASAP7_75t_SL g12715 ( 
.A(n_12441),
.B(n_1620),
.Y(n_12715)
);

AND2x2_ASAP7_75t_L g12716 ( 
.A(n_12642),
.B(n_1621),
.Y(n_12716)
);

AND2x2_ASAP7_75t_L g12717 ( 
.A(n_12646),
.B(n_1622),
.Y(n_12717)
);

INVx1_ASAP7_75t_L g12718 ( 
.A(n_12327),
.Y(n_12718)
);

OA21x2_ASAP7_75t_L g12719 ( 
.A1(n_12383),
.A2(n_1622),
.B(n_1623),
.Y(n_12719)
);

INVx3_ASAP7_75t_L g12720 ( 
.A(n_12321),
.Y(n_12720)
);

NOR2xp33_ASAP7_75t_L g12721 ( 
.A(n_12636),
.B(n_1622),
.Y(n_12721)
);

NAND3xp33_ASAP7_75t_L g12722 ( 
.A(n_12266),
.B(n_1623),
.C(n_1624),
.Y(n_12722)
);

BUFx3_ASAP7_75t_L g12723 ( 
.A(n_12422),
.Y(n_12723)
);

INVxp67_ASAP7_75t_L g12724 ( 
.A(n_12265),
.Y(n_12724)
);

AO21x2_ASAP7_75t_L g12725 ( 
.A1(n_12292),
.A2(n_1624),
.B(n_1625),
.Y(n_12725)
);

O2A1O1Ixp33_ASAP7_75t_L g12726 ( 
.A1(n_12648),
.A2(n_12364),
.B(n_12332),
.C(n_12541),
.Y(n_12726)
);

A2O1A1Ixp33_ASAP7_75t_L g12727 ( 
.A1(n_12556),
.A2(n_12548),
.B(n_12587),
.C(n_12520),
.Y(n_12727)
);

AND2x4_ASAP7_75t_L g12728 ( 
.A(n_12336),
.B(n_1625),
.Y(n_12728)
);

O2A1O1Ixp33_ASAP7_75t_SL g12729 ( 
.A1(n_12597),
.A2(n_1628),
.B(n_1626),
.C(n_1627),
.Y(n_12729)
);

AND2x2_ASAP7_75t_L g12730 ( 
.A(n_12652),
.B(n_1627),
.Y(n_12730)
);

NOR2xp33_ASAP7_75t_L g12731 ( 
.A(n_12408),
.B(n_12276),
.Y(n_12731)
);

OR2x2_ASAP7_75t_L g12732 ( 
.A(n_12274),
.B(n_1627),
.Y(n_12732)
);

OAI211xp5_ASAP7_75t_SL g12733 ( 
.A1(n_12609),
.A2(n_1636),
.B(n_1645),
.C(n_1628),
.Y(n_12733)
);

O2A1O1Ixp5_ASAP7_75t_L g12734 ( 
.A1(n_12367),
.A2(n_1630),
.B(n_1628),
.C(n_1629),
.Y(n_12734)
);

AO32x2_ASAP7_75t_L g12735 ( 
.A1(n_12449),
.A2(n_12535),
.A3(n_12357),
.B1(n_12280),
.B2(n_12437),
.Y(n_12735)
);

AND2x2_ASAP7_75t_L g12736 ( 
.A(n_12230),
.B(n_1629),
.Y(n_12736)
);

A2O1A1Ixp33_ASAP7_75t_L g12737 ( 
.A1(n_12559),
.A2(n_1632),
.B(n_1633),
.C(n_1631),
.Y(n_12737)
);

INVx2_ASAP7_75t_L g12738 ( 
.A(n_12410),
.Y(n_12738)
);

OR2x2_ASAP7_75t_L g12739 ( 
.A(n_12639),
.B(n_1630),
.Y(n_12739)
);

AOI22xp5_ASAP7_75t_L g12740 ( 
.A1(n_12348),
.A2(n_1634),
.B1(n_1632),
.B2(n_1633),
.Y(n_12740)
);

AOI221xp5_ASAP7_75t_L g12741 ( 
.A1(n_12301),
.A2(n_1635),
.B1(n_1632),
.B2(n_1634),
.C(n_1636),
.Y(n_12741)
);

AO32x2_ASAP7_75t_L g12742 ( 
.A1(n_12458),
.A2(n_1636),
.A3(n_1634),
.B1(n_1635),
.B2(n_1637),
.Y(n_12742)
);

AND2x2_ASAP7_75t_L g12743 ( 
.A(n_12242),
.B(n_1635),
.Y(n_12743)
);

AND2x2_ASAP7_75t_L g12744 ( 
.A(n_12629),
.B(n_12354),
.Y(n_12744)
);

OAI21xp5_ASAP7_75t_L g12745 ( 
.A1(n_12486),
.A2(n_12426),
.B(n_12419),
.Y(n_12745)
);

OAI21xp5_ASAP7_75t_L g12746 ( 
.A1(n_12381),
.A2(n_1638),
.B(n_1639),
.Y(n_12746)
);

OAI211xp5_ASAP7_75t_L g12747 ( 
.A1(n_12395),
.A2(n_1640),
.B(n_1638),
.C(n_1639),
.Y(n_12747)
);

OAI22xp5_ASAP7_75t_L g12748 ( 
.A1(n_12536),
.A2(n_1640),
.B1(n_1638),
.B2(n_1639),
.Y(n_12748)
);

AND2x2_ASAP7_75t_SL g12749 ( 
.A(n_12551),
.B(n_1640),
.Y(n_12749)
);

AND2x2_ASAP7_75t_L g12750 ( 
.A(n_12243),
.B(n_1641),
.Y(n_12750)
);

OA21x2_ASAP7_75t_L g12751 ( 
.A1(n_12281),
.A2(n_1641),
.B(n_1642),
.Y(n_12751)
);

AND2x2_ASAP7_75t_L g12752 ( 
.A(n_12622),
.B(n_1641),
.Y(n_12752)
);

INVx1_ASAP7_75t_L g12753 ( 
.A(n_12355),
.Y(n_12753)
);

NAND3xp33_ASAP7_75t_L g12754 ( 
.A(n_12345),
.B(n_1642),
.C(n_1643),
.Y(n_12754)
);

INVx5_ASAP7_75t_L g12755 ( 
.A(n_12302),
.Y(n_12755)
);

NAND2xp5_ASAP7_75t_L g12756 ( 
.A(n_12341),
.B(n_12460),
.Y(n_12756)
);

NAND2xp5_ASAP7_75t_L g12757 ( 
.A(n_12610),
.B(n_12245),
.Y(n_12757)
);

INVx2_ASAP7_75t_L g12758 ( 
.A(n_12410),
.Y(n_12758)
);

OAI22xp5_ASAP7_75t_SL g12759 ( 
.A1(n_12580),
.A2(n_1646),
.B1(n_1643),
.B2(n_1645),
.Y(n_12759)
);

OR2x2_ASAP7_75t_L g12760 ( 
.A(n_12297),
.B(n_1643),
.Y(n_12760)
);

OAI21xp5_ASAP7_75t_L g12761 ( 
.A1(n_12571),
.A2(n_1646),
.B(n_1647),
.Y(n_12761)
);

INVx2_ASAP7_75t_L g12762 ( 
.A(n_12433),
.Y(n_12762)
);

HB1xp67_ASAP7_75t_L g12763 ( 
.A(n_12396),
.Y(n_12763)
);

AND2x2_ASAP7_75t_L g12764 ( 
.A(n_12643),
.B(n_1646),
.Y(n_12764)
);

OAI21xp5_ASAP7_75t_L g12765 ( 
.A1(n_12558),
.A2(n_1647),
.B(n_1648),
.Y(n_12765)
);

HB1xp67_ASAP7_75t_L g12766 ( 
.A(n_12402),
.Y(n_12766)
);

AND2x2_ASAP7_75t_L g12767 ( 
.A(n_12651),
.B(n_1648),
.Y(n_12767)
);

A2O1A1Ixp33_ASAP7_75t_L g12768 ( 
.A1(n_12544),
.A2(n_1651),
.B(n_1652),
.C(n_1650),
.Y(n_12768)
);

NOR2x1_ASAP7_75t_SL g12769 ( 
.A(n_12373),
.B(n_1649),
.Y(n_12769)
);

AND2x2_ASAP7_75t_L g12770 ( 
.A(n_12304),
.B(n_1649),
.Y(n_12770)
);

A2O1A1Ixp33_ASAP7_75t_L g12771 ( 
.A1(n_12528),
.A2(n_1652),
.B(n_1653),
.C(n_1650),
.Y(n_12771)
);

AND2x2_ASAP7_75t_L g12772 ( 
.A(n_12339),
.B(n_1649),
.Y(n_12772)
);

OR2x2_ASAP7_75t_L g12773 ( 
.A(n_12476),
.B(n_1650),
.Y(n_12773)
);

AND2x2_ASAP7_75t_L g12774 ( 
.A(n_12465),
.B(n_1652),
.Y(n_12774)
);

OAI22xp5_ASAP7_75t_L g12775 ( 
.A1(n_12531),
.A2(n_1655),
.B1(n_1653),
.B2(n_1654),
.Y(n_12775)
);

INVx1_ASAP7_75t_L g12776 ( 
.A(n_12376),
.Y(n_12776)
);

AND2x2_ASAP7_75t_L g12777 ( 
.A(n_12445),
.B(n_1653),
.Y(n_12777)
);

INVx1_ASAP7_75t_L g12778 ( 
.A(n_12475),
.Y(n_12778)
);

INVx2_ASAP7_75t_L g12779 ( 
.A(n_12433),
.Y(n_12779)
);

NAND2xp33_ASAP7_75t_L g12780 ( 
.A(n_12605),
.B(n_1654),
.Y(n_12780)
);

AO32x2_ASAP7_75t_L g12781 ( 
.A1(n_12439),
.A2(n_1656),
.A3(n_1654),
.B1(n_1655),
.B2(n_1657),
.Y(n_12781)
);

INVx1_ASAP7_75t_L g12782 ( 
.A(n_12344),
.Y(n_12782)
);

NOR2xp33_ASAP7_75t_L g12783 ( 
.A(n_12575),
.B(n_12529),
.Y(n_12783)
);

AO32x2_ASAP7_75t_L g12784 ( 
.A1(n_12439),
.A2(n_1657),
.A3(n_1655),
.B1(n_1656),
.B2(n_1658),
.Y(n_12784)
);

AOI22xp5_ASAP7_75t_L g12785 ( 
.A1(n_12350),
.A2(n_1659),
.B1(n_1657),
.B2(n_1658),
.Y(n_12785)
);

AND2x2_ASAP7_75t_L g12786 ( 
.A(n_12488),
.B(n_1658),
.Y(n_12786)
);

INVx1_ASAP7_75t_L g12787 ( 
.A(n_12346),
.Y(n_12787)
);

CKINVDCx20_ASAP7_75t_R g12788 ( 
.A(n_12635),
.Y(n_12788)
);

AND2x2_ASAP7_75t_L g12789 ( 
.A(n_12507),
.B(n_1659),
.Y(n_12789)
);

OR2x6_ASAP7_75t_L g12790 ( 
.A(n_12302),
.B(n_1659),
.Y(n_12790)
);

AOI22xp33_ASAP7_75t_L g12791 ( 
.A1(n_12567),
.A2(n_1662),
.B1(n_1660),
.B2(n_1661),
.Y(n_12791)
);

OR2x6_ASAP7_75t_L g12792 ( 
.A(n_12284),
.B(n_1660),
.Y(n_12792)
);

AOI221xp5_ASAP7_75t_L g12793 ( 
.A1(n_12287),
.A2(n_1662),
.B1(n_1660),
.B2(n_1661),
.C(n_1663),
.Y(n_12793)
);

A2O1A1Ixp33_ASAP7_75t_L g12794 ( 
.A1(n_12532),
.A2(n_12534),
.B(n_12596),
.C(n_12550),
.Y(n_12794)
);

NOR2xp33_ASAP7_75t_L g12795 ( 
.A(n_12529),
.B(n_1661),
.Y(n_12795)
);

INVx3_ASAP7_75t_L g12796 ( 
.A(n_12385),
.Y(n_12796)
);

INVx4_ASAP7_75t_SL g12797 ( 
.A(n_12232),
.Y(n_12797)
);

O2A1O1Ixp33_ASAP7_75t_SL g12798 ( 
.A1(n_12461),
.A2(n_1665),
.B(n_1662),
.C(n_1664),
.Y(n_12798)
);

OAI22xp5_ASAP7_75t_L g12799 ( 
.A1(n_12506),
.A2(n_1666),
.B1(n_1664),
.B2(n_1665),
.Y(n_12799)
);

OAI211xp5_ASAP7_75t_L g12800 ( 
.A1(n_12615),
.A2(n_1667),
.B(n_1665),
.C(n_1666),
.Y(n_12800)
);

NOR2x1_ASAP7_75t_SL g12801 ( 
.A(n_12373),
.B(n_1668),
.Y(n_12801)
);

NAND2xp5_ASAP7_75t_L g12802 ( 
.A(n_12638),
.B(n_1668),
.Y(n_12802)
);

AND2x2_ASAP7_75t_L g12803 ( 
.A(n_12261),
.B(n_1668),
.Y(n_12803)
);

AO21x2_ASAP7_75t_L g12804 ( 
.A1(n_12625),
.A2(n_1669),
.B(n_1670),
.Y(n_12804)
);

AND2x2_ASAP7_75t_L g12805 ( 
.A(n_12526),
.B(n_1669),
.Y(n_12805)
);

OA21x2_ASAP7_75t_L g12806 ( 
.A1(n_12334),
.A2(n_1669),
.B(n_1670),
.Y(n_12806)
);

OR2x2_ASAP7_75t_L g12807 ( 
.A(n_12393),
.B(n_1670),
.Y(n_12807)
);

AND2x2_ASAP7_75t_L g12808 ( 
.A(n_12527),
.B(n_1671),
.Y(n_12808)
);

INVx1_ASAP7_75t_L g12809 ( 
.A(n_12384),
.Y(n_12809)
);

INVx2_ASAP7_75t_SL g12810 ( 
.A(n_12359),
.Y(n_12810)
);

BUFx6f_ASAP7_75t_L g12811 ( 
.A(n_12519),
.Y(n_12811)
);

OR2x2_ASAP7_75t_L g12812 ( 
.A(n_12400),
.B(n_12403),
.Y(n_12812)
);

OR2x2_ASAP7_75t_L g12813 ( 
.A(n_12407),
.B(n_1671),
.Y(n_12813)
);

OR2x2_ASAP7_75t_L g12814 ( 
.A(n_12416),
.B(n_1672),
.Y(n_12814)
);

NOR2xp33_ASAP7_75t_L g12815 ( 
.A(n_12509),
.B(n_1672),
.Y(n_12815)
);

AND2x4_ASAP7_75t_L g12816 ( 
.A(n_12414),
.B(n_1672),
.Y(n_12816)
);

NOR2xp33_ASAP7_75t_L g12817 ( 
.A(n_12617),
.B(n_1673),
.Y(n_12817)
);

OAI21x1_ASAP7_75t_L g12818 ( 
.A1(n_12401),
.A2(n_1675),
.B(n_1674),
.Y(n_12818)
);

INVx1_ASAP7_75t_L g12819 ( 
.A(n_12273),
.Y(n_12819)
);

AND2x2_ASAP7_75t_L g12820 ( 
.A(n_12311),
.B(n_1673),
.Y(n_12820)
);

NOR4xp25_ASAP7_75t_SL g12821 ( 
.A(n_12250),
.B(n_1675),
.C(n_1673),
.D(n_1674),
.Y(n_12821)
);

INVx1_ASAP7_75t_L g12822 ( 
.A(n_12360),
.Y(n_12822)
);

AO21x2_ASAP7_75t_L g12823 ( 
.A1(n_12627),
.A2(n_1675),
.B(n_1676),
.Y(n_12823)
);

OR2x2_ASAP7_75t_L g12824 ( 
.A(n_12423),
.B(n_12428),
.Y(n_12824)
);

AO21x2_ASAP7_75t_L g12825 ( 
.A1(n_12630),
.A2(n_1676),
.B(n_1677),
.Y(n_12825)
);

AOI21xp5_ASAP7_75t_L g12826 ( 
.A1(n_12537),
.A2(n_1677),
.B(n_1678),
.Y(n_12826)
);

OR2x2_ASAP7_75t_L g12827 ( 
.A(n_12430),
.B(n_1677),
.Y(n_12827)
);

AOI21x1_ASAP7_75t_L g12828 ( 
.A1(n_12417),
.A2(n_2441),
.B(n_1678),
.Y(n_12828)
);

AOI221xp5_ASAP7_75t_L g12829 ( 
.A1(n_12358),
.A2(n_1680),
.B1(n_1678),
.B2(n_1679),
.C(n_1681),
.Y(n_12829)
);

AND2x4_ASAP7_75t_L g12830 ( 
.A(n_12421),
.B(n_1679),
.Y(n_12830)
);

AO32x1_ASAP7_75t_L g12831 ( 
.A1(n_12343),
.A2(n_1696),
.A3(n_1705),
.B1(n_1688),
.B2(n_1680),
.Y(n_12831)
);

O2A1O1Ixp33_ASAP7_75t_L g12832 ( 
.A1(n_12608),
.A2(n_1682),
.B(n_1680),
.C(n_1681),
.Y(n_12832)
);

AND2x2_ASAP7_75t_L g12833 ( 
.A(n_12427),
.B(n_1682),
.Y(n_12833)
);

AND2x2_ASAP7_75t_L g12834 ( 
.A(n_12429),
.B(n_1683),
.Y(n_12834)
);

OR2x2_ASAP7_75t_L g12835 ( 
.A(n_12431),
.B(n_1683),
.Y(n_12835)
);

A2O1A1Ixp33_ASAP7_75t_L g12836 ( 
.A1(n_12572),
.A2(n_1685),
.B(n_1686),
.C(n_1684),
.Y(n_12836)
);

O2A1O1Ixp33_ASAP7_75t_L g12837 ( 
.A1(n_12238),
.A2(n_1686),
.B(n_1683),
.C(n_1685),
.Y(n_12837)
);

OAI21x1_ASAP7_75t_L g12838 ( 
.A1(n_12298),
.A2(n_1688),
.B(n_1687),
.Y(n_12838)
);

OAI22xp5_ASAP7_75t_L g12839 ( 
.A1(n_12503),
.A2(n_1688),
.B1(n_1685),
.B2(n_1687),
.Y(n_12839)
);

NOR2xp33_ASAP7_75t_L g12840 ( 
.A(n_12613),
.B(n_1687),
.Y(n_12840)
);

AND2x2_ASAP7_75t_L g12841 ( 
.A(n_12279),
.B(n_1689),
.Y(n_12841)
);

AOI22xp33_ASAP7_75t_L g12842 ( 
.A1(n_12283),
.A2(n_12573),
.B1(n_12227),
.B2(n_12375),
.Y(n_12842)
);

NAND2xp5_ASAP7_75t_L g12843 ( 
.A(n_12653),
.B(n_12656),
.Y(n_12843)
);

OA21x2_ASAP7_75t_L g12844 ( 
.A1(n_12286),
.A2(n_1689),
.B(n_1690),
.Y(n_12844)
);

AND2x2_ASAP7_75t_L g12845 ( 
.A(n_12378),
.B(n_1690),
.Y(n_12845)
);

OAI21xp5_ASAP7_75t_L g12846 ( 
.A1(n_12288),
.A2(n_1690),
.B(n_1691),
.Y(n_12846)
);

INVx1_ASAP7_75t_L g12847 ( 
.A(n_12365),
.Y(n_12847)
);

INVx4_ASAP7_75t_L g12848 ( 
.A(n_12397),
.Y(n_12848)
);

NAND2xp5_ASAP7_75t_L g12849 ( 
.A(n_12549),
.B(n_1691),
.Y(n_12849)
);

OR2x6_ASAP7_75t_L g12850 ( 
.A(n_12263),
.B(n_1691),
.Y(n_12850)
);

OAI21x1_ASAP7_75t_SL g12851 ( 
.A1(n_12270),
.A2(n_12640),
.B(n_12333),
.Y(n_12851)
);

AND2x2_ASAP7_75t_L g12852 ( 
.A(n_12553),
.B(n_1692),
.Y(n_12852)
);

AND2x2_ASAP7_75t_L g12853 ( 
.A(n_12555),
.B(n_1692),
.Y(n_12853)
);

NAND2xp5_ASAP7_75t_SL g12854 ( 
.A(n_12523),
.B(n_1693),
.Y(n_12854)
);

AND2x2_ASAP7_75t_L g12855 ( 
.A(n_12524),
.B(n_1693),
.Y(n_12855)
);

NOR2x1_ASAP7_75t_L g12856 ( 
.A(n_12411),
.B(n_1693),
.Y(n_12856)
);

NOR2x1_ASAP7_75t_SL g12857 ( 
.A(n_12415),
.B(n_12495),
.Y(n_12857)
);

INVx3_ASAP7_75t_L g12858 ( 
.A(n_12351),
.Y(n_12858)
);

NAND4xp25_ASAP7_75t_L g12859 ( 
.A(n_12252),
.B(n_1696),
.C(n_1694),
.D(n_1695),
.Y(n_12859)
);

INVx2_ASAP7_75t_L g12860 ( 
.A(n_12382),
.Y(n_12860)
);

OA21x2_ASAP7_75t_L g12861 ( 
.A1(n_12309),
.A2(n_1694),
.B(n_1695),
.Y(n_12861)
);

HB1xp67_ASAP7_75t_L g12862 ( 
.A(n_12452),
.Y(n_12862)
);

OAI22xp5_ASAP7_75t_L g12863 ( 
.A1(n_12557),
.A2(n_12545),
.B1(n_12574),
.B2(n_12530),
.Y(n_12863)
);

AND2x4_ASAP7_75t_L g12864 ( 
.A(n_12324),
.B(n_1695),
.Y(n_12864)
);

AND2x4_ASAP7_75t_L g12865 ( 
.A(n_12306),
.B(n_1696),
.Y(n_12865)
);

OR2x6_ASAP7_75t_L g12866 ( 
.A(n_12299),
.B(n_12467),
.Y(n_12866)
);

OAI21xp5_ASAP7_75t_L g12867 ( 
.A1(n_12325),
.A2(n_1697),
.B(n_1698),
.Y(n_12867)
);

NAND2xp33_ASAP7_75t_L g12868 ( 
.A(n_12614),
.B(n_1697),
.Y(n_12868)
);

AO32x2_ASAP7_75t_L g12869 ( 
.A1(n_12303),
.A2(n_1700),
.A3(n_1697),
.B1(n_1698),
.B2(n_1701),
.Y(n_12869)
);

AO32x2_ASAP7_75t_L g12870 ( 
.A1(n_12322),
.A2(n_1702),
.A3(n_1700),
.B1(n_1701),
.B2(n_1703),
.Y(n_12870)
);

NAND2xp33_ASAP7_75t_L g12871 ( 
.A(n_12618),
.B(n_1700),
.Y(n_12871)
);

BUFx3_ASAP7_75t_L g12872 ( 
.A(n_12468),
.Y(n_12872)
);

NAND2xp5_ASAP7_75t_L g12873 ( 
.A(n_12425),
.B(n_1701),
.Y(n_12873)
);

A2O1A1Ixp33_ASAP7_75t_L g12874 ( 
.A1(n_12505),
.A2(n_1704),
.B(n_1705),
.C(n_1703),
.Y(n_12874)
);

OAI21xp5_ASAP7_75t_L g12875 ( 
.A1(n_12595),
.A2(n_1702),
.B(n_1704),
.Y(n_12875)
);

NOR2xp33_ASAP7_75t_L g12876 ( 
.A(n_12440),
.B(n_1702),
.Y(n_12876)
);

O2A1O1Ixp33_ASAP7_75t_L g12877 ( 
.A1(n_12547),
.A2(n_1706),
.B(n_1704),
.C(n_1705),
.Y(n_12877)
);

INVx1_ASAP7_75t_L g12878 ( 
.A(n_12368),
.Y(n_12878)
);

AO32x2_ASAP7_75t_L g12879 ( 
.A1(n_12369),
.A2(n_1708),
.A3(n_1706),
.B1(n_1707),
.B2(n_1709),
.Y(n_12879)
);

NAND4xp25_ASAP7_75t_L g12880 ( 
.A(n_12253),
.B(n_1708),
.C(n_1706),
.D(n_1707),
.Y(n_12880)
);

INVx1_ASAP7_75t_L g12881 ( 
.A(n_12386),
.Y(n_12881)
);

NOR2xp33_ASAP7_75t_L g12882 ( 
.A(n_12569),
.B(n_1708),
.Y(n_12882)
);

AND2x2_ASAP7_75t_L g12883 ( 
.A(n_12435),
.B(n_1709),
.Y(n_12883)
);

NAND2xp33_ASAP7_75t_L g12884 ( 
.A(n_12603),
.B(n_1709),
.Y(n_12884)
);

AOI211xp5_ASAP7_75t_L g12885 ( 
.A1(n_12592),
.A2(n_1712),
.B(n_1710),
.C(n_1711),
.Y(n_12885)
);

OR2x2_ASAP7_75t_L g12886 ( 
.A(n_12436),
.B(n_1710),
.Y(n_12886)
);

AND2x2_ASAP7_75t_L g12887 ( 
.A(n_12566),
.B(n_12481),
.Y(n_12887)
);

OA21x2_ASAP7_75t_L g12888 ( 
.A1(n_12267),
.A2(n_1710),
.B(n_1711),
.Y(n_12888)
);

OR2x6_ASAP7_75t_L g12889 ( 
.A(n_12307),
.B(n_1711),
.Y(n_12889)
);

AND2x2_ASAP7_75t_L g12890 ( 
.A(n_12482),
.B(n_12257),
.Y(n_12890)
);

AND2x2_ASAP7_75t_L g12891 ( 
.A(n_12262),
.B(n_1712),
.Y(n_12891)
);

OAI21xp5_ASAP7_75t_L g12892 ( 
.A1(n_12600),
.A2(n_1713),
.B(n_1714),
.Y(n_12892)
);

O2A1O1Ixp33_ASAP7_75t_L g12893 ( 
.A1(n_12517),
.A2(n_1715),
.B(n_1713),
.C(n_1714),
.Y(n_12893)
);

INVx1_ASAP7_75t_L g12894 ( 
.A(n_12387),
.Y(n_12894)
);

OAI21xp5_ASAP7_75t_L g12895 ( 
.A1(n_12586),
.A2(n_12598),
.B(n_12579),
.Y(n_12895)
);

INVx1_ASAP7_75t_L g12896 ( 
.A(n_12391),
.Y(n_12896)
);

AND2x2_ASAP7_75t_L g12897 ( 
.A(n_12515),
.B(n_12313),
.Y(n_12897)
);

AOI221xp5_ASAP7_75t_L g12898 ( 
.A1(n_12585),
.A2(n_1717),
.B1(n_1715),
.B2(n_1716),
.C(n_1718),
.Y(n_12898)
);

AND2x2_ASAP7_75t_L g12899 ( 
.A(n_12319),
.B(n_1715),
.Y(n_12899)
);

AND2x2_ASAP7_75t_L g12900 ( 
.A(n_12320),
.B(n_12337),
.Y(n_12900)
);

OAI21xp5_ASAP7_75t_L g12901 ( 
.A1(n_12518),
.A2(n_1716),
.B(n_1717),
.Y(n_12901)
);

INVx1_ASAP7_75t_L g12902 ( 
.A(n_12271),
.Y(n_12902)
);

A2O1A1Ixp33_ASAP7_75t_L g12903 ( 
.A1(n_12611),
.A2(n_1720),
.B(n_1721),
.C(n_1719),
.Y(n_12903)
);

OR2x2_ASAP7_75t_L g12904 ( 
.A(n_12477),
.B(n_1716),
.Y(n_12904)
);

AOI22xp33_ASAP7_75t_SL g12905 ( 
.A1(n_12471),
.A2(n_1721),
.B1(n_1719),
.B2(n_1720),
.Y(n_12905)
);

NAND2xp5_ASAP7_75t_L g12906 ( 
.A(n_12604),
.B(n_1720),
.Y(n_12906)
);

OA21x2_ASAP7_75t_L g12907 ( 
.A1(n_12291),
.A2(n_1721),
.B(n_1722),
.Y(n_12907)
);

OAI21xp5_ASAP7_75t_L g12908 ( 
.A1(n_12588),
.A2(n_1722),
.B(n_1723),
.Y(n_12908)
);

AO21x2_ASAP7_75t_L g12909 ( 
.A1(n_12240),
.A2(n_1723),
.B(n_1724),
.Y(n_12909)
);

HB1xp67_ASAP7_75t_L g12910 ( 
.A(n_12259),
.Y(n_12910)
);

NOR2x1_ASAP7_75t_SL g12911 ( 
.A(n_12616),
.B(n_1723),
.Y(n_12911)
);

OR2x2_ASAP7_75t_L g12912 ( 
.A(n_12478),
.B(n_1724),
.Y(n_12912)
);

NOR2xp33_ASAP7_75t_L g12913 ( 
.A(n_12406),
.B(n_12329),
.Y(n_12913)
);

OR2x2_ASAP7_75t_L g12914 ( 
.A(n_12451),
.B(n_1724),
.Y(n_12914)
);

BUFx3_ASAP7_75t_L g12915 ( 
.A(n_12473),
.Y(n_12915)
);

AO21x2_ASAP7_75t_L g12916 ( 
.A1(n_12255),
.A2(n_1725),
.B(n_1726),
.Y(n_12916)
);

AND2x2_ASAP7_75t_L g12917 ( 
.A(n_12353),
.B(n_12366),
.Y(n_12917)
);

AND2x2_ASAP7_75t_L g12918 ( 
.A(n_12371),
.B(n_1725),
.Y(n_12918)
);

AND2x2_ASAP7_75t_L g12919 ( 
.A(n_12388),
.B(n_1726),
.Y(n_12919)
);

OA21x2_ASAP7_75t_L g12920 ( 
.A1(n_12268),
.A2(n_1726),
.B(n_1727),
.Y(n_12920)
);

NAND3xp33_ASAP7_75t_L g12921 ( 
.A(n_12483),
.B(n_1727),
.C(n_1728),
.Y(n_12921)
);

OAI21xp5_ASAP7_75t_L g12922 ( 
.A1(n_12479),
.A2(n_1727),
.B(n_1728),
.Y(n_12922)
);

AND2x6_ASAP7_75t_L g12923 ( 
.A(n_12389),
.B(n_1729),
.Y(n_12923)
);

AND2x4_ASAP7_75t_L g12924 ( 
.A(n_12504),
.B(n_1728),
.Y(n_12924)
);

INVx1_ASAP7_75t_L g12925 ( 
.A(n_12272),
.Y(n_12925)
);

AND2x2_ASAP7_75t_L g12926 ( 
.A(n_12349),
.B(n_1729),
.Y(n_12926)
);

AO32x2_ASAP7_75t_L g12927 ( 
.A1(n_12227),
.A2(n_1731),
.A3(n_1729),
.B1(n_1730),
.B2(n_1732),
.Y(n_12927)
);

INVxp33_ASAP7_75t_L g12928 ( 
.A(n_12649),
.Y(n_12928)
);

AND2x2_ASAP7_75t_L g12929 ( 
.A(n_12590),
.B(n_1730),
.Y(n_12929)
);

OAI21xp5_ASAP7_75t_L g12930 ( 
.A1(n_12470),
.A2(n_1730),
.B(n_1731),
.Y(n_12930)
);

INVx1_ASAP7_75t_L g12931 ( 
.A(n_12269),
.Y(n_12931)
);

A2O1A1Ixp33_ASAP7_75t_L g12932 ( 
.A1(n_12607),
.A2(n_1733),
.B(n_1734),
.C(n_1732),
.Y(n_12932)
);

AO21x2_ASAP7_75t_L g12933 ( 
.A1(n_12228),
.A2(n_1731),
.B(n_1733),
.Y(n_12933)
);

O2A1O1Ixp33_ASAP7_75t_SL g12934 ( 
.A1(n_12560),
.A2(n_1736),
.B(n_1734),
.C(n_1735),
.Y(n_12934)
);

AND2x2_ASAP7_75t_L g12935 ( 
.A(n_12462),
.B(n_1734),
.Y(n_12935)
);

A2O1A1Ixp33_ASAP7_75t_L g12936 ( 
.A1(n_12568),
.A2(n_1737),
.B(n_1738),
.C(n_1736),
.Y(n_12936)
);

AND2x2_ASAP7_75t_L g12937 ( 
.A(n_12463),
.B(n_1735),
.Y(n_12937)
);

OAI221xp5_ASAP7_75t_L g12938 ( 
.A1(n_12508),
.A2(n_1737),
.B1(n_1735),
.B2(n_1736),
.C(n_1738),
.Y(n_12938)
);

AND2x4_ASAP7_75t_L g12939 ( 
.A(n_12510),
.B(n_1739),
.Y(n_12939)
);

AOI22xp33_ASAP7_75t_L g12940 ( 
.A1(n_12356),
.A2(n_1741),
.B1(n_1739),
.B2(n_1740),
.Y(n_12940)
);

NAND2xp5_ASAP7_75t_L g12941 ( 
.A(n_12581),
.B(n_1739),
.Y(n_12941)
);

INVx2_ASAP7_75t_L g12942 ( 
.A(n_12447),
.Y(n_12942)
);

NAND4xp25_ASAP7_75t_L g12943 ( 
.A(n_12229),
.B(n_1742),
.C(n_1740),
.D(n_1741),
.Y(n_12943)
);

AO32x2_ASAP7_75t_L g12944 ( 
.A1(n_12443),
.A2(n_1742),
.A3(n_1740),
.B1(n_1741),
.B2(n_1743),
.Y(n_12944)
);

AND2x2_ASAP7_75t_L g12945 ( 
.A(n_12577),
.B(n_1742),
.Y(n_12945)
);

INVx2_ASAP7_75t_L g12946 ( 
.A(n_12522),
.Y(n_12946)
);

AOI22xp5_ASAP7_75t_L g12947 ( 
.A1(n_12540),
.A2(n_1745),
.B1(n_1743),
.B2(n_1744),
.Y(n_12947)
);

AND2x2_ASAP7_75t_L g12948 ( 
.A(n_12582),
.B(n_12362),
.Y(n_12948)
);

NOR2x1_ASAP7_75t_SL g12949 ( 
.A(n_12442),
.B(n_1743),
.Y(n_12949)
);

OAI211xp5_ASAP7_75t_SL g12950 ( 
.A1(n_12654),
.A2(n_1752),
.B(n_1760),
.C(n_1744),
.Y(n_12950)
);

OAI21xp5_ASAP7_75t_L g12951 ( 
.A1(n_12561),
.A2(n_12583),
.B(n_12546),
.Y(n_12951)
);

INVx3_ASAP7_75t_L g12952 ( 
.A(n_12446),
.Y(n_12952)
);

O2A1O1Ixp33_ASAP7_75t_SL g12953 ( 
.A1(n_12491),
.A2(n_1746),
.B(n_1744),
.C(n_1745),
.Y(n_12953)
);

AND2x2_ASAP7_75t_L g12954 ( 
.A(n_12372),
.B(n_1745),
.Y(n_12954)
);

AND2x4_ASAP7_75t_L g12955 ( 
.A(n_12434),
.B(n_1746),
.Y(n_12955)
);

AND2x2_ASAP7_75t_L g12956 ( 
.A(n_12438),
.B(n_1747),
.Y(n_12956)
);

OR2x2_ASAP7_75t_L g12957 ( 
.A(n_12563),
.B(n_1747),
.Y(n_12957)
);

AND2x2_ASAP7_75t_L g12958 ( 
.A(n_12285),
.B(n_12289),
.Y(n_12958)
);

OAI22xp5_ASAP7_75t_SL g12959 ( 
.A1(n_12589),
.A2(n_1750),
.B1(n_1748),
.B2(n_1749),
.Y(n_12959)
);

OAI22xp5_ASAP7_75t_L g12960 ( 
.A1(n_12498),
.A2(n_1750),
.B1(n_1748),
.B2(n_1749),
.Y(n_12960)
);

A2O1A1Ixp33_ASAP7_75t_L g12961 ( 
.A1(n_12293),
.A2(n_1753),
.B(n_1754),
.C(n_1752),
.Y(n_12961)
);

AND2x2_ASAP7_75t_L g12962 ( 
.A(n_12290),
.B(n_1751),
.Y(n_12962)
);

OAI21xp5_ASAP7_75t_L g12963 ( 
.A1(n_12525),
.A2(n_1751),
.B(n_1752),
.Y(n_12963)
);

OAI21xp5_ASAP7_75t_L g12964 ( 
.A1(n_12576),
.A2(n_1753),
.B(n_1754),
.Y(n_12964)
);

O2A1O1Ixp33_ASAP7_75t_L g12965 ( 
.A1(n_12606),
.A2(n_1756),
.B(n_1753),
.C(n_1755),
.Y(n_12965)
);

AND2x2_ASAP7_75t_L g12966 ( 
.A(n_12294),
.B(n_1755),
.Y(n_12966)
);

AO32x2_ASAP7_75t_L g12967 ( 
.A1(n_12340),
.A2(n_1757),
.A3(n_1755),
.B1(n_1756),
.B2(n_1758),
.Y(n_12967)
);

O2A1O1Ixp33_ASAP7_75t_SL g12968 ( 
.A1(n_12497),
.A2(n_1759),
.B(n_1757),
.C(n_1758),
.Y(n_12968)
);

OAI22xp5_ASAP7_75t_L g12969 ( 
.A1(n_12448),
.A2(n_1759),
.B1(n_1757),
.B2(n_1758),
.Y(n_12969)
);

OAI211xp5_ASAP7_75t_L g12970 ( 
.A1(n_12237),
.A2(n_1762),
.B(n_1759),
.C(n_1761),
.Y(n_12970)
);

A2O1A1Ixp33_ASAP7_75t_L g12971 ( 
.A1(n_12584),
.A2(n_1763),
.B(n_1764),
.C(n_1762),
.Y(n_12971)
);

OA21x2_ASAP7_75t_L g12972 ( 
.A1(n_12392),
.A2(n_1761),
.B(n_1763),
.Y(n_12972)
);

OA21x2_ASAP7_75t_L g12973 ( 
.A1(n_12317),
.A2(n_1764),
.B(n_1765),
.Y(n_12973)
);

NOR2x1_ASAP7_75t_SL g12974 ( 
.A(n_12432),
.B(n_1765),
.Y(n_12974)
);

INVxp33_ASAP7_75t_L g12975 ( 
.A(n_12494),
.Y(n_12975)
);

NAND2xp5_ASAP7_75t_L g12976 ( 
.A(n_12390),
.B(n_1765),
.Y(n_12976)
);

OR2x6_ASAP7_75t_L g12977 ( 
.A(n_12457),
.B(n_1766),
.Y(n_12977)
);

AND2x2_ASAP7_75t_L g12978 ( 
.A(n_12295),
.B(n_1766),
.Y(n_12978)
);

INVx1_ASAP7_75t_SL g12979 ( 
.A(n_12511),
.Y(n_12979)
);

OR2x2_ASAP7_75t_L g12980 ( 
.A(n_12300),
.B(n_1766),
.Y(n_12980)
);

NAND2xp5_ASAP7_75t_L g12981 ( 
.A(n_12390),
.B(n_1767),
.Y(n_12981)
);

INVx4_ASAP7_75t_L g12982 ( 
.A(n_12361),
.Y(n_12982)
);

INVx2_ASAP7_75t_L g12983 ( 
.A(n_12593),
.Y(n_12983)
);

AND2x2_ASAP7_75t_L g12984 ( 
.A(n_12667),
.B(n_12296),
.Y(n_12984)
);

HB1xp67_ASAP7_75t_L g12985 ( 
.A(n_12811),
.Y(n_12985)
);

BUFx3_ASAP7_75t_L g12986 ( 
.A(n_12660),
.Y(n_12986)
);

BUFx2_ASAP7_75t_L g12987 ( 
.A(n_12797),
.Y(n_12987)
);

INVx1_ASAP7_75t_L g12988 ( 
.A(n_12831),
.Y(n_12988)
);

INVx3_ASAP7_75t_L g12989 ( 
.A(n_12872),
.Y(n_12989)
);

INVx3_ASAP7_75t_L g12990 ( 
.A(n_12848),
.Y(n_12990)
);

INVx2_ASAP7_75t_L g12991 ( 
.A(n_12755),
.Y(n_12991)
);

AND2x2_ASAP7_75t_L g12992 ( 
.A(n_12697),
.B(n_12623),
.Y(n_12992)
);

OR2x2_ASAP7_75t_L g12993 ( 
.A(n_12703),
.B(n_12420),
.Y(n_12993)
);

BUFx2_ASAP7_75t_L g12994 ( 
.A(n_12723),
.Y(n_12994)
);

INVx2_ASAP7_75t_L g12995 ( 
.A(n_12755),
.Y(n_12995)
);

AND2x2_ASAP7_75t_L g12996 ( 
.A(n_12665),
.B(n_12631),
.Y(n_12996)
);

INVx2_ASAP7_75t_L g12997 ( 
.A(n_12974),
.Y(n_12997)
);

HB1xp67_ASAP7_75t_L g12998 ( 
.A(n_12811),
.Y(n_12998)
);

AND2x2_ASAP7_75t_L g12999 ( 
.A(n_12692),
.B(n_12632),
.Y(n_12999)
);

HB1xp67_ASAP7_75t_L g13000 ( 
.A(n_12900),
.Y(n_13000)
);

BUFx3_ASAP7_75t_L g13001 ( 
.A(n_12915),
.Y(n_13001)
);

INVx3_ASAP7_75t_L g13002 ( 
.A(n_12686),
.Y(n_13002)
);

INVx1_ASAP7_75t_L g13003 ( 
.A(n_12831),
.Y(n_13003)
);

NOR2x1_ASAP7_75t_L g13004 ( 
.A(n_12906),
.B(n_12459),
.Y(n_13004)
);

AND2x2_ASAP7_75t_L g13005 ( 
.A(n_12695),
.B(n_12633),
.Y(n_13005)
);

INVx1_ASAP7_75t_L g13006 ( 
.A(n_12672),
.Y(n_13006)
);

NAND2xp5_ASAP7_75t_L g13007 ( 
.A(n_12917),
.B(n_12982),
.Y(n_13007)
);

INVx2_ASAP7_75t_SL g13008 ( 
.A(n_12661),
.Y(n_13008)
);

AND2x2_ASAP7_75t_L g13009 ( 
.A(n_12720),
.B(n_12709),
.Y(n_13009)
);

INVxp67_ASAP7_75t_L g13010 ( 
.A(n_12693),
.Y(n_13010)
);

AND2x4_ASAP7_75t_L g13011 ( 
.A(n_12810),
.B(n_12489),
.Y(n_13011)
);

INVx1_ASAP7_75t_L g13012 ( 
.A(n_12732),
.Y(n_13012)
);

INVx2_ASAP7_75t_L g13013 ( 
.A(n_12769),
.Y(n_13013)
);

HB1xp67_ASAP7_75t_L g13014 ( 
.A(n_12766),
.Y(n_13014)
);

BUFx6f_ASAP7_75t_L g13015 ( 
.A(n_12777),
.Y(n_13015)
);

HB1xp67_ASAP7_75t_L g13016 ( 
.A(n_12952),
.Y(n_13016)
);

AND2x2_ASAP7_75t_L g13017 ( 
.A(n_12796),
.B(n_12641),
.Y(n_13017)
);

AND2x2_ASAP7_75t_L g13018 ( 
.A(n_12670),
.B(n_12644),
.Y(n_13018)
);

AND2x2_ASAP7_75t_L g13019 ( 
.A(n_12744),
.B(n_12239),
.Y(n_13019)
);

INVx2_ASAP7_75t_L g13020 ( 
.A(n_12801),
.Y(n_13020)
);

INVx2_ASAP7_75t_L g13021 ( 
.A(n_12866),
.Y(n_13021)
);

HB1xp67_ASAP7_75t_L g13022 ( 
.A(n_12724),
.Y(n_13022)
);

OR2x2_ASAP7_75t_L g13023 ( 
.A(n_12713),
.B(n_12241),
.Y(n_13023)
);

AND2x2_ASAP7_75t_L g13024 ( 
.A(n_12658),
.B(n_12637),
.Y(n_13024)
);

AND2x2_ASAP7_75t_L g13025 ( 
.A(n_12700),
.B(n_12244),
.Y(n_13025)
);

INVx1_ASAP7_75t_L g13026 ( 
.A(n_12739),
.Y(n_13026)
);

HB1xp67_ASAP7_75t_L g13027 ( 
.A(n_12897),
.Y(n_13027)
);

NAND2xp5_ASAP7_75t_L g13028 ( 
.A(n_12715),
.B(n_12323),
.Y(n_13028)
);

INVx2_ASAP7_75t_L g13029 ( 
.A(n_12889),
.Y(n_13029)
);

INVx1_ASAP7_75t_L g13030 ( 
.A(n_12742),
.Y(n_13030)
);

HB1xp67_ASAP7_75t_L g13031 ( 
.A(n_12757),
.Y(n_13031)
);

AND2x2_ASAP7_75t_L g13032 ( 
.A(n_12891),
.B(n_12246),
.Y(n_13032)
);

INVx1_ASAP7_75t_L g13033 ( 
.A(n_12742),
.Y(n_13033)
);

HB1xp67_ASAP7_75t_L g13034 ( 
.A(n_12682),
.Y(n_13034)
);

INVx1_ASAP7_75t_L g13035 ( 
.A(n_12688),
.Y(n_13035)
);

INVx1_ASAP7_75t_L g13036 ( 
.A(n_12676),
.Y(n_13036)
);

INVx1_ASAP7_75t_L g13037 ( 
.A(n_12676),
.Y(n_13037)
);

BUFx2_ASAP7_75t_L g13038 ( 
.A(n_12735),
.Y(n_13038)
);

AND2x2_ASAP7_75t_L g13039 ( 
.A(n_12926),
.B(n_12247),
.Y(n_13039)
);

INVx3_ASAP7_75t_L g13040 ( 
.A(n_12712),
.Y(n_13040)
);

NAND2x1_ASAP7_75t_L g13041 ( 
.A(n_12858),
.B(n_12248),
.Y(n_13041)
);

AND2x2_ASAP7_75t_L g13042 ( 
.A(n_12783),
.B(n_12249),
.Y(n_13042)
);

HB1xp67_ASAP7_75t_L g13043 ( 
.A(n_12862),
.Y(n_13043)
);

AND2x4_ASAP7_75t_L g13044 ( 
.A(n_12675),
.B(n_12480),
.Y(n_13044)
);

INVxp67_ASAP7_75t_SL g13045 ( 
.A(n_12657),
.Y(n_13045)
);

INVx2_ASAP7_75t_L g13046 ( 
.A(n_12889),
.Y(n_13046)
);

INVx1_ASAP7_75t_L g13047 ( 
.A(n_12869),
.Y(n_13047)
);

BUFx6f_ASAP7_75t_L g13048 ( 
.A(n_12680),
.Y(n_13048)
);

BUFx3_ASAP7_75t_L g13049 ( 
.A(n_12923),
.Y(n_13049)
);

BUFx3_ASAP7_75t_L g13050 ( 
.A(n_12923),
.Y(n_13050)
);

INVx1_ASAP7_75t_L g13051 ( 
.A(n_12869),
.Y(n_13051)
);

AOI22xp33_ASAP7_75t_SL g13052 ( 
.A1(n_12857),
.A2(n_12305),
.B1(n_12308),
.B2(n_12512),
.Y(n_13052)
);

BUFx2_ASAP7_75t_L g13053 ( 
.A(n_12735),
.Y(n_13053)
);

INVx2_ASAP7_75t_L g13054 ( 
.A(n_12792),
.Y(n_13054)
);

INVx2_ASAP7_75t_L g13055 ( 
.A(n_12949),
.Y(n_13055)
);

OR2x2_ASAP7_75t_L g13056 ( 
.A(n_12756),
.B(n_12413),
.Y(n_13056)
);

AND2x2_ASAP7_75t_L g13057 ( 
.A(n_12677),
.B(n_12538),
.Y(n_13057)
);

AND2x2_ASAP7_75t_L g13058 ( 
.A(n_12679),
.B(n_12731),
.Y(n_13058)
);

AND2x2_ASAP7_75t_L g13059 ( 
.A(n_12890),
.B(n_12738),
.Y(n_13059)
);

INVx5_ASAP7_75t_SL g13060 ( 
.A(n_12790),
.Y(n_13060)
);

AND2x2_ASAP7_75t_L g13061 ( 
.A(n_12758),
.B(n_12542),
.Y(n_13061)
);

INVx2_ASAP7_75t_L g13062 ( 
.A(n_12850),
.Y(n_13062)
);

INVx2_ASAP7_75t_L g13063 ( 
.A(n_12689),
.Y(n_13063)
);

BUFx3_ASAP7_75t_L g13064 ( 
.A(n_12923),
.Y(n_13064)
);

INVx2_ASAP7_75t_L g13065 ( 
.A(n_12977),
.Y(n_13065)
);

NOR2xp33_ASAP7_75t_L g13066 ( 
.A(n_12928),
.B(n_12310),
.Y(n_13066)
);

INVx3_ASAP7_75t_L g13067 ( 
.A(n_12728),
.Y(n_13067)
);

NOR4xp25_ASAP7_75t_SL g13068 ( 
.A(n_12794),
.B(n_12601),
.C(n_12444),
.D(n_12342),
.Y(n_13068)
);

INVx1_ASAP7_75t_L g13069 ( 
.A(n_12944),
.Y(n_13069)
);

OR2x2_ASAP7_75t_L g13070 ( 
.A(n_12668),
.B(n_12578),
.Y(n_13070)
);

NAND2xp5_ASAP7_75t_L g13071 ( 
.A(n_12979),
.B(n_12805),
.Y(n_13071)
);

AOI222xp33_ASAP7_75t_L g13072 ( 
.A1(n_12975),
.A2(n_12594),
.B1(n_12326),
.B2(n_12409),
.C1(n_12412),
.C2(n_12404),
.Y(n_13072)
);

AND2x2_ASAP7_75t_L g13073 ( 
.A(n_12762),
.B(n_12543),
.Y(n_13073)
);

INVx2_ASAP7_75t_L g13074 ( 
.A(n_12911),
.Y(n_13074)
);

INVx1_ASAP7_75t_L g13075 ( 
.A(n_12944),
.Y(n_13075)
);

INVx3_ASAP7_75t_L g13076 ( 
.A(n_12696),
.Y(n_13076)
);

AND2x2_ASAP7_75t_L g13077 ( 
.A(n_12779),
.B(n_12564),
.Y(n_13077)
);

BUFx3_ASAP7_75t_L g13078 ( 
.A(n_12899),
.Y(n_13078)
);

INVx1_ASAP7_75t_L g13079 ( 
.A(n_12773),
.Y(n_13079)
);

INVx1_ASAP7_75t_L g13080 ( 
.A(n_12967),
.Y(n_13080)
);

INVx1_ASAP7_75t_L g13081 ( 
.A(n_12967),
.Y(n_13081)
);

AND2x2_ASAP7_75t_L g13082 ( 
.A(n_12662),
.B(n_12521),
.Y(n_13082)
);

NOR2xp33_ASAP7_75t_L g13083 ( 
.A(n_12659),
.B(n_12493),
.Y(n_13083)
);

INVx4_ASAP7_75t_L g13084 ( 
.A(n_12736),
.Y(n_13084)
);

INVx2_ASAP7_75t_SL g13085 ( 
.A(n_12750),
.Y(n_13085)
);

INVx1_ASAP7_75t_L g13086 ( 
.A(n_12976),
.Y(n_13086)
);

INVx2_ASAP7_75t_L g13087 ( 
.A(n_12749),
.Y(n_13087)
);

NAND3xp33_ASAP7_75t_L g13088 ( 
.A(n_12694),
.B(n_12331),
.C(n_12379),
.Y(n_13088)
);

INVx2_ASAP7_75t_SL g13089 ( 
.A(n_12752),
.Y(n_13089)
);

INVx3_ASAP7_75t_L g13090 ( 
.A(n_12683),
.Y(n_13090)
);

NAND2xp5_ASAP7_75t_L g13091 ( 
.A(n_12808),
.B(n_12318),
.Y(n_13091)
);

INVx1_ASAP7_75t_L g13092 ( 
.A(n_12981),
.Y(n_13092)
);

INVx3_ASAP7_75t_L g13093 ( 
.A(n_12774),
.Y(n_13093)
);

OR2x2_ASAP7_75t_L g13094 ( 
.A(n_12763),
.B(n_12328),
.Y(n_13094)
);

INVx3_ASAP7_75t_L g13095 ( 
.A(n_12786),
.Y(n_13095)
);

HB1xp67_ASAP7_75t_L g13096 ( 
.A(n_12910),
.Y(n_13096)
);

OR2x2_ASAP7_75t_L g13097 ( 
.A(n_12812),
.B(n_12454),
.Y(n_13097)
);

INVx2_ASAP7_75t_L g13098 ( 
.A(n_12924),
.Y(n_13098)
);

INVx1_ASAP7_75t_L g13099 ( 
.A(n_12760),
.Y(n_13099)
);

INVx3_ASAP7_75t_L g13100 ( 
.A(n_12789),
.Y(n_13100)
);

INVx2_ASAP7_75t_L g13101 ( 
.A(n_12939),
.Y(n_13101)
);

AND2x2_ASAP7_75t_L g13102 ( 
.A(n_12704),
.B(n_12499),
.Y(n_13102)
);

INVx2_ASAP7_75t_L g13103 ( 
.A(n_12927),
.Y(n_13103)
);

AND2x2_ASAP7_75t_L g13104 ( 
.A(n_12705),
.B(n_12602),
.Y(n_13104)
);

OR2x2_ASAP7_75t_L g13105 ( 
.A(n_12824),
.B(n_12398),
.Y(n_13105)
);

INVx1_ASAP7_75t_L g13106 ( 
.A(n_12941),
.Y(n_13106)
);

AND2x2_ASAP7_75t_L g13107 ( 
.A(n_12708),
.B(n_12620),
.Y(n_13107)
);

INVx8_ASAP7_75t_L g13108 ( 
.A(n_12743),
.Y(n_13108)
);

INVx1_ASAP7_75t_L g13109 ( 
.A(n_12904),
.Y(n_13109)
);

OR2x2_ASAP7_75t_L g13110 ( 
.A(n_12863),
.B(n_12474),
.Y(n_13110)
);

INVx1_ASAP7_75t_L g13111 ( 
.A(n_12912),
.Y(n_13111)
);

BUFx2_ASAP7_75t_L g13112 ( 
.A(n_12710),
.Y(n_13112)
);

AND2x4_ASAP7_75t_L g13113 ( 
.A(n_12716),
.B(n_12282),
.Y(n_13113)
);

INVx1_ASAP7_75t_L g13114 ( 
.A(n_12807),
.Y(n_13114)
);

NAND2xp5_ASAP7_75t_L g13115 ( 
.A(n_12841),
.B(n_12424),
.Y(n_13115)
);

INVx1_ASAP7_75t_L g13116 ( 
.A(n_12813),
.Y(n_13116)
);

CKINVDCx20_ASAP7_75t_R g13117 ( 
.A(n_12788),
.Y(n_13117)
);

OR2x2_ASAP7_75t_L g13118 ( 
.A(n_12663),
.B(n_12456),
.Y(n_13118)
);

BUFx6f_ASAP7_75t_L g13119 ( 
.A(n_12770),
.Y(n_13119)
);

BUFx6f_ASAP7_75t_L g13120 ( 
.A(n_12673),
.Y(n_13120)
);

HB1xp67_ASAP7_75t_L g13121 ( 
.A(n_12701),
.Y(n_13121)
);

BUFx3_ASAP7_75t_L g13122 ( 
.A(n_12918),
.Y(n_13122)
);

INVx1_ASAP7_75t_L g13123 ( 
.A(n_12814),
.Y(n_13123)
);

OR2x2_ASAP7_75t_L g13124 ( 
.A(n_12702),
.B(n_12466),
.Y(n_13124)
);

INVx1_ASAP7_75t_L g13125 ( 
.A(n_12827),
.Y(n_13125)
);

INVx1_ASAP7_75t_L g13126 ( 
.A(n_12835),
.Y(n_13126)
);

AOI22xp33_ASAP7_75t_L g13127 ( 
.A1(n_12895),
.A2(n_12251),
.B1(n_12450),
.B2(n_12233),
.Y(n_13127)
);

OR2x2_ASAP7_75t_L g13128 ( 
.A(n_12664),
.B(n_12624),
.Y(n_13128)
);

INVx2_ASAP7_75t_L g13129 ( 
.A(n_12927),
.Y(n_13129)
);

INVx1_ASAP7_75t_L g13130 ( 
.A(n_12886),
.Y(n_13130)
);

HB1xp67_ASAP7_75t_L g13131 ( 
.A(n_12711),
.Y(n_13131)
);

OR2x2_ASAP7_75t_L g13132 ( 
.A(n_12778),
.B(n_12650),
.Y(n_13132)
);

OAI22xp33_ASAP7_75t_L g13133 ( 
.A1(n_12843),
.A2(n_1769),
.B1(n_1767),
.B2(n_1768),
.Y(n_13133)
);

AND2x2_ASAP7_75t_L g13134 ( 
.A(n_12717),
.B(n_1767),
.Y(n_13134)
);

INVx1_ASAP7_75t_L g13135 ( 
.A(n_12914),
.Y(n_13135)
);

INVx2_ASAP7_75t_L g13136 ( 
.A(n_12955),
.Y(n_13136)
);

BUFx6f_ASAP7_75t_L g13137 ( 
.A(n_12919),
.Y(n_13137)
);

INVx2_ASAP7_75t_L g13138 ( 
.A(n_12816),
.Y(n_13138)
);

HB1xp67_ASAP7_75t_L g13139 ( 
.A(n_12983),
.Y(n_13139)
);

AND2x2_ASAP7_75t_L g13140 ( 
.A(n_12730),
.B(n_12962),
.Y(n_13140)
);

AND2x2_ASAP7_75t_L g13141 ( 
.A(n_12966),
.B(n_1768),
.Y(n_13141)
);

INVx2_ASAP7_75t_L g13142 ( 
.A(n_12830),
.Y(n_13142)
);

NAND2xp5_ASAP7_75t_L g13143 ( 
.A(n_12933),
.B(n_2432),
.Y(n_13143)
);

AND2x2_ASAP7_75t_L g13144 ( 
.A(n_12978),
.B(n_1769),
.Y(n_13144)
);

INVx2_ASAP7_75t_L g13145 ( 
.A(n_12806),
.Y(n_13145)
);

NAND2x1p5_ASAP7_75t_L g13146 ( 
.A(n_12681),
.B(n_1769),
.Y(n_13146)
);

NAND2xp5_ASAP7_75t_L g13147 ( 
.A(n_12856),
.B(n_2433),
.Y(n_13147)
);

INVx2_ASAP7_75t_SL g13148 ( 
.A(n_12764),
.Y(n_13148)
);

INVx1_ASAP7_75t_L g13149 ( 
.A(n_12873),
.Y(n_13149)
);

OAI21xp5_ASAP7_75t_L g13150 ( 
.A1(n_12666),
.A2(n_1770),
.B(n_1771),
.Y(n_13150)
);

NAND2xp5_ASAP7_75t_L g13151 ( 
.A(n_12883),
.B(n_2434),
.Y(n_13151)
);

AOI33xp33_ASAP7_75t_L g13152 ( 
.A1(n_12726),
.A2(n_1772),
.A3(n_1774),
.B1(n_1770),
.B2(n_1771),
.B3(n_1773),
.Y(n_13152)
);

AND2x2_ASAP7_75t_L g13153 ( 
.A(n_12958),
.B(n_1772),
.Y(n_13153)
);

OR2x2_ASAP7_75t_L g13154 ( 
.A(n_12819),
.B(n_1773),
.Y(n_13154)
);

HB1xp67_ASAP7_75t_L g13155 ( 
.A(n_12948),
.Y(n_13155)
);

INVx1_ASAP7_75t_L g13156 ( 
.A(n_12879),
.Y(n_13156)
);

AND2x4_ASAP7_75t_L g13157 ( 
.A(n_12767),
.B(n_1773),
.Y(n_13157)
);

AND2x2_ASAP7_75t_L g13158 ( 
.A(n_12954),
.B(n_1774),
.Y(n_13158)
);

HB1xp67_ASAP7_75t_L g13159 ( 
.A(n_12887),
.Y(n_13159)
);

INVx1_ASAP7_75t_L g13160 ( 
.A(n_12879),
.Y(n_13160)
);

INVx2_ASAP7_75t_SL g13161 ( 
.A(n_12803),
.Y(n_13161)
);

OR2x2_ASAP7_75t_L g13162 ( 
.A(n_12847),
.B(n_1774),
.Y(n_13162)
);

INVx1_ASAP7_75t_L g13163 ( 
.A(n_12870),
.Y(n_13163)
);

OR2x2_ASAP7_75t_L g13164 ( 
.A(n_12878),
.B(n_1775),
.Y(n_13164)
);

INVx1_ASAP7_75t_L g13165 ( 
.A(n_12870),
.Y(n_13165)
);

INVx2_ASAP7_75t_L g13166 ( 
.A(n_12844),
.Y(n_13166)
);

INVx1_ASAP7_75t_L g13167 ( 
.A(n_12935),
.Y(n_13167)
);

INVx3_ASAP7_75t_L g13168 ( 
.A(n_12864),
.Y(n_13168)
);

INVx1_ASAP7_75t_L g13169 ( 
.A(n_12937),
.Y(n_13169)
);

NAND2xp5_ASAP7_75t_L g13170 ( 
.A(n_12913),
.B(n_2442),
.Y(n_13170)
);

BUFx2_ASAP7_75t_L g13171 ( 
.A(n_12881),
.Y(n_13171)
);

OR2x2_ASAP7_75t_L g13172 ( 
.A(n_12894),
.B(n_1775),
.Y(n_13172)
);

AND2x2_ASAP7_75t_L g13173 ( 
.A(n_12896),
.B(n_1776),
.Y(n_13173)
);

INVx2_ASAP7_75t_L g13174 ( 
.A(n_12861),
.Y(n_13174)
);

OAI22xp5_ASAP7_75t_L g13175 ( 
.A1(n_12687),
.A2(n_12842),
.B1(n_12947),
.B2(n_12722),
.Y(n_13175)
);

AND2x2_ASAP7_75t_L g13176 ( 
.A(n_12671),
.B(n_1776),
.Y(n_13176)
);

INVx3_ASAP7_75t_L g13177 ( 
.A(n_12865),
.Y(n_13177)
);

INVx1_ASAP7_75t_L g13178 ( 
.A(n_12802),
.Y(n_13178)
);

INVx1_ASAP7_75t_L g13179 ( 
.A(n_12980),
.Y(n_13179)
);

INVx2_ASAP7_75t_L g13180 ( 
.A(n_12888),
.Y(n_13180)
);

AND2x2_ASAP7_75t_L g13181 ( 
.A(n_12721),
.B(n_1777),
.Y(n_13181)
);

INVx1_ASAP7_75t_L g13182 ( 
.A(n_12957),
.Y(n_13182)
);

AO21x2_ASAP7_75t_L g13183 ( 
.A1(n_12851),
.A2(n_1777),
.B(n_1778),
.Y(n_13183)
);

NAND2xp5_ASAP7_75t_L g13184 ( 
.A(n_12852),
.B(n_2445),
.Y(n_13184)
);

INVx1_ASAP7_75t_L g13185 ( 
.A(n_12956),
.Y(n_13185)
);

AND2x2_ASAP7_75t_L g13186 ( 
.A(n_12817),
.B(n_1777),
.Y(n_13186)
);

NAND2xp5_ASAP7_75t_L g13187 ( 
.A(n_12853),
.B(n_2447),
.Y(n_13187)
);

AND2x2_ASAP7_75t_L g13188 ( 
.A(n_12840),
.B(n_1779),
.Y(n_13188)
);

A2O1A1Ixp33_ASAP7_75t_L g13189 ( 
.A1(n_12727),
.A2(n_1781),
.B(n_1779),
.C(n_1780),
.Y(n_13189)
);

HB1xp67_ASAP7_75t_L g13190 ( 
.A(n_12929),
.Y(n_13190)
);

INVx2_ASAP7_75t_L g13191 ( 
.A(n_12907),
.Y(n_13191)
);

INVx1_ASAP7_75t_L g13192 ( 
.A(n_12849),
.Y(n_13192)
);

NOR2xp33_ASAP7_75t_L g13193 ( 
.A(n_12729),
.B(n_1780),
.Y(n_13193)
);

INVx1_ASAP7_75t_L g13194 ( 
.A(n_12699),
.Y(n_13194)
);

AND2x2_ASAP7_75t_L g13195 ( 
.A(n_12772),
.B(n_1781),
.Y(n_13195)
);

INVx2_ASAP7_75t_SL g13196 ( 
.A(n_12845),
.Y(n_13196)
);

BUFx6f_ASAP7_75t_L g13197 ( 
.A(n_12795),
.Y(n_13197)
);

OR2x2_ASAP7_75t_L g13198 ( 
.A(n_12859),
.B(n_1781),
.Y(n_13198)
);

AND2x2_ASAP7_75t_L g13199 ( 
.A(n_12855),
.B(n_1782),
.Y(n_13199)
);

INVx2_ASAP7_75t_L g13200 ( 
.A(n_12781),
.Y(n_13200)
);

AND2x4_ASAP7_75t_L g13201 ( 
.A(n_12820),
.B(n_1782),
.Y(n_13201)
);

BUFx2_ASAP7_75t_L g13202 ( 
.A(n_12781),
.Y(n_13202)
);

INVx4_ASAP7_75t_L g13203 ( 
.A(n_12833),
.Y(n_13203)
);

NAND2xp33_ASAP7_75t_R g13204 ( 
.A(n_12821),
.B(n_1782),
.Y(n_13204)
);

INVx1_ASAP7_75t_L g13205 ( 
.A(n_12699),
.Y(n_13205)
);

AND2x2_ASAP7_75t_L g13206 ( 
.A(n_12868),
.B(n_1783),
.Y(n_13206)
);

INVx2_ASAP7_75t_L g13207 ( 
.A(n_12784),
.Y(n_13207)
);

AND2x4_ASAP7_75t_L g13208 ( 
.A(n_12834),
.B(n_1783),
.Y(n_13208)
);

AND2x4_ASAP7_75t_SL g13209 ( 
.A(n_12860),
.B(n_12945),
.Y(n_13209)
);

OA21x2_ASAP7_75t_L g13210 ( 
.A1(n_12745),
.A2(n_1783),
.B(n_1784),
.Y(n_13210)
);

INVx2_ASAP7_75t_L g13211 ( 
.A(n_12784),
.Y(n_13211)
);

AND2x2_ASAP7_75t_L g13212 ( 
.A(n_12822),
.B(n_1784),
.Y(n_13212)
);

INVx1_ASAP7_75t_L g13213 ( 
.A(n_12719),
.Y(n_13213)
);

INVx2_ASAP7_75t_L g13214 ( 
.A(n_12909),
.Y(n_13214)
);

INVx2_ASAP7_75t_SL g13215 ( 
.A(n_12854),
.Y(n_13215)
);

HB1xp67_ASAP7_75t_L g13216 ( 
.A(n_12908),
.Y(n_13216)
);

NAND2xp5_ASAP7_75t_L g13217 ( 
.A(n_12706),
.B(n_2431),
.Y(n_13217)
);

AND2x4_ASAP7_75t_L g13218 ( 
.A(n_12765),
.B(n_1784),
.Y(n_13218)
);

AOI22xp33_ASAP7_75t_L g13219 ( 
.A1(n_12809),
.A2(n_1787),
.B1(n_1785),
.B2(n_1786),
.Y(n_13219)
);

HB1xp67_ASAP7_75t_L g13220 ( 
.A(n_12718),
.Y(n_13220)
);

BUFx2_ASAP7_75t_L g13221 ( 
.A(n_12963),
.Y(n_13221)
);

AND2x2_ASAP7_75t_L g13222 ( 
.A(n_12761),
.B(n_1785),
.Y(n_13222)
);

AOI22xp5_ASAP7_75t_SL g13223 ( 
.A1(n_13038),
.A2(n_12691),
.B1(n_12876),
.B2(n_12799),
.Y(n_13223)
);

NAND2xp5_ASAP7_75t_L g13224 ( 
.A(n_13057),
.B(n_13078),
.Y(n_13224)
);

OAI21xp5_ASAP7_75t_SL g13225 ( 
.A1(n_13053),
.A2(n_12733),
.B(n_12707),
.Y(n_13225)
);

NAND2xp5_ASAP7_75t_L g13226 ( 
.A(n_13122),
.B(n_13161),
.Y(n_13226)
);

NAND2xp5_ASAP7_75t_L g13227 ( 
.A(n_13140),
.B(n_12836),
.Y(n_13227)
);

NAND2xp5_ASAP7_75t_L g13228 ( 
.A(n_13112),
.B(n_13085),
.Y(n_13228)
);

NOR2xp33_ASAP7_75t_L g13229 ( 
.A(n_13117),
.B(n_12780),
.Y(n_13229)
);

NAND2xp5_ASAP7_75t_L g13230 ( 
.A(n_13089),
.B(n_12714),
.Y(n_13230)
);

NAND2xp5_ASAP7_75t_L g13231 ( 
.A(n_13148),
.B(n_12804),
.Y(n_13231)
);

OAI21xp33_ASAP7_75t_L g13232 ( 
.A1(n_13001),
.A2(n_12925),
.B(n_12902),
.Y(n_13232)
);

NOR3xp33_ASAP7_75t_L g13233 ( 
.A(n_12991),
.B(n_12759),
.C(n_12698),
.Y(n_13233)
);

NAND2xp5_ASAP7_75t_L g13234 ( 
.A(n_13137),
.B(n_12823),
.Y(n_13234)
);

NAND2xp5_ASAP7_75t_L g13235 ( 
.A(n_13137),
.B(n_12825),
.Y(n_13235)
);

NAND2xp5_ASAP7_75t_L g13236 ( 
.A(n_13153),
.B(n_13196),
.Y(n_13236)
);

NAND2xp5_ASAP7_75t_L g13237 ( 
.A(n_13006),
.B(n_12674),
.Y(n_13237)
);

OAI22xp5_ASAP7_75t_L g13238 ( 
.A1(n_13052),
.A2(n_12921),
.B1(n_12771),
.B2(n_12785),
.Y(n_13238)
);

NAND2xp5_ASAP7_75t_L g13239 ( 
.A(n_13076),
.B(n_12725),
.Y(n_13239)
);

OAI21xp33_ASAP7_75t_L g13240 ( 
.A1(n_13025),
.A2(n_12931),
.B(n_12776),
.Y(n_13240)
);

OAI22xp5_ASAP7_75t_L g13241 ( 
.A1(n_12993),
.A2(n_12690),
.B1(n_12791),
.B2(n_12905),
.Y(n_13241)
);

NAND2xp5_ASAP7_75t_SL g13242 ( 
.A(n_13015),
.B(n_12951),
.Y(n_13242)
);

AND2x2_ASAP7_75t_L g13243 ( 
.A(n_12987),
.B(n_12986),
.Y(n_13243)
);

OA21x2_ASAP7_75t_L g13244 ( 
.A1(n_12988),
.A2(n_12826),
.B(n_12901),
.Y(n_13244)
);

NOR3xp33_ASAP7_75t_L g13245 ( 
.A(n_12995),
.B(n_12800),
.C(n_12747),
.Y(n_13245)
);

AND2x2_ASAP7_75t_L g13246 ( 
.A(n_13009),
.B(n_12753),
.Y(n_13246)
);

AOI221xp5_ASAP7_75t_L g13247 ( 
.A1(n_13121),
.A2(n_12832),
.B1(n_12837),
.B2(n_12734),
.C(n_12934),
.Y(n_13247)
);

INVx1_ASAP7_75t_L g13248 ( 
.A(n_13096),
.Y(n_13248)
);

NAND2xp5_ASAP7_75t_L g13249 ( 
.A(n_13157),
.B(n_12882),
.Y(n_13249)
);

AND2x2_ASAP7_75t_L g13250 ( 
.A(n_12994),
.B(n_12782),
.Y(n_13250)
);

OAI21xp5_ASAP7_75t_SL g13251 ( 
.A1(n_13010),
.A2(n_12880),
.B(n_12943),
.Y(n_13251)
);

NAND3xp33_ASAP7_75t_L g13252 ( 
.A(n_13131),
.B(n_12685),
.C(n_12678),
.Y(n_13252)
);

AND2x2_ASAP7_75t_L g13253 ( 
.A(n_13000),
.B(n_12787),
.Y(n_13253)
);

NAND2xp5_ASAP7_75t_SL g13254 ( 
.A(n_13015),
.B(n_12740),
.Y(n_13254)
);

AOI22xp33_ASAP7_75t_L g13255 ( 
.A1(n_13202),
.A2(n_12754),
.B1(n_12871),
.B2(n_12751),
.Y(n_13255)
);

NAND3xp33_ASAP7_75t_L g13256 ( 
.A(n_13068),
.B(n_12885),
.C(n_12793),
.Y(n_13256)
);

INVx1_ASAP7_75t_L g13257 ( 
.A(n_13027),
.Y(n_13257)
);

OAI221xp5_ASAP7_75t_L g13258 ( 
.A1(n_13045),
.A2(n_12829),
.B1(n_12741),
.B2(n_12737),
.C(n_12970),
.Y(n_13258)
);

NAND2xp5_ASAP7_75t_L g13259 ( 
.A(n_13167),
.B(n_12884),
.Y(n_13259)
);

NAND3xp33_ASAP7_75t_L g13260 ( 
.A(n_13031),
.B(n_12684),
.C(n_12898),
.Y(n_13260)
);

NOR2xp33_ASAP7_75t_L g13261 ( 
.A(n_13002),
.B(n_12953),
.Y(n_13261)
);

AND2x2_ASAP7_75t_L g13262 ( 
.A(n_12989),
.B(n_12922),
.Y(n_13262)
);

AND2x2_ASAP7_75t_L g13263 ( 
.A(n_13058),
.B(n_12990),
.Y(n_13263)
);

AND2x2_ASAP7_75t_L g13264 ( 
.A(n_13032),
.B(n_12930),
.Y(n_13264)
);

NAND4xp25_ASAP7_75t_L g13265 ( 
.A(n_13007),
.B(n_12964),
.C(n_12815),
.D(n_12893),
.Y(n_13265)
);

AND2x2_ASAP7_75t_L g13266 ( 
.A(n_13039),
.B(n_12942),
.Y(n_13266)
);

NAND2xp5_ASAP7_75t_L g13267 ( 
.A(n_13169),
.B(n_12968),
.Y(n_13267)
);

NAND2xp5_ASAP7_75t_L g13268 ( 
.A(n_13155),
.B(n_13044),
.Y(n_13268)
);

NAND3xp33_ASAP7_75t_L g13269 ( 
.A(n_13152),
.B(n_12932),
.C(n_12903),
.Y(n_13269)
);

NAND2xp5_ASAP7_75t_L g13270 ( 
.A(n_13090),
.B(n_12936),
.Y(n_13270)
);

NOR2xp33_ASAP7_75t_L g13271 ( 
.A(n_13084),
.B(n_12959),
.Y(n_13271)
);

AOI22xp33_ASAP7_75t_L g13272 ( 
.A1(n_13200),
.A2(n_12973),
.B1(n_12972),
.B2(n_12946),
.Y(n_13272)
);

NAND2xp5_ASAP7_75t_L g13273 ( 
.A(n_13093),
.B(n_12874),
.Y(n_13273)
);

OAI22xp5_ASAP7_75t_L g13274 ( 
.A1(n_13063),
.A2(n_12961),
.B1(n_12940),
.B2(n_12768),
.Y(n_13274)
);

NAND3xp33_ASAP7_75t_L g13275 ( 
.A(n_13175),
.B(n_12950),
.C(n_12892),
.Y(n_13275)
);

NAND2xp33_ASAP7_75t_SL g13276 ( 
.A(n_13041),
.B(n_12916),
.Y(n_13276)
);

NAND2xp5_ASAP7_75t_SL g13277 ( 
.A(n_13048),
.B(n_12746),
.Y(n_13277)
);

OAI21xp5_ASAP7_75t_SL g13278 ( 
.A1(n_13003),
.A2(n_12877),
.B(n_12965),
.Y(n_13278)
);

NAND2xp5_ASAP7_75t_SL g13279 ( 
.A(n_13048),
.B(n_12828),
.Y(n_13279)
);

NAND2xp5_ASAP7_75t_L g13280 ( 
.A(n_13095),
.B(n_12920),
.Y(n_13280)
);

NAND2xp5_ASAP7_75t_L g13281 ( 
.A(n_13100),
.B(n_12875),
.Y(n_13281)
);

NAND2xp5_ASAP7_75t_L g13282 ( 
.A(n_13203),
.B(n_12971),
.Y(n_13282)
);

NAND2xp5_ASAP7_75t_L g13283 ( 
.A(n_13120),
.B(n_12846),
.Y(n_13283)
);

NAND2xp5_ASAP7_75t_L g13284 ( 
.A(n_13120),
.B(n_12839),
.Y(n_13284)
);

NAND3xp33_ASAP7_75t_L g13285 ( 
.A(n_13189),
.B(n_12867),
.C(n_12669),
.Y(n_13285)
);

AND2x2_ASAP7_75t_L g13286 ( 
.A(n_12985),
.B(n_12748),
.Y(n_13286)
);

NAND2xp33_ASAP7_75t_SL g13287 ( 
.A(n_13159),
.B(n_12775),
.Y(n_13287)
);

NAND2xp5_ASAP7_75t_L g13288 ( 
.A(n_13185),
.B(n_12798),
.Y(n_13288)
);

OAI21xp5_ASAP7_75t_SL g13289 ( 
.A1(n_12984),
.A2(n_12960),
.B(n_12938),
.Y(n_13289)
);

NAND2xp33_ASAP7_75t_SL g13290 ( 
.A(n_13008),
.B(n_12969),
.Y(n_13290)
);

NAND3xp33_ASAP7_75t_L g13291 ( 
.A(n_13216),
.B(n_12838),
.C(n_12818),
.Y(n_13291)
);

NOR2xp33_ASAP7_75t_L g13292 ( 
.A(n_12997),
.B(n_1787),
.Y(n_13292)
);

AND2x2_ASAP7_75t_L g13293 ( 
.A(n_12998),
.B(n_1787),
.Y(n_13293)
);

AOI22xp33_ASAP7_75t_L g13294 ( 
.A1(n_13207),
.A2(n_1790),
.B1(n_1788),
.B2(n_1789),
.Y(n_13294)
);

INVx2_ASAP7_75t_L g13295 ( 
.A(n_13146),
.Y(n_13295)
);

AND2x2_ASAP7_75t_L g13296 ( 
.A(n_13059),
.B(n_1788),
.Y(n_13296)
);

NAND3xp33_ASAP7_75t_L g13297 ( 
.A(n_13119),
.B(n_1790),
.C(n_1789),
.Y(n_13297)
);

NAND2xp5_ASAP7_75t_L g13298 ( 
.A(n_13099),
.B(n_13182),
.Y(n_13298)
);

OR2x2_ASAP7_75t_L g13299 ( 
.A(n_13071),
.B(n_1788),
.Y(n_13299)
);

AOI221x1_ASAP7_75t_SL g13300 ( 
.A1(n_13011),
.A2(n_1791),
.B1(n_1789),
.B2(n_1790),
.C(n_1792),
.Y(n_13300)
);

NAND3xp33_ASAP7_75t_L g13301 ( 
.A(n_13119),
.B(n_1793),
.C(n_1792),
.Y(n_13301)
);

NAND2xp5_ASAP7_75t_L g13302 ( 
.A(n_13193),
.B(n_1791),
.Y(n_13302)
);

NOR2xp33_ASAP7_75t_L g13303 ( 
.A(n_13040),
.B(n_1791),
.Y(n_13303)
);

NAND2xp5_ASAP7_75t_L g13304 ( 
.A(n_13026),
.B(n_1792),
.Y(n_13304)
);

NAND2xp5_ASAP7_75t_L g13305 ( 
.A(n_13012),
.B(n_1793),
.Y(n_13305)
);

OAI21xp5_ASAP7_75t_SL g13306 ( 
.A1(n_13013),
.A2(n_1794),
.B(n_1795),
.Y(n_13306)
);

NOR2xp33_ASAP7_75t_SL g13307 ( 
.A(n_13020),
.B(n_1794),
.Y(n_13307)
);

NAND2xp5_ASAP7_75t_SL g13308 ( 
.A(n_13055),
.B(n_1795),
.Y(n_13308)
);

AND2x2_ASAP7_75t_L g13309 ( 
.A(n_13034),
.B(n_1795),
.Y(n_13309)
);

AND2x2_ASAP7_75t_SL g13310 ( 
.A(n_13074),
.B(n_1796),
.Y(n_13310)
);

NAND3xp33_ASAP7_75t_L g13311 ( 
.A(n_13072),
.B(n_1798),
.C(n_1797),
.Y(n_13311)
);

NAND2xp5_ASAP7_75t_L g13312 ( 
.A(n_13060),
.B(n_1796),
.Y(n_13312)
);

NAND2xp5_ASAP7_75t_L g13313 ( 
.A(n_13215),
.B(n_1796),
.Y(n_13313)
);

OAI22xp33_ASAP7_75t_L g13314 ( 
.A1(n_13110),
.A2(n_1799),
.B1(n_1797),
.B2(n_1798),
.Y(n_13314)
);

AND2x2_ASAP7_75t_L g13315 ( 
.A(n_13016),
.B(n_1797),
.Y(n_13315)
);

NAND2xp5_ASAP7_75t_L g13316 ( 
.A(n_13212),
.B(n_1798),
.Y(n_13316)
);

OAI221xp5_ASAP7_75t_SL g13317 ( 
.A1(n_13056),
.A2(n_1801),
.B1(n_1799),
.B2(n_1800),
.C(n_1802),
.Y(n_13317)
);

AND2x2_ASAP7_75t_L g13318 ( 
.A(n_12992),
.B(n_1800),
.Y(n_13318)
);

OAI21xp5_ASAP7_75t_SL g13319 ( 
.A1(n_13022),
.A2(n_1801),
.B(n_1803),
.Y(n_13319)
);

AND2x2_ASAP7_75t_L g13320 ( 
.A(n_12999),
.B(n_1803),
.Y(n_13320)
);

HB1xp67_ASAP7_75t_L g13321 ( 
.A(n_13183),
.Y(n_13321)
);

OAI21xp5_ASAP7_75t_SL g13322 ( 
.A1(n_13024),
.A2(n_1803),
.B(n_1804),
.Y(n_13322)
);

NAND2xp5_ASAP7_75t_L g13323 ( 
.A(n_13035),
.B(n_1804),
.Y(n_13323)
);

OAI221xp5_ASAP7_75t_SL g13324 ( 
.A1(n_13094),
.A2(n_1806),
.B1(n_1804),
.B2(n_1805),
.C(n_1807),
.Y(n_13324)
);

INVx1_ASAP7_75t_L g13325 ( 
.A(n_13190),
.Y(n_13325)
);

NAND2xp5_ASAP7_75t_L g13326 ( 
.A(n_13079),
.B(n_1805),
.Y(n_13326)
);

AOI221xp5_ASAP7_75t_L g13327 ( 
.A1(n_13163),
.A2(n_1807),
.B1(n_1805),
.B2(n_1806),
.C(n_1808),
.Y(n_13327)
);

AOI21xp5_ASAP7_75t_SL g13328 ( 
.A1(n_13028),
.A2(n_1810),
.B(n_1809),
.Y(n_13328)
);

OAI221xp5_ASAP7_75t_SL g13329 ( 
.A1(n_13105),
.A2(n_1812),
.B1(n_1808),
.B2(n_1811),
.C(n_1813),
.Y(n_13329)
);

OAI21xp33_ASAP7_75t_L g13330 ( 
.A1(n_13021),
.A2(n_1808),
.B(n_1811),
.Y(n_13330)
);

OAI221xp5_ASAP7_75t_L g13331 ( 
.A1(n_13165),
.A2(n_1813),
.B1(n_1811),
.B2(n_1812),
.C(n_1815),
.Y(n_13331)
);

AND2x2_ASAP7_75t_L g13332 ( 
.A(n_13019),
.B(n_1815),
.Y(n_13332)
);

AND2x2_ASAP7_75t_L g13333 ( 
.A(n_13017),
.B(n_1815),
.Y(n_13333)
);

OAI21xp5_ASAP7_75t_L g13334 ( 
.A1(n_13004),
.A2(n_13088),
.B(n_13083),
.Y(n_13334)
);

NAND2xp5_ASAP7_75t_SL g13335 ( 
.A(n_13067),
.B(n_1816),
.Y(n_13335)
);

AOI211xp5_ASAP7_75t_L g13336 ( 
.A1(n_13066),
.A2(n_1824),
.B(n_1832),
.C(n_1816),
.Y(n_13336)
);

NAND2xp5_ASAP7_75t_L g13337 ( 
.A(n_13173),
.B(n_1817),
.Y(n_13337)
);

NOR2xp33_ASAP7_75t_R g13338 ( 
.A(n_13204),
.B(n_2432),
.Y(n_13338)
);

OAI22xp5_ASAP7_75t_L g13339 ( 
.A1(n_13070),
.A2(n_1820),
.B1(n_1818),
.B2(n_1819),
.Y(n_13339)
);

NOR3xp33_ASAP7_75t_L g13340 ( 
.A(n_13086),
.B(n_1818),
.C(n_1819),
.Y(n_13340)
);

OAI211xp5_ASAP7_75t_L g13341 ( 
.A1(n_13043),
.A2(n_1820),
.B(n_1818),
.C(n_1819),
.Y(n_13341)
);

NAND2xp5_ASAP7_75t_L g13342 ( 
.A(n_13109),
.B(n_1820),
.Y(n_13342)
);

NAND3xp33_ASAP7_75t_L g13343 ( 
.A(n_13139),
.B(n_13014),
.C(n_13197),
.Y(n_13343)
);

OAI21xp33_ASAP7_75t_L g13344 ( 
.A1(n_13042),
.A2(n_1821),
.B(n_1822),
.Y(n_13344)
);

NAND3xp33_ASAP7_75t_L g13345 ( 
.A(n_13197),
.B(n_1823),
.C(n_1822),
.Y(n_13345)
);

NOR3xp33_ASAP7_75t_SL g13346 ( 
.A(n_13149),
.B(n_1821),
.C(n_1822),
.Y(n_13346)
);

OAI221xp5_ASAP7_75t_SL g13347 ( 
.A1(n_13036),
.A2(n_1825),
.B1(n_1823),
.B2(n_1824),
.C(n_1826),
.Y(n_13347)
);

NOR3xp33_ASAP7_75t_L g13348 ( 
.A(n_13092),
.B(n_1823),
.C(n_1825),
.Y(n_13348)
);

NAND2xp5_ASAP7_75t_SL g13349 ( 
.A(n_12996),
.B(n_1825),
.Y(n_13349)
);

AND2x2_ASAP7_75t_L g13350 ( 
.A(n_13018),
.B(n_1826),
.Y(n_13350)
);

OAI21xp5_ASAP7_75t_L g13351 ( 
.A1(n_13133),
.A2(n_13217),
.B(n_13150),
.Y(n_13351)
);

AND2x2_ASAP7_75t_L g13352 ( 
.A(n_13005),
.B(n_1827),
.Y(n_13352)
);

OAI21xp5_ASAP7_75t_SL g13353 ( 
.A1(n_13171),
.A2(n_1827),
.B(n_1828),
.Y(n_13353)
);

NAND2xp5_ASAP7_75t_L g13354 ( 
.A(n_13111),
.B(n_1827),
.Y(n_13354)
);

NAND2xp5_ASAP7_75t_L g13355 ( 
.A(n_13114),
.B(n_1828),
.Y(n_13355)
);

NAND4xp25_ASAP7_75t_L g13356 ( 
.A(n_13023),
.B(n_1830),
.C(n_1828),
.D(n_1829),
.Y(n_13356)
);

NAND2xp5_ASAP7_75t_L g13357 ( 
.A(n_13116),
.B(n_1829),
.Y(n_13357)
);

OAI21xp5_ASAP7_75t_SL g13358 ( 
.A1(n_13061),
.A2(n_1829),
.B(n_1830),
.Y(n_13358)
);

AND2x2_ASAP7_75t_L g13359 ( 
.A(n_13073),
.B(n_1830),
.Y(n_13359)
);

OAI22xp5_ASAP7_75t_L g13360 ( 
.A1(n_13124),
.A2(n_1833),
.B1(n_1831),
.B2(n_1832),
.Y(n_13360)
);

NAND2xp5_ASAP7_75t_L g13361 ( 
.A(n_13123),
.B(n_1831),
.Y(n_13361)
);

AOI22xp33_ASAP7_75t_L g13362 ( 
.A1(n_13211),
.A2(n_1834),
.B1(n_1832),
.B2(n_1833),
.Y(n_13362)
);

AND2x2_ASAP7_75t_L g13363 ( 
.A(n_13077),
.B(n_1833),
.Y(n_13363)
);

AND2x2_ASAP7_75t_L g13364 ( 
.A(n_13104),
.B(n_1835),
.Y(n_13364)
);

NAND3xp33_ASAP7_75t_L g13365 ( 
.A(n_13037),
.B(n_1837),
.C(n_1836),
.Y(n_13365)
);

AND2x2_ASAP7_75t_L g13366 ( 
.A(n_13107),
.B(n_1835),
.Y(n_13366)
);

NAND2xp5_ASAP7_75t_L g13367 ( 
.A(n_13125),
.B(n_1835),
.Y(n_13367)
);

AOI21xp5_ASAP7_75t_SL g13368 ( 
.A1(n_13154),
.A2(n_1838),
.B(n_1837),
.Y(n_13368)
);

AND2x2_ASAP7_75t_L g13369 ( 
.A(n_13220),
.B(n_1836),
.Y(n_13369)
);

OAI22xp5_ASAP7_75t_L g13370 ( 
.A1(n_13108),
.A2(n_13198),
.B1(n_13221),
.B2(n_13097),
.Y(n_13370)
);

NAND2xp5_ASAP7_75t_L g13371 ( 
.A(n_13126),
.B(n_1836),
.Y(n_13371)
);

NAND2xp5_ASAP7_75t_L g13372 ( 
.A(n_13130),
.B(n_1837),
.Y(n_13372)
);

OA211x2_ASAP7_75t_L g13373 ( 
.A1(n_13091),
.A2(n_1840),
.B(n_1838),
.C(n_1839),
.Y(n_13373)
);

NAND2xp5_ASAP7_75t_L g13374 ( 
.A(n_13135),
.B(n_1838),
.Y(n_13374)
);

NAND2xp5_ASAP7_75t_L g13375 ( 
.A(n_13179),
.B(n_1839),
.Y(n_13375)
);

NAND2xp5_ASAP7_75t_L g13376 ( 
.A(n_13218),
.B(n_1839),
.Y(n_13376)
);

NAND2xp5_ASAP7_75t_SL g13377 ( 
.A(n_13082),
.B(n_1840),
.Y(n_13377)
);

HB1xp67_ASAP7_75t_L g13378 ( 
.A(n_13108),
.Y(n_13378)
);

NAND2xp5_ASAP7_75t_L g13379 ( 
.A(n_13186),
.B(n_1841),
.Y(n_13379)
);

NAND3xp33_ASAP7_75t_L g13380 ( 
.A(n_13047),
.B(n_1844),
.C(n_1843),
.Y(n_13380)
);

AND2x2_ASAP7_75t_L g13381 ( 
.A(n_13209),
.B(n_1842),
.Y(n_13381)
);

AND2x2_ASAP7_75t_L g13382 ( 
.A(n_13141),
.B(n_1842),
.Y(n_13382)
);

AND2x2_ASAP7_75t_L g13383 ( 
.A(n_13144),
.B(n_1842),
.Y(n_13383)
);

NAND3xp33_ASAP7_75t_L g13384 ( 
.A(n_13051),
.B(n_1846),
.C(n_1845),
.Y(n_13384)
);

AOI221xp5_ASAP7_75t_L g13385 ( 
.A1(n_13030),
.A2(n_1846),
.B1(n_1843),
.B2(n_1845),
.C(n_1847),
.Y(n_13385)
);

AOI22xp33_ASAP7_75t_L g13386 ( 
.A1(n_13194),
.A2(n_1848),
.B1(n_1846),
.B2(n_1847),
.Y(n_13386)
);

AND2x2_ASAP7_75t_L g13387 ( 
.A(n_13158),
.B(n_1848),
.Y(n_13387)
);

NAND2xp5_ASAP7_75t_L g13388 ( 
.A(n_13188),
.B(n_1849),
.Y(n_13388)
);

NAND2xp5_ASAP7_75t_L g13389 ( 
.A(n_13102),
.B(n_1849),
.Y(n_13389)
);

OAI22xp5_ASAP7_75t_L g13390 ( 
.A1(n_13170),
.A2(n_1851),
.B1(n_1849),
.B2(n_1850),
.Y(n_13390)
);

AND2x2_ASAP7_75t_L g13391 ( 
.A(n_13168),
.B(n_1850),
.Y(n_13391)
);

NAND4xp25_ASAP7_75t_L g13392 ( 
.A(n_13178),
.B(n_1852),
.C(n_1850),
.D(n_1851),
.Y(n_13392)
);

AND2x2_ASAP7_75t_L g13393 ( 
.A(n_13177),
.B(n_1851),
.Y(n_13393)
);

NAND3xp33_ASAP7_75t_L g13394 ( 
.A(n_13069),
.B(n_1854),
.C(n_1853),
.Y(n_13394)
);

NAND2xp5_ASAP7_75t_L g13395 ( 
.A(n_13134),
.B(n_1852),
.Y(n_13395)
);

NAND2xp5_ASAP7_75t_L g13396 ( 
.A(n_13206),
.B(n_1852),
.Y(n_13396)
);

AND2x2_ASAP7_75t_L g13397 ( 
.A(n_13062),
.B(n_1853),
.Y(n_13397)
);

AOI221xp5_ASAP7_75t_L g13398 ( 
.A1(n_13033),
.A2(n_1856),
.B1(n_1854),
.B2(n_1855),
.C(n_1857),
.Y(n_13398)
);

NAND2xp5_ASAP7_75t_L g13399 ( 
.A(n_13210),
.B(n_1855),
.Y(n_13399)
);

OAI221xp5_ASAP7_75t_SL g13400 ( 
.A1(n_13205),
.A2(n_1857),
.B1(n_1855),
.B2(n_1856),
.C(n_1859),
.Y(n_13400)
);

NAND3xp33_ASAP7_75t_L g13401 ( 
.A(n_13075),
.B(n_1859),
.C(n_1857),
.Y(n_13401)
);

NAND2xp5_ASAP7_75t_L g13402 ( 
.A(n_13106),
.B(n_1856),
.Y(n_13402)
);

NAND2xp5_ASAP7_75t_L g13403 ( 
.A(n_13176),
.B(n_1859),
.Y(n_13403)
);

NAND2xp5_ASAP7_75t_L g13404 ( 
.A(n_13181),
.B(n_1860),
.Y(n_13404)
);

AND2x2_ASAP7_75t_L g13405 ( 
.A(n_13065),
.B(n_1861),
.Y(n_13405)
);

AND2x2_ASAP7_75t_L g13406 ( 
.A(n_13222),
.B(n_1861),
.Y(n_13406)
);

NAND3xp33_ASAP7_75t_L g13407 ( 
.A(n_13080),
.B(n_1864),
.C(n_1863),
.Y(n_13407)
);

NAND2xp5_ASAP7_75t_L g13408 ( 
.A(n_13201),
.B(n_1862),
.Y(n_13408)
);

AOI22xp33_ASAP7_75t_SL g13409 ( 
.A1(n_13081),
.A2(n_1864),
.B1(n_1862),
.B2(n_1863),
.Y(n_13409)
);

AND2x2_ASAP7_75t_L g13410 ( 
.A(n_13049),
.B(n_13050),
.Y(n_13410)
);

AND2x2_ASAP7_75t_SL g13411 ( 
.A(n_13054),
.B(n_1862),
.Y(n_13411)
);

NAND2xp5_ASAP7_75t_L g13412 ( 
.A(n_13136),
.B(n_1863),
.Y(n_13412)
);

NAND2xp5_ASAP7_75t_L g13413 ( 
.A(n_13195),
.B(n_1865),
.Y(n_13413)
);

AND2x2_ASAP7_75t_L g13414 ( 
.A(n_13064),
.B(n_1865),
.Y(n_13414)
);

NAND3xp33_ASAP7_75t_L g13415 ( 
.A(n_13192),
.B(n_13160),
.C(n_13156),
.Y(n_13415)
);

NAND2xp5_ASAP7_75t_L g13416 ( 
.A(n_13199),
.B(n_1865),
.Y(n_13416)
);

AND2x2_ASAP7_75t_L g13417 ( 
.A(n_13162),
.B(n_1866),
.Y(n_13417)
);

NOR2xp33_ASAP7_75t_L g13418 ( 
.A(n_13151),
.B(n_1866),
.Y(n_13418)
);

OAI21xp33_ASAP7_75t_L g13419 ( 
.A1(n_13132),
.A2(n_1866),
.B(n_1867),
.Y(n_13419)
);

NAND2xp5_ASAP7_75t_L g13420 ( 
.A(n_13143),
.B(n_13147),
.Y(n_13420)
);

AND2x2_ASAP7_75t_L g13421 ( 
.A(n_13243),
.B(n_13029),
.Y(n_13421)
);

AND2x2_ASAP7_75t_SL g13422 ( 
.A(n_13310),
.B(n_13046),
.Y(n_13422)
);

NAND2xp5_ASAP7_75t_L g13423 ( 
.A(n_13300),
.B(n_13098),
.Y(n_13423)
);

INVx1_ASAP7_75t_L g13424 ( 
.A(n_13321),
.Y(n_13424)
);

AND2x2_ASAP7_75t_L g13425 ( 
.A(n_13263),
.B(n_13087),
.Y(n_13425)
);

AND2x4_ASAP7_75t_SL g13426 ( 
.A(n_13378),
.B(n_13208),
.Y(n_13426)
);

AND2x2_ASAP7_75t_L g13427 ( 
.A(n_13246),
.B(n_13101),
.Y(n_13427)
);

INVx1_ASAP7_75t_L g13428 ( 
.A(n_13382),
.Y(n_13428)
);

AND2x2_ASAP7_75t_L g13429 ( 
.A(n_13320),
.B(n_13138),
.Y(n_13429)
);

AND2x2_ASAP7_75t_L g13430 ( 
.A(n_13318),
.B(n_13142),
.Y(n_13430)
);

AND2x2_ASAP7_75t_L g13431 ( 
.A(n_13332),
.B(n_13164),
.Y(n_13431)
);

AND2x2_ASAP7_75t_L g13432 ( 
.A(n_13250),
.B(n_13172),
.Y(n_13432)
);

AND2x2_ASAP7_75t_L g13433 ( 
.A(n_13262),
.B(n_13113),
.Y(n_13433)
);

NAND2xp5_ASAP7_75t_L g13434 ( 
.A(n_13359),
.B(n_13213),
.Y(n_13434)
);

INVx1_ASAP7_75t_L g13435 ( 
.A(n_13383),
.Y(n_13435)
);

INVx2_ASAP7_75t_L g13436 ( 
.A(n_13411),
.Y(n_13436)
);

INVx1_ASAP7_75t_L g13437 ( 
.A(n_13387),
.Y(n_13437)
);

INVx2_ASAP7_75t_L g13438 ( 
.A(n_13363),
.Y(n_13438)
);

INVx3_ASAP7_75t_L g13439 ( 
.A(n_13381),
.Y(n_13439)
);

AND2x2_ASAP7_75t_L g13440 ( 
.A(n_13224),
.B(n_13118),
.Y(n_13440)
);

HB1xp67_ASAP7_75t_L g13441 ( 
.A(n_13296),
.Y(n_13441)
);

INVx1_ASAP7_75t_L g13442 ( 
.A(n_13309),
.Y(n_13442)
);

INVx2_ASAP7_75t_L g13443 ( 
.A(n_13350),
.Y(n_13443)
);

AND2x2_ASAP7_75t_L g13444 ( 
.A(n_13352),
.B(n_13103),
.Y(n_13444)
);

INVx1_ASAP7_75t_L g13445 ( 
.A(n_13406),
.Y(n_13445)
);

NAND2xp5_ASAP7_75t_L g13446 ( 
.A(n_13364),
.B(n_13145),
.Y(n_13446)
);

AND2x2_ASAP7_75t_L g13447 ( 
.A(n_13315),
.B(n_13129),
.Y(n_13447)
);

NOR2xp33_ASAP7_75t_L g13448 ( 
.A(n_13229),
.B(n_13184),
.Y(n_13448)
);

INVx4_ASAP7_75t_L g13449 ( 
.A(n_13293),
.Y(n_13449)
);

HB1xp67_ASAP7_75t_L g13450 ( 
.A(n_13366),
.Y(n_13450)
);

INVx1_ASAP7_75t_L g13451 ( 
.A(n_13395),
.Y(n_13451)
);

INVx1_ASAP7_75t_L g13452 ( 
.A(n_13413),
.Y(n_13452)
);

INVx1_ASAP7_75t_L g13453 ( 
.A(n_13416),
.Y(n_13453)
);

INVx1_ASAP7_75t_L g13454 ( 
.A(n_13417),
.Y(n_13454)
);

AND2x2_ASAP7_75t_L g13455 ( 
.A(n_13253),
.B(n_13166),
.Y(n_13455)
);

HB1xp67_ASAP7_75t_L g13456 ( 
.A(n_13266),
.Y(n_13456)
);

AND2x2_ASAP7_75t_L g13457 ( 
.A(n_13325),
.B(n_13174),
.Y(n_13457)
);

INVx1_ASAP7_75t_L g13458 ( 
.A(n_13379),
.Y(n_13458)
);

HB1xp67_ASAP7_75t_L g13459 ( 
.A(n_13410),
.Y(n_13459)
);

AND2x4_ASAP7_75t_L g13460 ( 
.A(n_13343),
.B(n_13187),
.Y(n_13460)
);

INVx1_ASAP7_75t_L g13461 ( 
.A(n_13388),
.Y(n_13461)
);

INVx2_ASAP7_75t_L g13462 ( 
.A(n_13333),
.Y(n_13462)
);

AND2x4_ASAP7_75t_L g13463 ( 
.A(n_13226),
.B(n_13115),
.Y(n_13463)
);

AND2x2_ASAP7_75t_L g13464 ( 
.A(n_13257),
.B(n_13191),
.Y(n_13464)
);

AND2x2_ASAP7_75t_L g13465 ( 
.A(n_13268),
.B(n_13180),
.Y(n_13465)
);

NAND2xp5_ASAP7_75t_L g13466 ( 
.A(n_13264),
.B(n_13219),
.Y(n_13466)
);

INVx2_ASAP7_75t_L g13467 ( 
.A(n_13295),
.Y(n_13467)
);

INVx2_ASAP7_75t_SL g13468 ( 
.A(n_13228),
.Y(n_13468)
);

OR2x2_ASAP7_75t_L g13469 ( 
.A(n_13415),
.B(n_13128),
.Y(n_13469)
);

OR2x2_ASAP7_75t_L g13470 ( 
.A(n_13236),
.B(n_13214),
.Y(n_13470)
);

AND2x4_ASAP7_75t_L g13471 ( 
.A(n_13242),
.B(n_13127),
.Y(n_13471)
);

CKINVDCx16_ASAP7_75t_R g13472 ( 
.A(n_13338),
.Y(n_13472)
);

AND2x2_ASAP7_75t_L g13473 ( 
.A(n_13286),
.B(n_13369),
.Y(n_13473)
);

AOI22xp5_ASAP7_75t_L g13474 ( 
.A1(n_13256),
.A2(n_1869),
.B1(n_1867),
.B2(n_1868),
.Y(n_13474)
);

HB1xp67_ASAP7_75t_L g13475 ( 
.A(n_13312),
.Y(n_13475)
);

INVx3_ASAP7_75t_L g13476 ( 
.A(n_13391),
.Y(n_13476)
);

AND2x2_ASAP7_75t_L g13477 ( 
.A(n_13261),
.B(n_2432),
.Y(n_13477)
);

AND2x2_ASAP7_75t_L g13478 ( 
.A(n_13248),
.B(n_2434),
.Y(n_13478)
);

OR2x2_ASAP7_75t_L g13479 ( 
.A(n_13298),
.B(n_1867),
.Y(n_13479)
);

AND2x2_ASAP7_75t_L g13480 ( 
.A(n_13349),
.B(n_2435),
.Y(n_13480)
);

AND2x2_ASAP7_75t_L g13481 ( 
.A(n_13292),
.B(n_2435),
.Y(n_13481)
);

INVx2_ASAP7_75t_SL g13482 ( 
.A(n_13308),
.Y(n_13482)
);

NAND2xp5_ASAP7_75t_L g13483 ( 
.A(n_13358),
.B(n_1868),
.Y(n_13483)
);

INVx1_ASAP7_75t_L g13484 ( 
.A(n_13393),
.Y(n_13484)
);

AND2x2_ASAP7_75t_L g13485 ( 
.A(n_13245),
.B(n_13271),
.Y(n_13485)
);

AND2x2_ASAP7_75t_L g13486 ( 
.A(n_13244),
.B(n_2436),
.Y(n_13486)
);

INVx2_ASAP7_75t_L g13487 ( 
.A(n_13414),
.Y(n_13487)
);

NAND2xp5_ASAP7_75t_L g13488 ( 
.A(n_13322),
.B(n_1868),
.Y(n_13488)
);

BUFx2_ASAP7_75t_L g13489 ( 
.A(n_13287),
.Y(n_13489)
);

INVx2_ASAP7_75t_L g13490 ( 
.A(n_13299),
.Y(n_13490)
);

AND2x2_ASAP7_75t_L g13491 ( 
.A(n_13244),
.B(n_2439),
.Y(n_13491)
);

AND2x2_ASAP7_75t_L g13492 ( 
.A(n_13233),
.B(n_2441),
.Y(n_13492)
);

NOR2xp33_ASAP7_75t_SL g13493 ( 
.A(n_13324),
.B(n_1869),
.Y(n_13493)
);

INVx1_ASAP7_75t_L g13494 ( 
.A(n_13403),
.Y(n_13494)
);

INVx1_ASAP7_75t_L g13495 ( 
.A(n_13404),
.Y(n_13495)
);

BUFx3_ASAP7_75t_L g13496 ( 
.A(n_13389),
.Y(n_13496)
);

INVx2_ASAP7_75t_L g13497 ( 
.A(n_13249),
.Y(n_13497)
);

AND2x2_ASAP7_75t_L g13498 ( 
.A(n_13251),
.B(n_2442),
.Y(n_13498)
);

INVx3_ASAP7_75t_L g13499 ( 
.A(n_13397),
.Y(n_13499)
);

AND2x2_ASAP7_75t_L g13500 ( 
.A(n_13303),
.B(n_2442),
.Y(n_13500)
);

AND2x4_ASAP7_75t_L g13501 ( 
.A(n_13335),
.B(n_1869),
.Y(n_13501)
);

INVx1_ASAP7_75t_L g13502 ( 
.A(n_13316),
.Y(n_13502)
);

INVx2_ASAP7_75t_L g13503 ( 
.A(n_13405),
.Y(n_13503)
);

HB1xp67_ASAP7_75t_L g13504 ( 
.A(n_13279),
.Y(n_13504)
);

NAND2xp5_ASAP7_75t_L g13505 ( 
.A(n_13353),
.B(n_1870),
.Y(n_13505)
);

OAI22xp33_ASAP7_75t_L g13506 ( 
.A1(n_13225),
.A2(n_1872),
.B1(n_1870),
.B2(n_1871),
.Y(n_13506)
);

INVx2_ASAP7_75t_L g13507 ( 
.A(n_13373),
.Y(n_13507)
);

HB1xp67_ASAP7_75t_L g13508 ( 
.A(n_13259),
.Y(n_13508)
);

INVx1_ASAP7_75t_L g13509 ( 
.A(n_13337),
.Y(n_13509)
);

INVx2_ASAP7_75t_L g13510 ( 
.A(n_13368),
.Y(n_13510)
);

INVxp67_ASAP7_75t_L g13511 ( 
.A(n_13307),
.Y(n_13511)
);

BUFx2_ASAP7_75t_L g13512 ( 
.A(n_13290),
.Y(n_13512)
);

AND2x2_ASAP7_75t_L g13513 ( 
.A(n_13289),
.B(n_2445),
.Y(n_13513)
);

NOR2xp33_ASAP7_75t_L g13514 ( 
.A(n_13356),
.B(n_1871),
.Y(n_13514)
);

INVx1_ASAP7_75t_L g13515 ( 
.A(n_13408),
.Y(n_13515)
);

INVxp67_ASAP7_75t_L g13516 ( 
.A(n_13276),
.Y(n_13516)
);

AND2x2_ASAP7_75t_L g13517 ( 
.A(n_13232),
.B(n_2447),
.Y(n_13517)
);

AND2x2_ASAP7_75t_L g13518 ( 
.A(n_13240),
.B(n_2448),
.Y(n_13518)
);

INVx1_ASAP7_75t_L g13519 ( 
.A(n_13396),
.Y(n_13519)
);

INVx1_ASAP7_75t_L g13520 ( 
.A(n_13399),
.Y(n_13520)
);

NAND2xp5_ASAP7_75t_L g13521 ( 
.A(n_13319),
.B(n_1871),
.Y(n_13521)
);

INVx3_ASAP7_75t_L g13522 ( 
.A(n_13313),
.Y(n_13522)
);

NAND2xp5_ASAP7_75t_L g13523 ( 
.A(n_13247),
.B(n_13306),
.Y(n_13523)
);

AND2x2_ASAP7_75t_L g13524 ( 
.A(n_13230),
.B(n_2449),
.Y(n_13524)
);

INVx2_ASAP7_75t_L g13525 ( 
.A(n_13234),
.Y(n_13525)
);

NAND2xp5_ASAP7_75t_L g13526 ( 
.A(n_13346),
.B(n_1872),
.Y(n_13526)
);

OAI22xp5_ASAP7_75t_L g13527 ( 
.A1(n_13275),
.A2(n_1874),
.B1(n_1872),
.B2(n_1873),
.Y(n_13527)
);

AND2x2_ASAP7_75t_L g13528 ( 
.A(n_13370),
.B(n_2422),
.Y(n_13528)
);

AND2x4_ASAP7_75t_L g13529 ( 
.A(n_13277),
.B(n_1873),
.Y(n_13529)
);

HB1xp67_ASAP7_75t_L g13530 ( 
.A(n_13280),
.Y(n_13530)
);

AND2x2_ASAP7_75t_L g13531 ( 
.A(n_13223),
.B(n_2422),
.Y(n_13531)
);

BUFx2_ASAP7_75t_L g13532 ( 
.A(n_13231),
.Y(n_13532)
);

AND2x2_ASAP7_75t_L g13533 ( 
.A(n_13409),
.B(n_13334),
.Y(n_13533)
);

NAND2xp5_ASAP7_75t_L g13534 ( 
.A(n_13418),
.B(n_1873),
.Y(n_13534)
);

NAND2xp5_ASAP7_75t_L g13535 ( 
.A(n_13336),
.B(n_1874),
.Y(n_13535)
);

AND2x2_ASAP7_75t_L g13536 ( 
.A(n_13377),
.B(n_2425),
.Y(n_13536)
);

INVx1_ASAP7_75t_L g13537 ( 
.A(n_13376),
.Y(n_13537)
);

AND2x2_ASAP7_75t_L g13538 ( 
.A(n_13281),
.B(n_2425),
.Y(n_13538)
);

AND2x2_ASAP7_75t_L g13539 ( 
.A(n_13267),
.B(n_2425),
.Y(n_13539)
);

INVx2_ASAP7_75t_L g13540 ( 
.A(n_13235),
.Y(n_13540)
);

AND2x2_ASAP7_75t_L g13541 ( 
.A(n_13284),
.B(n_2426),
.Y(n_13541)
);

OR2x2_ASAP7_75t_L g13542 ( 
.A(n_13265),
.B(n_1875),
.Y(n_13542)
);

INVxp67_ASAP7_75t_L g13543 ( 
.A(n_13227),
.Y(n_13543)
);

HB1xp67_ASAP7_75t_L g13544 ( 
.A(n_13302),
.Y(n_13544)
);

AND2x2_ASAP7_75t_L g13545 ( 
.A(n_13344),
.B(n_2426),
.Y(n_13545)
);

NOR2xp33_ASAP7_75t_L g13546 ( 
.A(n_13392),
.B(n_1875),
.Y(n_13546)
);

OR2x2_ASAP7_75t_L g13547 ( 
.A(n_13323),
.B(n_1875),
.Y(n_13547)
);

INVx2_ASAP7_75t_L g13548 ( 
.A(n_13283),
.Y(n_13548)
);

INVx1_ASAP7_75t_L g13549 ( 
.A(n_13420),
.Y(n_13549)
);

AND2x2_ASAP7_75t_L g13550 ( 
.A(n_13351),
.B(n_2427),
.Y(n_13550)
);

OR2x2_ASAP7_75t_L g13551 ( 
.A(n_13304),
.B(n_1876),
.Y(n_13551)
);

AND2x2_ASAP7_75t_L g13552 ( 
.A(n_13238),
.B(n_2427),
.Y(n_13552)
);

AND2x4_ASAP7_75t_L g13553 ( 
.A(n_13297),
.B(n_13301),
.Y(n_13553)
);

INVx1_ASAP7_75t_L g13554 ( 
.A(n_13412),
.Y(n_13554)
);

NAND2xp5_ASAP7_75t_L g13555 ( 
.A(n_13340),
.B(n_1876),
.Y(n_13555)
);

INVx1_ASAP7_75t_L g13556 ( 
.A(n_13305),
.Y(n_13556)
);

OR2x2_ASAP7_75t_L g13557 ( 
.A(n_13326),
.B(n_1878),
.Y(n_13557)
);

INVx1_ASAP7_75t_L g13558 ( 
.A(n_13342),
.Y(n_13558)
);

INVx1_ASAP7_75t_L g13559 ( 
.A(n_13354),
.Y(n_13559)
);

INVx1_ASAP7_75t_L g13560 ( 
.A(n_13355),
.Y(n_13560)
);

AND2x2_ASAP7_75t_L g13561 ( 
.A(n_13282),
.B(n_2430),
.Y(n_13561)
);

INVx1_ASAP7_75t_L g13562 ( 
.A(n_13357),
.Y(n_13562)
);

INVx1_ASAP7_75t_L g13563 ( 
.A(n_13361),
.Y(n_13563)
);

INVx1_ASAP7_75t_L g13564 ( 
.A(n_13367),
.Y(n_13564)
);

INVx1_ASAP7_75t_SL g13565 ( 
.A(n_13239),
.Y(n_13565)
);

AND2x2_ASAP7_75t_L g13566 ( 
.A(n_13254),
.B(n_2430),
.Y(n_13566)
);

HB1xp67_ASAP7_75t_L g13567 ( 
.A(n_13270),
.Y(n_13567)
);

INVx1_ASAP7_75t_L g13568 ( 
.A(n_13371),
.Y(n_13568)
);

AND2x2_ASAP7_75t_L g13569 ( 
.A(n_13372),
.B(n_2430),
.Y(n_13569)
);

NAND2xp5_ASAP7_75t_L g13570 ( 
.A(n_13348),
.B(n_1879),
.Y(n_13570)
);

NAND2xp5_ASAP7_75t_L g13571 ( 
.A(n_13341),
.B(n_1879),
.Y(n_13571)
);

NAND2xp5_ASAP7_75t_L g13572 ( 
.A(n_13328),
.B(n_1879),
.Y(n_13572)
);

INVx1_ASAP7_75t_L g13573 ( 
.A(n_13374),
.Y(n_13573)
);

AND2x2_ASAP7_75t_L g13574 ( 
.A(n_13375),
.B(n_2434),
.Y(n_13574)
);

NAND2xp5_ASAP7_75t_L g13575 ( 
.A(n_13278),
.B(n_1880),
.Y(n_13575)
);

AND2x2_ASAP7_75t_L g13576 ( 
.A(n_13386),
.B(n_2436),
.Y(n_13576)
);

INVx1_ASAP7_75t_SL g13577 ( 
.A(n_13288),
.Y(n_13577)
);

INVx2_ASAP7_75t_L g13578 ( 
.A(n_13402),
.Y(n_13578)
);

OR2x2_ASAP7_75t_L g13579 ( 
.A(n_13365),
.B(n_1880),
.Y(n_13579)
);

AND2x2_ASAP7_75t_L g13580 ( 
.A(n_13273),
.B(n_2444),
.Y(n_13580)
);

INVx1_ASAP7_75t_L g13581 ( 
.A(n_13380),
.Y(n_13581)
);

INVx2_ASAP7_75t_SL g13582 ( 
.A(n_13345),
.Y(n_13582)
);

AND2x2_ASAP7_75t_L g13583 ( 
.A(n_13237),
.B(n_2444),
.Y(n_13583)
);

INVx1_ASAP7_75t_L g13584 ( 
.A(n_13384),
.Y(n_13584)
);

AND2x2_ASAP7_75t_SL g13585 ( 
.A(n_13255),
.B(n_1881),
.Y(n_13585)
);

BUFx2_ASAP7_75t_SL g13586 ( 
.A(n_13421),
.Y(n_13586)
);

INVx3_ASAP7_75t_L g13587 ( 
.A(n_13426),
.Y(n_13587)
);

INVx1_ASAP7_75t_L g13588 ( 
.A(n_13456),
.Y(n_13588)
);

HB1xp67_ASAP7_75t_L g13589 ( 
.A(n_13512),
.Y(n_13589)
);

INVx2_ASAP7_75t_L g13590 ( 
.A(n_13422),
.Y(n_13590)
);

INVx2_ASAP7_75t_L g13591 ( 
.A(n_13472),
.Y(n_13591)
);

INVx2_ASAP7_75t_L g13592 ( 
.A(n_13449),
.Y(n_13592)
);

OAI21x1_ASAP7_75t_L g13593 ( 
.A1(n_13486),
.A2(n_13360),
.B(n_13272),
.Y(n_13593)
);

NAND2x1_ASAP7_75t_L g13594 ( 
.A(n_13425),
.B(n_13427),
.Y(n_13594)
);

NAND2xp5_ASAP7_75t_SL g13595 ( 
.A(n_13489),
.B(n_13473),
.Y(n_13595)
);

INVx1_ASAP7_75t_L g13596 ( 
.A(n_13450),
.Y(n_13596)
);

INVx2_ASAP7_75t_L g13597 ( 
.A(n_13510),
.Y(n_13597)
);

INVx2_ASAP7_75t_L g13598 ( 
.A(n_13431),
.Y(n_13598)
);

INVx2_ASAP7_75t_L g13599 ( 
.A(n_13436),
.Y(n_13599)
);

INVx2_ASAP7_75t_SL g13600 ( 
.A(n_13459),
.Y(n_13600)
);

NAND3xp33_ASAP7_75t_SL g13601 ( 
.A(n_13491),
.B(n_13252),
.C(n_13311),
.Y(n_13601)
);

INVx2_ASAP7_75t_L g13602 ( 
.A(n_13499),
.Y(n_13602)
);

INVx1_ASAP7_75t_L g13603 ( 
.A(n_13441),
.Y(n_13603)
);

INVx2_ASAP7_75t_L g13604 ( 
.A(n_13432),
.Y(n_13604)
);

OAI21x1_ASAP7_75t_L g13605 ( 
.A1(n_13446),
.A2(n_13241),
.B(n_13294),
.Y(n_13605)
);

NAND3xp33_ASAP7_75t_L g13606 ( 
.A(n_13504),
.B(n_13531),
.C(n_13469),
.Y(n_13606)
);

INVx2_ASAP7_75t_L g13607 ( 
.A(n_13444),
.Y(n_13607)
);

INVx1_ASAP7_75t_L g13608 ( 
.A(n_13447),
.Y(n_13608)
);

INVx2_ASAP7_75t_L g13609 ( 
.A(n_13476),
.Y(n_13609)
);

INVx1_ASAP7_75t_L g13610 ( 
.A(n_13434),
.Y(n_13610)
);

OAI21xp33_ASAP7_75t_L g13611 ( 
.A1(n_13485),
.A2(n_13419),
.B(n_13260),
.Y(n_13611)
);

INVx2_ASAP7_75t_L g13612 ( 
.A(n_13429),
.Y(n_13612)
);

INVx1_ASAP7_75t_L g13613 ( 
.A(n_13544),
.Y(n_13613)
);

OA21x2_ASAP7_75t_L g13614 ( 
.A1(n_13516),
.A2(n_13401),
.B(n_13394),
.Y(n_13614)
);

INVx1_ASAP7_75t_L g13615 ( 
.A(n_13430),
.Y(n_13615)
);

OAI21xp5_ASAP7_75t_L g13616 ( 
.A1(n_13513),
.A2(n_13407),
.B(n_13269),
.Y(n_13616)
);

INVx2_ASAP7_75t_L g13617 ( 
.A(n_13507),
.Y(n_13617)
);

INVx2_ASAP7_75t_L g13618 ( 
.A(n_13496),
.Y(n_13618)
);

INVx1_ASAP7_75t_L g13619 ( 
.A(n_13572),
.Y(n_13619)
);

INVx1_ASAP7_75t_L g13620 ( 
.A(n_13445),
.Y(n_13620)
);

HB1xp67_ASAP7_75t_L g13621 ( 
.A(n_13455),
.Y(n_13621)
);

INVx2_ASAP7_75t_L g13622 ( 
.A(n_13438),
.Y(n_13622)
);

INVx2_ASAP7_75t_SL g13623 ( 
.A(n_13433),
.Y(n_13623)
);

NAND2xp5_ASAP7_75t_L g13624 ( 
.A(n_13428),
.B(n_13314),
.Y(n_13624)
);

INVx2_ASAP7_75t_L g13625 ( 
.A(n_13439),
.Y(n_13625)
);

OA21x2_ASAP7_75t_L g13626 ( 
.A1(n_13424),
.A2(n_13362),
.B(n_13327),
.Y(n_13626)
);

INVx1_ASAP7_75t_L g13627 ( 
.A(n_13435),
.Y(n_13627)
);

INVx1_ASAP7_75t_L g13628 ( 
.A(n_13437),
.Y(n_13628)
);

INVx1_ASAP7_75t_L g13629 ( 
.A(n_13566),
.Y(n_13629)
);

NAND2xp5_ASAP7_75t_L g13630 ( 
.A(n_13501),
.B(n_13330),
.Y(n_13630)
);

INVx2_ASAP7_75t_SL g13631 ( 
.A(n_13440),
.Y(n_13631)
);

INVx3_ASAP7_75t_L g13632 ( 
.A(n_13529),
.Y(n_13632)
);

NAND2xp5_ASAP7_75t_L g13633 ( 
.A(n_13454),
.B(n_13385),
.Y(n_13633)
);

OAI21xp5_ASAP7_75t_L g13634 ( 
.A1(n_13533),
.A2(n_13285),
.B(n_13258),
.Y(n_13634)
);

INVx2_ASAP7_75t_L g13635 ( 
.A(n_13443),
.Y(n_13635)
);

INVx2_ASAP7_75t_L g13636 ( 
.A(n_13462),
.Y(n_13636)
);

BUFx3_ASAP7_75t_L g13637 ( 
.A(n_13484),
.Y(n_13637)
);

AND2x2_ASAP7_75t_L g13638 ( 
.A(n_13465),
.B(n_13398),
.Y(n_13638)
);

INVx2_ASAP7_75t_L g13639 ( 
.A(n_13503),
.Y(n_13639)
);

INVx2_ASAP7_75t_L g13640 ( 
.A(n_13481),
.Y(n_13640)
);

NAND2xp5_ASAP7_75t_L g13641 ( 
.A(n_13487),
.B(n_13339),
.Y(n_13641)
);

NAND2xp5_ASAP7_75t_SL g13642 ( 
.A(n_13471),
.B(n_13274),
.Y(n_13642)
);

BUFx3_ASAP7_75t_L g13643 ( 
.A(n_13442),
.Y(n_13643)
);

INVx4_ASAP7_75t_L g13644 ( 
.A(n_13478),
.Y(n_13644)
);

BUFx2_ASAP7_75t_L g13645 ( 
.A(n_13457),
.Y(n_13645)
);

INVx4_ASAP7_75t_SL g13646 ( 
.A(n_13498),
.Y(n_13646)
);

INVx1_ASAP7_75t_L g13647 ( 
.A(n_13583),
.Y(n_13647)
);

INVx1_ASAP7_75t_L g13648 ( 
.A(n_13550),
.Y(n_13648)
);

INVx1_ASAP7_75t_L g13649 ( 
.A(n_13475),
.Y(n_13649)
);

NAND3xp33_ASAP7_75t_SL g13650 ( 
.A(n_13577),
.B(n_13291),
.C(n_13331),
.Y(n_13650)
);

INVx2_ASAP7_75t_L g13651 ( 
.A(n_13500),
.Y(n_13651)
);

INVx5_ASAP7_75t_L g13652 ( 
.A(n_13524),
.Y(n_13652)
);

INVx2_ASAP7_75t_L g13653 ( 
.A(n_13490),
.Y(n_13653)
);

NOR2x1p5_ASAP7_75t_L g13654 ( 
.A(n_13423),
.B(n_13347),
.Y(n_13654)
);

INVx2_ASAP7_75t_L g13655 ( 
.A(n_13553),
.Y(n_13655)
);

INVx2_ASAP7_75t_L g13656 ( 
.A(n_13479),
.Y(n_13656)
);

INVx2_ASAP7_75t_L g13657 ( 
.A(n_13536),
.Y(n_13657)
);

NAND3x1_ASAP7_75t_L g13658 ( 
.A(n_13464),
.B(n_13400),
.C(n_13317),
.Y(n_13658)
);

NAND3xp33_ASAP7_75t_SL g13659 ( 
.A(n_13523),
.B(n_13390),
.C(n_13329),
.Y(n_13659)
);

BUFx2_ASAP7_75t_L g13660 ( 
.A(n_13460),
.Y(n_13660)
);

BUFx2_ASAP7_75t_L g13661 ( 
.A(n_13477),
.Y(n_13661)
);

AND2x4_ASAP7_75t_L g13662 ( 
.A(n_13482),
.B(n_1881),
.Y(n_13662)
);

NAND2xp5_ASAP7_75t_SL g13663 ( 
.A(n_13468),
.B(n_1881),
.Y(n_13663)
);

INVx2_ASAP7_75t_L g13664 ( 
.A(n_13580),
.Y(n_13664)
);

INVx2_ASAP7_75t_L g13665 ( 
.A(n_13547),
.Y(n_13665)
);

INVx2_ASAP7_75t_L g13666 ( 
.A(n_13551),
.Y(n_13666)
);

INVx1_ASAP7_75t_L g13667 ( 
.A(n_13567),
.Y(n_13667)
);

INVx1_ASAP7_75t_SL g13668 ( 
.A(n_13470),
.Y(n_13668)
);

INVx1_ASAP7_75t_L g13669 ( 
.A(n_13526),
.Y(n_13669)
);

AO21x1_ASAP7_75t_SL g13670 ( 
.A1(n_13508),
.A2(n_1882),
.B(n_1883),
.Y(n_13670)
);

INVx1_ASAP7_75t_L g13671 ( 
.A(n_13534),
.Y(n_13671)
);

INVx1_ASAP7_75t_L g13672 ( 
.A(n_13483),
.Y(n_13672)
);

BUFx3_ASAP7_75t_L g13673 ( 
.A(n_13480),
.Y(n_13673)
);

OAI21x1_ASAP7_75t_L g13674 ( 
.A1(n_13575),
.A2(n_1882),
.B(n_1883),
.Y(n_13674)
);

INVx1_ASAP7_75t_L g13675 ( 
.A(n_13541),
.Y(n_13675)
);

OR2x6_ASAP7_75t_SL g13676 ( 
.A(n_13542),
.B(n_1882),
.Y(n_13676)
);

INVx1_ASAP7_75t_L g13677 ( 
.A(n_13488),
.Y(n_13677)
);

NAND2xp5_ASAP7_75t_L g13678 ( 
.A(n_13561),
.B(n_1883),
.Y(n_13678)
);

INVx2_ASAP7_75t_L g13679 ( 
.A(n_13557),
.Y(n_13679)
);

INVx3_ASAP7_75t_L g13680 ( 
.A(n_13463),
.Y(n_13680)
);

INVx1_ASAP7_75t_L g13681 ( 
.A(n_13521),
.Y(n_13681)
);

INVx2_ASAP7_75t_SL g13682 ( 
.A(n_13528),
.Y(n_13682)
);

INVx1_ASAP7_75t_L g13683 ( 
.A(n_13505),
.Y(n_13683)
);

INVx2_ASAP7_75t_L g13684 ( 
.A(n_13569),
.Y(n_13684)
);

OA21x2_ASAP7_75t_L g13685 ( 
.A1(n_13511),
.A2(n_2417),
.B(n_2416),
.Y(n_13685)
);

INVx2_ASAP7_75t_SL g13686 ( 
.A(n_13538),
.Y(n_13686)
);

AND2x4_ASAP7_75t_L g13687 ( 
.A(n_13539),
.B(n_1884),
.Y(n_13687)
);

BUFx2_ASAP7_75t_L g13688 ( 
.A(n_13518),
.Y(n_13688)
);

OAI21x1_ASAP7_75t_L g13689 ( 
.A1(n_13467),
.A2(n_1884),
.B(n_1885),
.Y(n_13689)
);

NAND3xp33_ASAP7_75t_SL g13690 ( 
.A(n_13565),
.B(n_1884),
.C(n_1885),
.Y(n_13690)
);

AOI21x1_ASAP7_75t_L g13691 ( 
.A1(n_13532),
.A2(n_2418),
.B(n_2417),
.Y(n_13691)
);

INVx1_ASAP7_75t_L g13692 ( 
.A(n_13574),
.Y(n_13692)
);

INVx2_ASAP7_75t_L g13693 ( 
.A(n_13579),
.Y(n_13693)
);

INVx2_ASAP7_75t_L g13694 ( 
.A(n_13582),
.Y(n_13694)
);

HB1xp67_ASAP7_75t_L g13695 ( 
.A(n_13492),
.Y(n_13695)
);

INVx2_ASAP7_75t_L g13696 ( 
.A(n_13497),
.Y(n_13696)
);

INVx1_ASAP7_75t_L g13697 ( 
.A(n_13552),
.Y(n_13697)
);

OA21x2_ASAP7_75t_L g13698 ( 
.A1(n_13474),
.A2(n_2419),
.B(n_2417),
.Y(n_13698)
);

OA21x2_ASAP7_75t_L g13699 ( 
.A1(n_13571),
.A2(n_13466),
.B(n_13581),
.Y(n_13699)
);

HB1xp67_ASAP7_75t_L g13700 ( 
.A(n_13530),
.Y(n_13700)
);

INVx1_ASAP7_75t_L g13701 ( 
.A(n_13535),
.Y(n_13701)
);

INVx4_ASAP7_75t_L g13702 ( 
.A(n_13517),
.Y(n_13702)
);

OR2x2_ASAP7_75t_L g13703 ( 
.A(n_13584),
.B(n_1885),
.Y(n_13703)
);

NOR2xp33_ASAP7_75t_L g13704 ( 
.A(n_13522),
.B(n_1886),
.Y(n_13704)
);

OAI21xp5_ASAP7_75t_SL g13705 ( 
.A1(n_13448),
.A2(n_1886),
.B(n_1887),
.Y(n_13705)
);

INVx1_ASAP7_75t_L g13706 ( 
.A(n_13555),
.Y(n_13706)
);

INVx1_ASAP7_75t_L g13707 ( 
.A(n_13570),
.Y(n_13707)
);

BUFx2_ASAP7_75t_L g13708 ( 
.A(n_13549),
.Y(n_13708)
);

AND4x1_ASAP7_75t_L g13709 ( 
.A(n_13493),
.B(n_13514),
.C(n_13546),
.D(n_13461),
.Y(n_13709)
);

AND2x2_ASAP7_75t_L g13710 ( 
.A(n_13556),
.B(n_1886),
.Y(n_13710)
);

INVx1_ASAP7_75t_L g13711 ( 
.A(n_13545),
.Y(n_13711)
);

INVx2_ASAP7_75t_L g13712 ( 
.A(n_13578),
.Y(n_13712)
);

INVx1_ASAP7_75t_L g13713 ( 
.A(n_13502),
.Y(n_13713)
);

INVx1_ASAP7_75t_SL g13714 ( 
.A(n_13585),
.Y(n_13714)
);

INVx1_ASAP7_75t_L g13715 ( 
.A(n_13509),
.Y(n_13715)
);

NAND2xp5_ASAP7_75t_SL g13716 ( 
.A(n_13506),
.B(n_1887),
.Y(n_13716)
);

HB1xp67_ASAP7_75t_L g13717 ( 
.A(n_13527),
.Y(n_13717)
);

INVx5_ASAP7_75t_L g13718 ( 
.A(n_13525),
.Y(n_13718)
);

NAND2xp5_ASAP7_75t_L g13719 ( 
.A(n_13652),
.B(n_13543),
.Y(n_13719)
);

INVx2_ASAP7_75t_L g13720 ( 
.A(n_13587),
.Y(n_13720)
);

AND2x2_ASAP7_75t_L g13721 ( 
.A(n_13586),
.B(n_13558),
.Y(n_13721)
);

AND2x2_ASAP7_75t_L g13722 ( 
.A(n_13621),
.B(n_13559),
.Y(n_13722)
);

INVx1_ASAP7_75t_L g13723 ( 
.A(n_13661),
.Y(n_13723)
);

NAND2x1p5_ASAP7_75t_L g13724 ( 
.A(n_13591),
.B(n_13515),
.Y(n_13724)
);

INVx1_ASAP7_75t_L g13725 ( 
.A(n_13645),
.Y(n_13725)
);

INVx2_ASAP7_75t_L g13726 ( 
.A(n_13652),
.Y(n_13726)
);

AND2x2_ASAP7_75t_L g13727 ( 
.A(n_13631),
.B(n_13560),
.Y(n_13727)
);

OR2x2_ASAP7_75t_L g13728 ( 
.A(n_13589),
.B(n_13562),
.Y(n_13728)
);

AND2x2_ASAP7_75t_L g13729 ( 
.A(n_13623),
.B(n_13563),
.Y(n_13729)
);

INVx1_ASAP7_75t_L g13730 ( 
.A(n_13660),
.Y(n_13730)
);

INVx1_ASAP7_75t_L g13731 ( 
.A(n_13700),
.Y(n_13731)
);

OR2x2_ASAP7_75t_L g13732 ( 
.A(n_13607),
.B(n_13564),
.Y(n_13732)
);

INVx1_ASAP7_75t_L g13733 ( 
.A(n_13691),
.Y(n_13733)
);

HB1xp67_ASAP7_75t_L g13734 ( 
.A(n_13594),
.Y(n_13734)
);

INVx1_ASAP7_75t_L g13735 ( 
.A(n_13612),
.Y(n_13735)
);

OR2x2_ASAP7_75t_L g13736 ( 
.A(n_13598),
.B(n_13568),
.Y(n_13736)
);

INVx1_ASAP7_75t_SL g13737 ( 
.A(n_13646),
.Y(n_13737)
);

INVx1_ASAP7_75t_L g13738 ( 
.A(n_13608),
.Y(n_13738)
);

INVx2_ASAP7_75t_L g13739 ( 
.A(n_13646),
.Y(n_13739)
);

INVx2_ASAP7_75t_L g13740 ( 
.A(n_13687),
.Y(n_13740)
);

NAND2xp5_ASAP7_75t_L g13741 ( 
.A(n_13644),
.B(n_13686),
.Y(n_13741)
);

OR2x2_ASAP7_75t_L g13742 ( 
.A(n_13600),
.B(n_13573),
.Y(n_13742)
);

AND2x2_ASAP7_75t_L g13743 ( 
.A(n_13604),
.B(n_13458),
.Y(n_13743)
);

INVx2_ASAP7_75t_L g13744 ( 
.A(n_13685),
.Y(n_13744)
);

AND2x2_ASAP7_75t_L g13745 ( 
.A(n_13680),
.B(n_13494),
.Y(n_13745)
);

NAND2xp5_ASAP7_75t_L g13746 ( 
.A(n_13682),
.B(n_13495),
.Y(n_13746)
);

INVx1_ASAP7_75t_SL g13747 ( 
.A(n_13668),
.Y(n_13747)
);

AND2x2_ASAP7_75t_L g13748 ( 
.A(n_13615),
.B(n_13451),
.Y(n_13748)
);

INVx1_ASAP7_75t_L g13749 ( 
.A(n_13688),
.Y(n_13749)
);

AND2x2_ASAP7_75t_L g13750 ( 
.A(n_13595),
.B(n_13452),
.Y(n_13750)
);

AND2x2_ASAP7_75t_L g13751 ( 
.A(n_13618),
.B(n_13453),
.Y(n_13751)
);

OR2x2_ASAP7_75t_L g13752 ( 
.A(n_13606),
.B(n_13548),
.Y(n_13752)
);

NOR2x1p5_ASAP7_75t_L g13753 ( 
.A(n_13643),
.B(n_13520),
.Y(n_13753)
);

NAND2xp5_ASAP7_75t_SL g13754 ( 
.A(n_13718),
.B(n_13540),
.Y(n_13754)
);

NAND2xp5_ASAP7_75t_L g13755 ( 
.A(n_13647),
.B(n_13519),
.Y(n_13755)
);

AND2x2_ASAP7_75t_L g13756 ( 
.A(n_13592),
.B(n_13537),
.Y(n_13756)
);

INVx1_ASAP7_75t_L g13757 ( 
.A(n_13695),
.Y(n_13757)
);

NAND2xp5_ASAP7_75t_L g13758 ( 
.A(n_13662),
.B(n_13554),
.Y(n_13758)
);

INVx1_ASAP7_75t_L g13759 ( 
.A(n_13664),
.Y(n_13759)
);

OR2x2_ASAP7_75t_L g13760 ( 
.A(n_13596),
.B(n_13576),
.Y(n_13760)
);

INVx1_ASAP7_75t_L g13761 ( 
.A(n_13678),
.Y(n_13761)
);

INVx1_ASAP7_75t_L g13762 ( 
.A(n_13675),
.Y(n_13762)
);

NAND2x1p5_ASAP7_75t_L g13763 ( 
.A(n_13632),
.B(n_1887),
.Y(n_13763)
);

INVx1_ASAP7_75t_L g13764 ( 
.A(n_13676),
.Y(n_13764)
);

NAND2x1p5_ASAP7_75t_L g13765 ( 
.A(n_13694),
.B(n_1888),
.Y(n_13765)
);

INVx2_ASAP7_75t_L g13766 ( 
.A(n_13673),
.Y(n_13766)
);

INVxp67_ASAP7_75t_L g13767 ( 
.A(n_13670),
.Y(n_13767)
);

INVxp67_ASAP7_75t_SL g13768 ( 
.A(n_13658),
.Y(n_13768)
);

AND2x2_ASAP7_75t_L g13769 ( 
.A(n_13602),
.B(n_1888),
.Y(n_13769)
);

NAND2xp5_ASAP7_75t_L g13770 ( 
.A(n_13684),
.B(n_1888),
.Y(n_13770)
);

INVx1_ASAP7_75t_L g13771 ( 
.A(n_13640),
.Y(n_13771)
);

AND2x2_ASAP7_75t_L g13772 ( 
.A(n_13625),
.B(n_1889),
.Y(n_13772)
);

INVx1_ASAP7_75t_L g13773 ( 
.A(n_13708),
.Y(n_13773)
);

INVx2_ASAP7_75t_L g13774 ( 
.A(n_13651),
.Y(n_13774)
);

OR2x2_ASAP7_75t_L g13775 ( 
.A(n_13603),
.B(n_2424),
.Y(n_13775)
);

NAND2xp5_ASAP7_75t_L g13776 ( 
.A(n_13692),
.B(n_1889),
.Y(n_13776)
);

INVxp67_ASAP7_75t_SL g13777 ( 
.A(n_13642),
.Y(n_13777)
);

INVx2_ASAP7_75t_L g13778 ( 
.A(n_13699),
.Y(n_13778)
);

INVx1_ASAP7_75t_L g13779 ( 
.A(n_13648),
.Y(n_13779)
);

INVx1_ASAP7_75t_L g13780 ( 
.A(n_13697),
.Y(n_13780)
);

INVx1_ASAP7_75t_L g13781 ( 
.A(n_13710),
.Y(n_13781)
);

AND3x1_ASAP7_75t_L g13782 ( 
.A(n_13609),
.B(n_1889),
.C(n_1890),
.Y(n_13782)
);

AND2x2_ASAP7_75t_L g13783 ( 
.A(n_13637),
.B(n_1890),
.Y(n_13783)
);

NOR2xp33_ASAP7_75t_L g13784 ( 
.A(n_13702),
.B(n_1890),
.Y(n_13784)
);

INVx1_ASAP7_75t_L g13785 ( 
.A(n_13655),
.Y(n_13785)
);

INVx1_ASAP7_75t_L g13786 ( 
.A(n_13665),
.Y(n_13786)
);

INVx1_ASAP7_75t_L g13787 ( 
.A(n_13666),
.Y(n_13787)
);

AND2x4_ASAP7_75t_L g13788 ( 
.A(n_13649),
.B(n_13613),
.Y(n_13788)
);

INVx1_ASAP7_75t_L g13789 ( 
.A(n_13679),
.Y(n_13789)
);

NOR2xp67_ASAP7_75t_SL g13790 ( 
.A(n_13667),
.B(n_1891),
.Y(n_13790)
);

INVx2_ASAP7_75t_SL g13791 ( 
.A(n_13590),
.Y(n_13791)
);

NAND2xp5_ASAP7_75t_L g13792 ( 
.A(n_13705),
.B(n_13619),
.Y(n_13792)
);

AND2x2_ASAP7_75t_L g13793 ( 
.A(n_13588),
.B(n_1891),
.Y(n_13793)
);

NAND2xp5_ASAP7_75t_L g13794 ( 
.A(n_13656),
.B(n_1891),
.Y(n_13794)
);

INVx2_ASAP7_75t_L g13795 ( 
.A(n_13698),
.Y(n_13795)
);

NAND2xp5_ASAP7_75t_L g13796 ( 
.A(n_13629),
.B(n_1892),
.Y(n_13796)
);

OR2x2_ASAP7_75t_L g13797 ( 
.A(n_13663),
.B(n_2429),
.Y(n_13797)
);

OR2x6_ASAP7_75t_L g13798 ( 
.A(n_13597),
.B(n_13599),
.Y(n_13798)
);

INVx1_ASAP7_75t_L g13799 ( 
.A(n_13614),
.Y(n_13799)
);

AND2x2_ASAP7_75t_L g13800 ( 
.A(n_13610),
.B(n_1892),
.Y(n_13800)
);

OR2x2_ASAP7_75t_L g13801 ( 
.A(n_13620),
.B(n_2429),
.Y(n_13801)
);

BUFx2_ASAP7_75t_L g13802 ( 
.A(n_13622),
.Y(n_13802)
);

AND2x2_ASAP7_75t_L g13803 ( 
.A(n_13627),
.B(n_1892),
.Y(n_13803)
);

AND2x4_ASAP7_75t_L g13804 ( 
.A(n_13635),
.B(n_1894),
.Y(n_13804)
);

AND2x2_ASAP7_75t_L g13805 ( 
.A(n_13628),
.B(n_1894),
.Y(n_13805)
);

NAND2xp5_ASAP7_75t_L g13806 ( 
.A(n_13718),
.B(n_1894),
.Y(n_13806)
);

INVx2_ASAP7_75t_L g13807 ( 
.A(n_13689),
.Y(n_13807)
);

AND2x2_ASAP7_75t_L g13808 ( 
.A(n_13636),
.B(n_1895),
.Y(n_13808)
);

INVx1_ASAP7_75t_L g13809 ( 
.A(n_13703),
.Y(n_13809)
);

INVx2_ASAP7_75t_L g13810 ( 
.A(n_13674),
.Y(n_13810)
);

NAND2xp5_ASAP7_75t_L g13811 ( 
.A(n_13638),
.B(n_1895),
.Y(n_13811)
);

INVx1_ASAP7_75t_L g13812 ( 
.A(n_13653),
.Y(n_13812)
);

INVx2_ASAP7_75t_L g13813 ( 
.A(n_13657),
.Y(n_13813)
);

NAND2xp5_ASAP7_75t_L g13814 ( 
.A(n_13704),
.B(n_1895),
.Y(n_13814)
);

OR2x2_ASAP7_75t_L g13815 ( 
.A(n_13713),
.B(n_2444),
.Y(n_13815)
);

NAND2xp5_ASAP7_75t_L g13816 ( 
.A(n_13671),
.B(n_13634),
.Y(n_13816)
);

NOR2x1p5_ASAP7_75t_L g13817 ( 
.A(n_13715),
.B(n_1896),
.Y(n_13817)
);

INVx3_ASAP7_75t_L g13818 ( 
.A(n_13639),
.Y(n_13818)
);

NAND2x1p5_ASAP7_75t_L g13819 ( 
.A(n_13709),
.B(n_1896),
.Y(n_13819)
);

INVx1_ASAP7_75t_L g13820 ( 
.A(n_13714),
.Y(n_13820)
);

INVx2_ASAP7_75t_SL g13821 ( 
.A(n_13617),
.Y(n_13821)
);

OR2x2_ASAP7_75t_L g13822 ( 
.A(n_13717),
.B(n_2448),
.Y(n_13822)
);

AND2x2_ASAP7_75t_L g13823 ( 
.A(n_13654),
.B(n_1896),
.Y(n_13823)
);

INVx1_ASAP7_75t_L g13824 ( 
.A(n_13690),
.Y(n_13824)
);

AND2x2_ASAP7_75t_L g13825 ( 
.A(n_13669),
.B(n_1897),
.Y(n_13825)
);

INVx2_ASAP7_75t_L g13826 ( 
.A(n_13696),
.Y(n_13826)
);

NAND2xp5_ASAP7_75t_L g13827 ( 
.A(n_13693),
.B(n_1897),
.Y(n_13827)
);

AND2x2_ASAP7_75t_L g13828 ( 
.A(n_13616),
.B(n_13626),
.Y(n_13828)
);

INVx1_ASAP7_75t_L g13829 ( 
.A(n_13624),
.Y(n_13829)
);

OR2x2_ASAP7_75t_L g13830 ( 
.A(n_13659),
.B(n_2412),
.Y(n_13830)
);

INVx1_ASAP7_75t_L g13831 ( 
.A(n_13641),
.Y(n_13831)
);

INVx1_ASAP7_75t_L g13832 ( 
.A(n_13593),
.Y(n_13832)
);

AND2x2_ASAP7_75t_L g13833 ( 
.A(n_13605),
.B(n_1897),
.Y(n_13833)
);

AND2x2_ASAP7_75t_L g13834 ( 
.A(n_13683),
.B(n_1898),
.Y(n_13834)
);

INVx2_ASAP7_75t_L g13835 ( 
.A(n_13712),
.Y(n_13835)
);

INVx2_ASAP7_75t_L g13836 ( 
.A(n_13711),
.Y(n_13836)
);

OR2x2_ASAP7_75t_L g13837 ( 
.A(n_13650),
.B(n_2414),
.Y(n_13837)
);

NAND2xp5_ASAP7_75t_L g13838 ( 
.A(n_13611),
.B(n_1899),
.Y(n_13838)
);

INVx2_ASAP7_75t_SL g13839 ( 
.A(n_13630),
.Y(n_13839)
);

OR2x2_ASAP7_75t_L g13840 ( 
.A(n_13601),
.B(n_13633),
.Y(n_13840)
);

INVx2_ASAP7_75t_L g13841 ( 
.A(n_13681),
.Y(n_13841)
);

AND2x2_ASAP7_75t_L g13842 ( 
.A(n_13672),
.B(n_13677),
.Y(n_13842)
);

AND2x2_ASAP7_75t_L g13843 ( 
.A(n_13706),
.B(n_1899),
.Y(n_13843)
);

AND2x2_ASAP7_75t_L g13844 ( 
.A(n_13707),
.B(n_1900),
.Y(n_13844)
);

AND2x2_ASAP7_75t_L g13845 ( 
.A(n_13701),
.B(n_1900),
.Y(n_13845)
);

OR2x2_ASAP7_75t_L g13846 ( 
.A(n_13716),
.B(n_2415),
.Y(n_13846)
);

OR2x2_ASAP7_75t_L g13847 ( 
.A(n_13645),
.B(n_2416),
.Y(n_13847)
);

OR2x6_ASAP7_75t_L g13848 ( 
.A(n_13591),
.B(n_1900),
.Y(n_13848)
);

INVx1_ASAP7_75t_L g13849 ( 
.A(n_13777),
.Y(n_13849)
);

INVx3_ASAP7_75t_L g13850 ( 
.A(n_13720),
.Y(n_13850)
);

INVx2_ASAP7_75t_L g13851 ( 
.A(n_13763),
.Y(n_13851)
);

AND2x2_ASAP7_75t_L g13852 ( 
.A(n_13747),
.B(n_1901),
.Y(n_13852)
);

AND2x2_ASAP7_75t_L g13853 ( 
.A(n_13767),
.B(n_1901),
.Y(n_13853)
);

HB1xp67_ASAP7_75t_L g13854 ( 
.A(n_13848),
.Y(n_13854)
);

INVx2_ASAP7_75t_L g13855 ( 
.A(n_13765),
.Y(n_13855)
);

INVx2_ASAP7_75t_SL g13856 ( 
.A(n_13753),
.Y(n_13856)
);

AND2x2_ASAP7_75t_L g13857 ( 
.A(n_13737),
.B(n_1901),
.Y(n_13857)
);

OR2x2_ASAP7_75t_L g13858 ( 
.A(n_13719),
.B(n_13802),
.Y(n_13858)
);

NAND2xp5_ASAP7_75t_L g13859 ( 
.A(n_13764),
.B(n_1902),
.Y(n_13859)
);

NAND3xp33_ASAP7_75t_L g13860 ( 
.A(n_13828),
.B(n_1902),
.C(n_1904),
.Y(n_13860)
);

O2A1O1Ixp33_ASAP7_75t_L g13861 ( 
.A1(n_13778),
.A2(n_1905),
.B(n_1902),
.C(n_1904),
.Y(n_13861)
);

NAND2xp5_ASAP7_75t_L g13862 ( 
.A(n_13744),
.B(n_1906),
.Y(n_13862)
);

AND2x2_ASAP7_75t_L g13863 ( 
.A(n_13722),
.B(n_1906),
.Y(n_13863)
);

NAND2xp5_ASAP7_75t_L g13864 ( 
.A(n_13804),
.B(n_1906),
.Y(n_13864)
);

INVx2_ASAP7_75t_L g13865 ( 
.A(n_13819),
.Y(n_13865)
);

AND2x2_ASAP7_75t_L g13866 ( 
.A(n_13750),
.B(n_1907),
.Y(n_13866)
);

AND2x2_ASAP7_75t_L g13867 ( 
.A(n_13721),
.B(n_1907),
.Y(n_13867)
);

INVx1_ASAP7_75t_L g13868 ( 
.A(n_13847),
.Y(n_13868)
);

INVx1_ASAP7_75t_L g13869 ( 
.A(n_13848),
.Y(n_13869)
);

INVx1_ASAP7_75t_L g13870 ( 
.A(n_13840),
.Y(n_13870)
);

AOI221xp5_ASAP7_75t_L g13871 ( 
.A1(n_13799),
.A2(n_13832),
.B1(n_13733),
.B2(n_13768),
.C(n_13816),
.Y(n_13871)
);

AND2x2_ASAP7_75t_L g13872 ( 
.A(n_13743),
.B(n_1907),
.Y(n_13872)
);

NAND2xp5_ASAP7_75t_L g13873 ( 
.A(n_13734),
.B(n_1908),
.Y(n_13873)
);

NAND2xp5_ASAP7_75t_L g13874 ( 
.A(n_13739),
.B(n_1908),
.Y(n_13874)
);

NAND2xp5_ASAP7_75t_L g13875 ( 
.A(n_13818),
.B(n_1909),
.Y(n_13875)
);

INVx1_ASAP7_75t_L g13876 ( 
.A(n_13782),
.Y(n_13876)
);

AND2x2_ASAP7_75t_L g13877 ( 
.A(n_13729),
.B(n_1909),
.Y(n_13877)
);

NAND2xp5_ASAP7_75t_L g13878 ( 
.A(n_13817),
.B(n_1909),
.Y(n_13878)
);

INVx1_ASAP7_75t_L g13879 ( 
.A(n_13822),
.Y(n_13879)
);

OR2x2_ASAP7_75t_L g13880 ( 
.A(n_13724),
.B(n_1910),
.Y(n_13880)
);

AND2x2_ASAP7_75t_L g13881 ( 
.A(n_13745),
.B(n_13723),
.Y(n_13881)
);

AND2x2_ASAP7_75t_L g13882 ( 
.A(n_13727),
.B(n_1910),
.Y(n_13882)
);

AND2x2_ASAP7_75t_L g13883 ( 
.A(n_13730),
.B(n_1910),
.Y(n_13883)
);

AND2x2_ASAP7_75t_L g13884 ( 
.A(n_13725),
.B(n_1911),
.Y(n_13884)
);

AND2x4_ASAP7_75t_SL g13885 ( 
.A(n_13766),
.B(n_1911),
.Y(n_13885)
);

NOR2xp33_ASAP7_75t_L g13886 ( 
.A(n_13726),
.B(n_13785),
.Y(n_13886)
);

NAND2xp5_ASAP7_75t_L g13887 ( 
.A(n_13781),
.B(n_1912),
.Y(n_13887)
);

NAND2x1_ASAP7_75t_SL g13888 ( 
.A(n_13773),
.B(n_1912),
.Y(n_13888)
);

AND2x2_ASAP7_75t_L g13889 ( 
.A(n_13749),
.B(n_1912),
.Y(n_13889)
);

INVx1_ASAP7_75t_L g13890 ( 
.A(n_13824),
.Y(n_13890)
);

OR2x2_ASAP7_75t_L g13891 ( 
.A(n_13728),
.B(n_1913),
.Y(n_13891)
);

AND2x2_ASAP7_75t_L g13892 ( 
.A(n_13751),
.B(n_1913),
.Y(n_13892)
);

NAND3xp33_ASAP7_75t_L g13893 ( 
.A(n_13790),
.B(n_1913),
.C(n_1914),
.Y(n_13893)
);

NAND2xp5_ASAP7_75t_L g13894 ( 
.A(n_13783),
.B(n_1914),
.Y(n_13894)
);

OR2x2_ASAP7_75t_L g13895 ( 
.A(n_13752),
.B(n_1914),
.Y(n_13895)
);

OR2x2_ASAP7_75t_L g13896 ( 
.A(n_13741),
.B(n_1915),
.Y(n_13896)
);

OR2x2_ASAP7_75t_L g13897 ( 
.A(n_13736),
.B(n_1915),
.Y(n_13897)
);

INVx1_ASAP7_75t_L g13898 ( 
.A(n_13833),
.Y(n_13898)
);

NAND2xp5_ASAP7_75t_L g13899 ( 
.A(n_13808),
.B(n_1915),
.Y(n_13899)
);

INVx1_ASAP7_75t_L g13900 ( 
.A(n_13795),
.Y(n_13900)
);

INVx2_ASAP7_75t_L g13901 ( 
.A(n_13740),
.Y(n_13901)
);

AND2x4_ASAP7_75t_L g13902 ( 
.A(n_13839),
.B(n_1916),
.Y(n_13902)
);

INVx1_ASAP7_75t_L g13903 ( 
.A(n_13806),
.Y(n_13903)
);

AND2x2_ASAP7_75t_L g13904 ( 
.A(n_13748),
.B(n_1916),
.Y(n_13904)
);

INVxp67_ASAP7_75t_L g13905 ( 
.A(n_13784),
.Y(n_13905)
);

AND2x4_ASAP7_75t_SL g13906 ( 
.A(n_13820),
.B(n_1916),
.Y(n_13906)
);

INVxp67_ASAP7_75t_L g13907 ( 
.A(n_13798),
.Y(n_13907)
);

INVx1_ASAP7_75t_L g13908 ( 
.A(n_13798),
.Y(n_13908)
);

AOI22xp33_ASAP7_75t_L g13909 ( 
.A1(n_13809),
.A2(n_1919),
.B1(n_1917),
.B2(n_1918),
.Y(n_13909)
);

INVx1_ASAP7_75t_L g13910 ( 
.A(n_13837),
.Y(n_13910)
);

AND2x2_ASAP7_75t_L g13911 ( 
.A(n_13756),
.B(n_1917),
.Y(n_13911)
);

INVx2_ASAP7_75t_L g13912 ( 
.A(n_13801),
.Y(n_13912)
);

INVx1_ASAP7_75t_L g13913 ( 
.A(n_13823),
.Y(n_13913)
);

OR2x2_ASAP7_75t_L g13914 ( 
.A(n_13760),
.B(n_1917),
.Y(n_13914)
);

NAND2xp5_ASAP7_75t_L g13915 ( 
.A(n_13834),
.B(n_1918),
.Y(n_13915)
);

INVx1_ASAP7_75t_L g13916 ( 
.A(n_13811),
.Y(n_13916)
);

BUFx2_ASAP7_75t_L g13917 ( 
.A(n_13774),
.Y(n_13917)
);

INVx1_ASAP7_75t_L g13918 ( 
.A(n_13792),
.Y(n_13918)
);

INVx2_ASAP7_75t_SL g13919 ( 
.A(n_13742),
.Y(n_13919)
);

NAND2xp5_ASAP7_75t_L g13920 ( 
.A(n_13831),
.B(n_1918),
.Y(n_13920)
);

OR2x2_ASAP7_75t_L g13921 ( 
.A(n_13732),
.B(n_1919),
.Y(n_13921)
);

INVx1_ASAP7_75t_L g13922 ( 
.A(n_13843),
.Y(n_13922)
);

AND2x2_ASAP7_75t_L g13923 ( 
.A(n_13757),
.B(n_1919),
.Y(n_13923)
);

HB1xp67_ASAP7_75t_L g13924 ( 
.A(n_13803),
.Y(n_13924)
);

NOR2x1_ASAP7_75t_L g13925 ( 
.A(n_13754),
.B(n_1920),
.Y(n_13925)
);

NOR2xp33_ASAP7_75t_L g13926 ( 
.A(n_13826),
.B(n_2421),
.Y(n_13926)
);

AND2x2_ASAP7_75t_L g13927 ( 
.A(n_13735),
.B(n_1920),
.Y(n_13927)
);

NAND2xp5_ASAP7_75t_L g13928 ( 
.A(n_13844),
.B(n_1920),
.Y(n_13928)
);

INVx1_ASAP7_75t_L g13929 ( 
.A(n_13758),
.Y(n_13929)
);

OR2x2_ASAP7_75t_L g13930 ( 
.A(n_13746),
.B(n_1921),
.Y(n_13930)
);

NAND2xp5_ASAP7_75t_L g13931 ( 
.A(n_13825),
.B(n_1921),
.Y(n_13931)
);

NOR2xp33_ASAP7_75t_L g13932 ( 
.A(n_13835),
.B(n_13812),
.Y(n_13932)
);

AND2x4_ASAP7_75t_L g13933 ( 
.A(n_13836),
.B(n_1921),
.Y(n_13933)
);

INVx1_ASAP7_75t_L g13934 ( 
.A(n_13845),
.Y(n_13934)
);

AND2x2_ASAP7_75t_L g13935 ( 
.A(n_13779),
.B(n_1922),
.Y(n_13935)
);

NOR2x1_ASAP7_75t_L g13936 ( 
.A(n_13731),
.B(n_1922),
.Y(n_13936)
);

INVx1_ASAP7_75t_L g13937 ( 
.A(n_13805),
.Y(n_13937)
);

INVx1_ASAP7_75t_L g13938 ( 
.A(n_13800),
.Y(n_13938)
);

INVxp67_ASAP7_75t_SL g13939 ( 
.A(n_13755),
.Y(n_13939)
);

OR2x2_ASAP7_75t_L g13940 ( 
.A(n_13775),
.B(n_1922),
.Y(n_13940)
);

O2A1O1Ixp33_ASAP7_75t_L g13941 ( 
.A1(n_13830),
.A2(n_1925),
.B(n_1923),
.C(n_1924),
.Y(n_13941)
);

INVx1_ASAP7_75t_L g13942 ( 
.A(n_13769),
.Y(n_13942)
);

OR2x2_ASAP7_75t_L g13943 ( 
.A(n_13780),
.B(n_1923),
.Y(n_13943)
);

INVx1_ASAP7_75t_L g13944 ( 
.A(n_13772),
.Y(n_13944)
);

NAND2xp5_ASAP7_75t_L g13945 ( 
.A(n_13842),
.B(n_1923),
.Y(n_13945)
);

INVx2_ASAP7_75t_SL g13946 ( 
.A(n_13793),
.Y(n_13946)
);

NAND2xp5_ASAP7_75t_L g13947 ( 
.A(n_13761),
.B(n_1924),
.Y(n_13947)
);

OR2x2_ASAP7_75t_L g13948 ( 
.A(n_13771),
.B(n_1925),
.Y(n_13948)
);

INVx1_ASAP7_75t_L g13949 ( 
.A(n_13815),
.Y(n_13949)
);

AND2x2_ASAP7_75t_L g13950 ( 
.A(n_13788),
.B(n_1925),
.Y(n_13950)
);

OR2x2_ASAP7_75t_L g13951 ( 
.A(n_13791),
.B(n_1926),
.Y(n_13951)
);

INVx2_ASAP7_75t_SL g13952 ( 
.A(n_13797),
.Y(n_13952)
);

INVx1_ASAP7_75t_L g13953 ( 
.A(n_13829),
.Y(n_13953)
);

INVx2_ASAP7_75t_L g13954 ( 
.A(n_13846),
.Y(n_13954)
);

INVx1_ASAP7_75t_L g13955 ( 
.A(n_13786),
.Y(n_13955)
);

NOR3xp33_ASAP7_75t_L g13956 ( 
.A(n_13838),
.B(n_1926),
.C(n_1927),
.Y(n_13956)
);

INVx1_ASAP7_75t_L g13957 ( 
.A(n_13787),
.Y(n_13957)
);

AND2x2_ASAP7_75t_L g13958 ( 
.A(n_13762),
.B(n_1926),
.Y(n_13958)
);

INVxp67_ASAP7_75t_L g13959 ( 
.A(n_13789),
.Y(n_13959)
);

INVx1_ASAP7_75t_L g13960 ( 
.A(n_13814),
.Y(n_13960)
);

NAND2xp5_ASAP7_75t_L g13961 ( 
.A(n_13759),
.B(n_1927),
.Y(n_13961)
);

INVx1_ASAP7_75t_L g13962 ( 
.A(n_13794),
.Y(n_13962)
);

INVx2_ASAP7_75t_SL g13963 ( 
.A(n_13813),
.Y(n_13963)
);

INVx1_ASAP7_75t_L g13964 ( 
.A(n_13770),
.Y(n_13964)
);

INVx1_ASAP7_75t_L g13965 ( 
.A(n_13776),
.Y(n_13965)
);

INVx1_ASAP7_75t_L g13966 ( 
.A(n_13827),
.Y(n_13966)
);

AND2x2_ASAP7_75t_L g13967 ( 
.A(n_13738),
.B(n_13821),
.Y(n_13967)
);

INVx2_ASAP7_75t_L g13968 ( 
.A(n_13841),
.Y(n_13968)
);

INVx1_ASAP7_75t_SL g13969 ( 
.A(n_13796),
.Y(n_13969)
);

AND2x2_ASAP7_75t_L g13970 ( 
.A(n_13810),
.B(n_1927),
.Y(n_13970)
);

INVx1_ASAP7_75t_L g13971 ( 
.A(n_13807),
.Y(n_13971)
);

INVx1_ASAP7_75t_L g13972 ( 
.A(n_13777),
.Y(n_13972)
);

NOR2x1p5_ASAP7_75t_SL g13973 ( 
.A(n_13778),
.B(n_1928),
.Y(n_13973)
);

HB1xp67_ASAP7_75t_L g13974 ( 
.A(n_13848),
.Y(n_13974)
);

HB1xp67_ASAP7_75t_L g13975 ( 
.A(n_13848),
.Y(n_13975)
);

AND2x2_ASAP7_75t_L g13976 ( 
.A(n_13720),
.B(n_1928),
.Y(n_13976)
);

AOI21xp5_ASAP7_75t_L g13977 ( 
.A1(n_13777),
.A2(n_1928),
.B(n_1929),
.Y(n_13977)
);

INVx2_ASAP7_75t_L g13978 ( 
.A(n_13763),
.Y(n_13978)
);

INVx1_ASAP7_75t_L g13979 ( 
.A(n_13777),
.Y(n_13979)
);

NOR2xp33_ASAP7_75t_L g13980 ( 
.A(n_13767),
.B(n_2411),
.Y(n_13980)
);

NAND2xp5_ASAP7_75t_L g13981 ( 
.A(n_13777),
.B(n_1929),
.Y(n_13981)
);

INVx2_ASAP7_75t_SL g13982 ( 
.A(n_13753),
.Y(n_13982)
);

INVxp67_ASAP7_75t_L g13983 ( 
.A(n_13782),
.Y(n_13983)
);

INVx1_ASAP7_75t_L g13984 ( 
.A(n_13777),
.Y(n_13984)
);

AND2x2_ASAP7_75t_L g13985 ( 
.A(n_13720),
.B(n_1929),
.Y(n_13985)
);

INVx1_ASAP7_75t_L g13986 ( 
.A(n_13777),
.Y(n_13986)
);

INVx1_ASAP7_75t_L g13987 ( 
.A(n_13777),
.Y(n_13987)
);

AND2x2_ASAP7_75t_L g13988 ( 
.A(n_13720),
.B(n_1930),
.Y(n_13988)
);

INVx1_ASAP7_75t_L g13989 ( 
.A(n_13777),
.Y(n_13989)
);

INVx1_ASAP7_75t_L g13990 ( 
.A(n_13777),
.Y(n_13990)
);

OR2x2_ASAP7_75t_L g13991 ( 
.A(n_13747),
.B(n_1930),
.Y(n_13991)
);

INVx1_ASAP7_75t_L g13992 ( 
.A(n_13777),
.Y(n_13992)
);

INVx1_ASAP7_75t_L g13993 ( 
.A(n_13777),
.Y(n_13993)
);

INVx1_ASAP7_75t_L g13994 ( 
.A(n_13777),
.Y(n_13994)
);

INVx2_ASAP7_75t_L g13995 ( 
.A(n_13763),
.Y(n_13995)
);

OR2x2_ASAP7_75t_L g13996 ( 
.A(n_13747),
.B(n_1930),
.Y(n_13996)
);

AND2x4_ASAP7_75t_L g13997 ( 
.A(n_13720),
.B(n_1931),
.Y(n_13997)
);

INVx1_ASAP7_75t_L g13998 ( 
.A(n_13888),
.Y(n_13998)
);

AND2x2_ASAP7_75t_L g13999 ( 
.A(n_13850),
.B(n_13881),
.Y(n_13999)
);

INVx1_ASAP7_75t_L g14000 ( 
.A(n_13973),
.Y(n_14000)
);

AOI22xp5_ASAP7_75t_L g14001 ( 
.A1(n_13900),
.A2(n_1933),
.B1(n_1931),
.B2(n_1932),
.Y(n_14001)
);

NAND2xp5_ASAP7_75t_L g14002 ( 
.A(n_13902),
.B(n_1932),
.Y(n_14002)
);

CKINVDCx16_ASAP7_75t_R g14003 ( 
.A(n_13870),
.Y(n_14003)
);

OR2x2_ASAP7_75t_L g14004 ( 
.A(n_13880),
.B(n_1932),
.Y(n_14004)
);

INVx1_ASAP7_75t_L g14005 ( 
.A(n_13854),
.Y(n_14005)
);

NAND2xp5_ASAP7_75t_L g14006 ( 
.A(n_13892),
.B(n_1933),
.Y(n_14006)
);

NAND2xp5_ASAP7_75t_L g14007 ( 
.A(n_13904),
.B(n_1934),
.Y(n_14007)
);

NAND2xp5_ASAP7_75t_L g14008 ( 
.A(n_13911),
.B(n_1934),
.Y(n_14008)
);

INVx1_ASAP7_75t_SL g14009 ( 
.A(n_13917),
.Y(n_14009)
);

AND2x2_ASAP7_75t_L g14010 ( 
.A(n_13852),
.B(n_1935),
.Y(n_14010)
);

AOI211xp5_ASAP7_75t_SL g14011 ( 
.A1(n_13849),
.A2(n_2421),
.B(n_2423),
.C(n_2420),
.Y(n_14011)
);

NAND2x1_ASAP7_75t_L g14012 ( 
.A(n_13925),
.B(n_1935),
.Y(n_14012)
);

AND2x2_ASAP7_75t_L g14013 ( 
.A(n_13919),
.B(n_1935),
.Y(n_14013)
);

INVx1_ASAP7_75t_L g14014 ( 
.A(n_13974),
.Y(n_14014)
);

OR2x2_ASAP7_75t_L g14015 ( 
.A(n_13963),
.B(n_1936),
.Y(n_14015)
);

INVx1_ASAP7_75t_L g14016 ( 
.A(n_13975),
.Y(n_14016)
);

OR2x2_ASAP7_75t_L g14017 ( 
.A(n_13858),
.B(n_1936),
.Y(n_14017)
);

HB1xp67_ASAP7_75t_L g14018 ( 
.A(n_13924),
.Y(n_14018)
);

AND2x2_ASAP7_75t_L g14019 ( 
.A(n_13972),
.B(n_1936),
.Y(n_14019)
);

INVx1_ASAP7_75t_SL g14020 ( 
.A(n_13863),
.Y(n_14020)
);

NAND2xp5_ASAP7_75t_L g14021 ( 
.A(n_13872),
.B(n_1937),
.Y(n_14021)
);

AND2x2_ASAP7_75t_L g14022 ( 
.A(n_13979),
.B(n_1937),
.Y(n_14022)
);

INVx1_ASAP7_75t_L g14023 ( 
.A(n_13866),
.Y(n_14023)
);

INVx1_ASAP7_75t_L g14024 ( 
.A(n_13936),
.Y(n_14024)
);

OR2x6_ASAP7_75t_L g14025 ( 
.A(n_13907),
.B(n_1938),
.Y(n_14025)
);

OR2x2_ASAP7_75t_L g14026 ( 
.A(n_13984),
.B(n_1939),
.Y(n_14026)
);

AND2x2_ASAP7_75t_SL g14027 ( 
.A(n_13906),
.B(n_1939),
.Y(n_14027)
);

INVx1_ASAP7_75t_L g14028 ( 
.A(n_13877),
.Y(n_14028)
);

INVxp67_ASAP7_75t_L g14029 ( 
.A(n_13876),
.Y(n_14029)
);

INVx2_ASAP7_75t_L g14030 ( 
.A(n_13885),
.Y(n_14030)
);

INVx1_ASAP7_75t_L g14031 ( 
.A(n_13882),
.Y(n_14031)
);

NAND2xp5_ASAP7_75t_L g14032 ( 
.A(n_13997),
.B(n_1940),
.Y(n_14032)
);

INVx1_ASAP7_75t_L g14033 ( 
.A(n_13867),
.Y(n_14033)
);

INVx1_ASAP7_75t_L g14034 ( 
.A(n_13898),
.Y(n_14034)
);

NAND2xp5_ASAP7_75t_L g14035 ( 
.A(n_13946),
.B(n_1940),
.Y(n_14035)
);

INVx1_ASAP7_75t_L g14036 ( 
.A(n_13950),
.Y(n_14036)
);

AOI211x1_ASAP7_75t_L g14037 ( 
.A1(n_13860),
.A2(n_1942),
.B(n_1940),
.C(n_1941),
.Y(n_14037)
);

NAND2xp5_ASAP7_75t_L g14038 ( 
.A(n_13933),
.B(n_1941),
.Y(n_14038)
);

NAND2xp5_ASAP7_75t_SL g14039 ( 
.A(n_13986),
.B(n_1941),
.Y(n_14039)
);

AND2x4_ASAP7_75t_L g14040 ( 
.A(n_13967),
.B(n_1942),
.Y(n_14040)
);

OR2x2_ASAP7_75t_L g14041 ( 
.A(n_13987),
.B(n_1943),
.Y(n_14041)
);

AND2x2_ASAP7_75t_L g14042 ( 
.A(n_13989),
.B(n_1943),
.Y(n_14042)
);

NOR2xp33_ASAP7_75t_L g14043 ( 
.A(n_13908),
.B(n_1943),
.Y(n_14043)
);

INVxp67_ASAP7_75t_L g14044 ( 
.A(n_13932),
.Y(n_14044)
);

AND2x2_ASAP7_75t_L g14045 ( 
.A(n_13990),
.B(n_1944),
.Y(n_14045)
);

AND2x2_ASAP7_75t_L g14046 ( 
.A(n_13992),
.B(n_1944),
.Y(n_14046)
);

INVx2_ASAP7_75t_SL g14047 ( 
.A(n_13991),
.Y(n_14047)
);

INVx2_ASAP7_75t_L g14048 ( 
.A(n_13897),
.Y(n_14048)
);

INVx1_ASAP7_75t_L g14049 ( 
.A(n_13921),
.Y(n_14049)
);

AND2x2_ASAP7_75t_L g14050 ( 
.A(n_13993),
.B(n_1944),
.Y(n_14050)
);

NAND2xp5_ASAP7_75t_L g14051 ( 
.A(n_13939),
.B(n_1945),
.Y(n_14051)
);

OR2x2_ASAP7_75t_L g14052 ( 
.A(n_13994),
.B(n_1945),
.Y(n_14052)
);

AND2x2_ASAP7_75t_L g14053 ( 
.A(n_13857),
.B(n_1945),
.Y(n_14053)
);

AND2x2_ASAP7_75t_L g14054 ( 
.A(n_13853),
.B(n_1946),
.Y(n_14054)
);

OR2x2_ASAP7_75t_L g14055 ( 
.A(n_13891),
.B(n_13996),
.Y(n_14055)
);

AND2x2_ASAP7_75t_L g14056 ( 
.A(n_13884),
.B(n_1946),
.Y(n_14056)
);

INVx2_ASAP7_75t_L g14057 ( 
.A(n_13940),
.Y(n_14057)
);

OR2x2_ASAP7_75t_L g14058 ( 
.A(n_13951),
.B(n_1946),
.Y(n_14058)
);

OR2x2_ASAP7_75t_L g14059 ( 
.A(n_13945),
.B(n_1947),
.Y(n_14059)
);

OR2x2_ASAP7_75t_L g14060 ( 
.A(n_13981),
.B(n_1947),
.Y(n_14060)
);

NAND2xp5_ASAP7_75t_L g14061 ( 
.A(n_13868),
.B(n_1947),
.Y(n_14061)
);

AND2x2_ASAP7_75t_L g14062 ( 
.A(n_13889),
.B(n_1948),
.Y(n_14062)
);

INVx1_ASAP7_75t_L g14063 ( 
.A(n_13976),
.Y(n_14063)
);

INVx1_ASAP7_75t_L g14064 ( 
.A(n_13985),
.Y(n_14064)
);

NAND2xp5_ASAP7_75t_L g14065 ( 
.A(n_13988),
.B(n_13851),
.Y(n_14065)
);

OR2x6_ASAP7_75t_L g14066 ( 
.A(n_13901),
.B(n_1948),
.Y(n_14066)
);

INVx1_ASAP7_75t_L g14067 ( 
.A(n_13914),
.Y(n_14067)
);

AND2x2_ASAP7_75t_L g14068 ( 
.A(n_13968),
.B(n_1948),
.Y(n_14068)
);

INVx1_ASAP7_75t_L g14069 ( 
.A(n_13927),
.Y(n_14069)
);

OR2x2_ASAP7_75t_L g14070 ( 
.A(n_13873),
.B(n_1949),
.Y(n_14070)
);

OR2x2_ASAP7_75t_L g14071 ( 
.A(n_13930),
.B(n_1949),
.Y(n_14071)
);

INVx2_ASAP7_75t_L g14072 ( 
.A(n_13895),
.Y(n_14072)
);

AND2x2_ASAP7_75t_L g14073 ( 
.A(n_13856),
.B(n_1950),
.Y(n_14073)
);

INVx2_ASAP7_75t_L g14074 ( 
.A(n_13978),
.Y(n_14074)
);

INVx1_ASAP7_75t_L g14075 ( 
.A(n_13883),
.Y(n_14075)
);

CKINVDCx16_ASAP7_75t_R g14076 ( 
.A(n_13923),
.Y(n_14076)
);

AND2x2_ASAP7_75t_L g14077 ( 
.A(n_13982),
.B(n_1950),
.Y(n_14077)
);

NOR2xp33_ASAP7_75t_L g14078 ( 
.A(n_13995),
.B(n_1951),
.Y(n_14078)
);

OAI21xp5_ASAP7_75t_L g14079 ( 
.A1(n_13959),
.A2(n_1951),
.B(n_1952),
.Y(n_14079)
);

INVx1_ASAP7_75t_L g14080 ( 
.A(n_13915),
.Y(n_14080)
);

NAND2xp5_ASAP7_75t_L g14081 ( 
.A(n_13855),
.B(n_1951),
.Y(n_14081)
);

INVx1_ASAP7_75t_L g14082 ( 
.A(n_13928),
.Y(n_14082)
);

INVx1_ASAP7_75t_L g14083 ( 
.A(n_13931),
.Y(n_14083)
);

INVx1_ASAP7_75t_L g14084 ( 
.A(n_13935),
.Y(n_14084)
);

AND2x4_ASAP7_75t_SL g14085 ( 
.A(n_13865),
.B(n_1952),
.Y(n_14085)
);

INVxp67_ASAP7_75t_SL g14086 ( 
.A(n_13862),
.Y(n_14086)
);

INVx1_ASAP7_75t_L g14087 ( 
.A(n_13958),
.Y(n_14087)
);

AND2x2_ASAP7_75t_L g14088 ( 
.A(n_13886),
.B(n_1952),
.Y(n_14088)
);

INVx1_ASAP7_75t_L g14089 ( 
.A(n_13869),
.Y(n_14089)
);

INVx1_ASAP7_75t_L g14090 ( 
.A(n_13899),
.Y(n_14090)
);

AND2x2_ASAP7_75t_L g14091 ( 
.A(n_13918),
.B(n_1953),
.Y(n_14091)
);

INVx2_ASAP7_75t_L g14092 ( 
.A(n_13948),
.Y(n_14092)
);

HB1xp67_ASAP7_75t_L g14093 ( 
.A(n_13879),
.Y(n_14093)
);

INVx1_ASAP7_75t_L g14094 ( 
.A(n_13864),
.Y(n_14094)
);

NOR2xp33_ASAP7_75t_L g14095 ( 
.A(n_13937),
.B(n_1954),
.Y(n_14095)
);

AND2x2_ASAP7_75t_L g14096 ( 
.A(n_13955),
.B(n_1954),
.Y(n_14096)
);

INVx1_ASAP7_75t_L g14097 ( 
.A(n_13894),
.Y(n_14097)
);

INVx2_ASAP7_75t_SL g14098 ( 
.A(n_13896),
.Y(n_14098)
);

INVx1_ASAP7_75t_L g14099 ( 
.A(n_13983),
.Y(n_14099)
);

NAND2xp5_ASAP7_75t_L g14100 ( 
.A(n_13922),
.B(n_1954),
.Y(n_14100)
);

AND2x2_ASAP7_75t_L g14101 ( 
.A(n_13957),
.B(n_1955),
.Y(n_14101)
);

NAND3xp33_ASAP7_75t_L g14102 ( 
.A(n_13871),
.B(n_2428),
.C(n_2426),
.Y(n_14102)
);

INVx1_ASAP7_75t_L g14103 ( 
.A(n_13970),
.Y(n_14103)
);

AOI22xp5_ASAP7_75t_L g14104 ( 
.A1(n_13910),
.A2(n_1957),
.B1(n_1955),
.B2(n_1956),
.Y(n_14104)
);

CKINVDCx8_ASAP7_75t_R g14105 ( 
.A(n_13980),
.Y(n_14105)
);

INVx1_ASAP7_75t_L g14106 ( 
.A(n_13878),
.Y(n_14106)
);

NAND2xp5_ASAP7_75t_L g14107 ( 
.A(n_13934),
.B(n_13938),
.Y(n_14107)
);

INVx1_ASAP7_75t_L g14108 ( 
.A(n_13943),
.Y(n_14108)
);

INVx1_ASAP7_75t_L g14109 ( 
.A(n_13912),
.Y(n_14109)
);

INVx1_ASAP7_75t_L g14110 ( 
.A(n_13942),
.Y(n_14110)
);

OR2x2_ASAP7_75t_L g14111 ( 
.A(n_13953),
.B(n_1956),
.Y(n_14111)
);

AND2x2_ASAP7_75t_L g14112 ( 
.A(n_13929),
.B(n_1957),
.Y(n_14112)
);

INVxp67_ASAP7_75t_SL g14113 ( 
.A(n_13861),
.Y(n_14113)
);

OR2x2_ASAP7_75t_L g14114 ( 
.A(n_13875),
.B(n_1958),
.Y(n_14114)
);

OR2x2_ASAP7_75t_L g14115 ( 
.A(n_13874),
.B(n_1958),
.Y(n_14115)
);

NAND2xp5_ASAP7_75t_L g14116 ( 
.A(n_13969),
.B(n_1959),
.Y(n_14116)
);

OR2x2_ASAP7_75t_L g14117 ( 
.A(n_13859),
.B(n_1959),
.Y(n_14117)
);

AND2x2_ASAP7_75t_L g14118 ( 
.A(n_13890),
.B(n_1959),
.Y(n_14118)
);

OR2x2_ASAP7_75t_L g14119 ( 
.A(n_13961),
.B(n_1960),
.Y(n_14119)
);

NAND2xp5_ASAP7_75t_L g14120 ( 
.A(n_13949),
.B(n_1960),
.Y(n_14120)
);

NOR2xp33_ASAP7_75t_L g14121 ( 
.A(n_13893),
.B(n_1961),
.Y(n_14121)
);

NAND2xp5_ASAP7_75t_L g14122 ( 
.A(n_13952),
.B(n_1961),
.Y(n_14122)
);

AND2x2_ASAP7_75t_L g14123 ( 
.A(n_13903),
.B(n_1961),
.Y(n_14123)
);

AOI22xp33_ASAP7_75t_L g14124 ( 
.A1(n_13913),
.A2(n_1964),
.B1(n_1962),
.B2(n_1963),
.Y(n_14124)
);

INVx1_ASAP7_75t_L g14125 ( 
.A(n_13944),
.Y(n_14125)
);

NAND2xp5_ASAP7_75t_L g14126 ( 
.A(n_13977),
.B(n_1962),
.Y(n_14126)
);

NAND2xp5_ASAP7_75t_L g14127 ( 
.A(n_13926),
.B(n_1963),
.Y(n_14127)
);

INVx1_ASAP7_75t_L g14128 ( 
.A(n_13920),
.Y(n_14128)
);

INVx1_ASAP7_75t_L g14129 ( 
.A(n_13916),
.Y(n_14129)
);

INVx1_ASAP7_75t_L g14130 ( 
.A(n_13999),
.Y(n_14130)
);

NAND4xp25_ASAP7_75t_L g14131 ( 
.A(n_14009),
.B(n_13941),
.C(n_13965),
.D(n_13954),
.Y(n_14131)
);

OAI22xp5_ASAP7_75t_L g14132 ( 
.A1(n_14003),
.A2(n_13909),
.B1(n_13887),
.B2(n_13905),
.Y(n_14132)
);

INVx2_ASAP7_75t_L g14133 ( 
.A(n_14027),
.Y(n_14133)
);

AOI22xp33_ASAP7_75t_L g14134 ( 
.A1(n_14000),
.A2(n_13971),
.B1(n_13966),
.B2(n_13962),
.Y(n_14134)
);

OAI21xp5_ASAP7_75t_SL g14135 ( 
.A1(n_14018),
.A2(n_13947),
.B(n_13964),
.Y(n_14135)
);

NAND2xp5_ASAP7_75t_L g14136 ( 
.A(n_13998),
.B(n_13956),
.Y(n_14136)
);

NOR2xp33_ASAP7_75t_L g14137 ( 
.A(n_14024),
.B(n_13960),
.Y(n_14137)
);

INVx1_ASAP7_75t_L g14138 ( 
.A(n_14093),
.Y(n_14138)
);

NOR2xp33_ASAP7_75t_L g14139 ( 
.A(n_14020),
.B(n_1963),
.Y(n_14139)
);

INVx1_ASAP7_75t_L g14140 ( 
.A(n_14066),
.Y(n_14140)
);

AOI22xp5_ASAP7_75t_L g14141 ( 
.A1(n_14099),
.A2(n_1966),
.B1(n_1964),
.B2(n_1965),
.Y(n_14141)
);

NAND2xp5_ASAP7_75t_L g14142 ( 
.A(n_14011),
.B(n_2416),
.Y(n_14142)
);

AOI21xp33_ASAP7_75t_SL g14143 ( 
.A1(n_14076),
.A2(n_2421),
.B(n_2420),
.Y(n_14143)
);

INVx1_ASAP7_75t_L g14144 ( 
.A(n_14066),
.Y(n_14144)
);

OA21x2_ASAP7_75t_L g14145 ( 
.A1(n_14102),
.A2(n_1964),
.B(n_1966),
.Y(n_14145)
);

AOI22xp33_ASAP7_75t_L g14146 ( 
.A1(n_14072),
.A2(n_1968),
.B1(n_1969),
.B2(n_1967),
.Y(n_14146)
);

AOI22xp5_ASAP7_75t_L g14147 ( 
.A1(n_14029),
.A2(n_1968),
.B1(n_1966),
.B2(n_1967),
.Y(n_14147)
);

AOI21xp5_ASAP7_75t_L g14148 ( 
.A1(n_14039),
.A2(n_1970),
.B(n_1969),
.Y(n_14148)
);

NAND2xp5_ASAP7_75t_SL g14149 ( 
.A(n_14040),
.B(n_1967),
.Y(n_14149)
);

INVx2_ASAP7_75t_L g14150 ( 
.A(n_14012),
.Y(n_14150)
);

BUFx2_ASAP7_75t_L g14151 ( 
.A(n_14088),
.Y(n_14151)
);

HB1xp67_ASAP7_75t_L g14152 ( 
.A(n_14025),
.Y(n_14152)
);

OAI322xp33_ASAP7_75t_L g14153 ( 
.A1(n_14005),
.A2(n_1975),
.A3(n_1974),
.B1(n_1972),
.B2(n_1970),
.C1(n_1971),
.C2(n_1973),
.Y(n_14153)
);

AND2x4_ASAP7_75t_L g14154 ( 
.A(n_14034),
.B(n_1971),
.Y(n_14154)
);

INVx1_ASAP7_75t_SL g14155 ( 
.A(n_14053),
.Y(n_14155)
);

INVx2_ASAP7_75t_SL g14156 ( 
.A(n_14017),
.Y(n_14156)
);

AOI221xp5_ASAP7_75t_L g14157 ( 
.A1(n_14014),
.A2(n_1973),
.B1(n_1971),
.B2(n_1972),
.C(n_1974),
.Y(n_14157)
);

INVx2_ASAP7_75t_L g14158 ( 
.A(n_14055),
.Y(n_14158)
);

INVx2_ASAP7_75t_L g14159 ( 
.A(n_14056),
.Y(n_14159)
);

NAND4xp25_ASAP7_75t_L g14160 ( 
.A(n_14107),
.B(n_1975),
.C(n_1972),
.D(n_1974),
.Y(n_14160)
);

AND2x4_ASAP7_75t_L g14161 ( 
.A(n_14073),
.B(n_1975),
.Y(n_14161)
);

INVx1_ASAP7_75t_SL g14162 ( 
.A(n_14054),
.Y(n_14162)
);

INVx1_ASAP7_75t_L g14163 ( 
.A(n_14062),
.Y(n_14163)
);

INVx2_ASAP7_75t_L g14164 ( 
.A(n_14010),
.Y(n_14164)
);

OAI32xp33_ASAP7_75t_L g14165 ( 
.A1(n_14015),
.A2(n_14044),
.A3(n_14051),
.B1(n_14109),
.B2(n_14125),
.Y(n_14165)
);

INVx1_ASAP7_75t_L g14166 ( 
.A(n_14085),
.Y(n_14166)
);

INVx1_ASAP7_75t_SL g14167 ( 
.A(n_14013),
.Y(n_14167)
);

AND2x2_ASAP7_75t_L g14168 ( 
.A(n_14077),
.B(n_1976),
.Y(n_14168)
);

OR2x2_ASAP7_75t_L g14169 ( 
.A(n_14026),
.B(n_1976),
.Y(n_14169)
);

INVx2_ASAP7_75t_L g14170 ( 
.A(n_14058),
.Y(n_14170)
);

NOR2xp33_ASAP7_75t_L g14171 ( 
.A(n_14033),
.B(n_1976),
.Y(n_14171)
);

INVx1_ASAP7_75t_L g14172 ( 
.A(n_14025),
.Y(n_14172)
);

AOI22xp5_ASAP7_75t_L g14173 ( 
.A1(n_14047),
.A2(n_1979),
.B1(n_1977),
.B2(n_1978),
.Y(n_14173)
);

INVx1_ASAP7_75t_L g14174 ( 
.A(n_14037),
.Y(n_14174)
);

NAND2x1p5_ASAP7_75t_L g14175 ( 
.A(n_14030),
.B(n_1977),
.Y(n_14175)
);

INVx1_ASAP7_75t_L g14176 ( 
.A(n_14071),
.Y(n_14176)
);

NAND2xp5_ASAP7_75t_L g14177 ( 
.A(n_14098),
.B(n_2412),
.Y(n_14177)
);

INVx1_ASAP7_75t_L g14178 ( 
.A(n_14091),
.Y(n_14178)
);

INVx2_ASAP7_75t_L g14179 ( 
.A(n_14004),
.Y(n_14179)
);

NOR2xp67_ASAP7_75t_L g14180 ( 
.A(n_14110),
.B(n_1978),
.Y(n_14180)
);

AND2x4_ASAP7_75t_L g14181 ( 
.A(n_14129),
.B(n_1978),
.Y(n_14181)
);

INVx1_ASAP7_75t_L g14182 ( 
.A(n_14007),
.Y(n_14182)
);

OAI21xp5_ASAP7_75t_SL g14183 ( 
.A1(n_14016),
.A2(n_14118),
.B(n_14122),
.Y(n_14183)
);

INVx1_ASAP7_75t_L g14184 ( 
.A(n_14006),
.Y(n_14184)
);

INVxp33_ASAP7_75t_L g14185 ( 
.A(n_14043),
.Y(n_14185)
);

NAND2xp5_ASAP7_75t_L g14186 ( 
.A(n_14028),
.B(n_2413),
.Y(n_14186)
);

INVx1_ASAP7_75t_L g14187 ( 
.A(n_14008),
.Y(n_14187)
);

INVx2_ASAP7_75t_L g14188 ( 
.A(n_14048),
.Y(n_14188)
);

INVx1_ASAP7_75t_SL g14189 ( 
.A(n_14068),
.Y(n_14189)
);

INVx2_ASAP7_75t_L g14190 ( 
.A(n_14023),
.Y(n_14190)
);

NAND2xp5_ASAP7_75t_L g14191 ( 
.A(n_14031),
.B(n_2414),
.Y(n_14191)
);

AND2x2_ASAP7_75t_L g14192 ( 
.A(n_14019),
.B(n_1979),
.Y(n_14192)
);

NOR2xp33_ASAP7_75t_L g14193 ( 
.A(n_14105),
.B(n_1979),
.Y(n_14193)
);

INVx1_ASAP7_75t_L g14194 ( 
.A(n_14021),
.Y(n_14194)
);

AO21x1_ASAP7_75t_L g14195 ( 
.A1(n_14095),
.A2(n_2423),
.B(n_2420),
.Y(n_14195)
);

NAND2x1p5_ASAP7_75t_L g14196 ( 
.A(n_14036),
.B(n_1980),
.Y(n_14196)
);

AOI21xp33_ASAP7_75t_L g14197 ( 
.A1(n_14086),
.A2(n_2424),
.B(n_2423),
.Y(n_14197)
);

OR2x2_ASAP7_75t_L g14198 ( 
.A(n_14041),
.B(n_1980),
.Y(n_14198)
);

INVx2_ASAP7_75t_L g14199 ( 
.A(n_14111),
.Y(n_14199)
);

AOI21xp5_ASAP7_75t_L g14200 ( 
.A1(n_14002),
.A2(n_1982),
.B(n_1981),
.Y(n_14200)
);

INVx1_ASAP7_75t_L g14201 ( 
.A(n_14022),
.Y(n_14201)
);

INVx2_ASAP7_75t_L g14202 ( 
.A(n_14052),
.Y(n_14202)
);

O2A1O1Ixp33_ASAP7_75t_SL g14203 ( 
.A1(n_14035),
.A2(n_1982),
.B(n_1980),
.C(n_1981),
.Y(n_14203)
);

INVx1_ASAP7_75t_L g14204 ( 
.A(n_14042),
.Y(n_14204)
);

INVx1_ASAP7_75t_L g14205 ( 
.A(n_14045),
.Y(n_14205)
);

INVx1_ASAP7_75t_SL g14206 ( 
.A(n_14046),
.Y(n_14206)
);

HB1xp67_ASAP7_75t_L g14207 ( 
.A(n_14050),
.Y(n_14207)
);

AOI22xp5_ASAP7_75t_L g14208 ( 
.A1(n_14075),
.A2(n_1984),
.B1(n_1981),
.B2(n_1983),
.Y(n_14208)
);

INVx1_ASAP7_75t_L g14209 ( 
.A(n_14096),
.Y(n_14209)
);

NAND2xp5_ASAP7_75t_L g14210 ( 
.A(n_14123),
.B(n_2443),
.Y(n_14210)
);

AND2x2_ASAP7_75t_L g14211 ( 
.A(n_14074),
.B(n_1983),
.Y(n_14211)
);

AND2x2_ASAP7_75t_L g14212 ( 
.A(n_14101),
.B(n_1984),
.Y(n_14212)
);

OA21x2_ASAP7_75t_L g14213 ( 
.A1(n_14079),
.A2(n_14100),
.B(n_14081),
.Y(n_14213)
);

NAND2xp5_ASAP7_75t_L g14214 ( 
.A(n_14067),
.B(n_2402),
.Y(n_14214)
);

NAND2xp33_ASAP7_75t_L g14215 ( 
.A(n_14112),
.B(n_1985),
.Y(n_14215)
);

OR2x2_ASAP7_75t_L g14216 ( 
.A(n_14061),
.B(n_1985),
.Y(n_14216)
);

AOI32xp33_ASAP7_75t_L g14217 ( 
.A1(n_14089),
.A2(n_1987),
.A3(n_1985),
.B1(n_1986),
.B2(n_1988),
.Y(n_14217)
);

INVx1_ASAP7_75t_L g14218 ( 
.A(n_14057),
.Y(n_14218)
);

INVx1_ASAP7_75t_L g14219 ( 
.A(n_14032),
.Y(n_14219)
);

INVx1_ASAP7_75t_L g14220 ( 
.A(n_14038),
.Y(n_14220)
);

AND2x2_ASAP7_75t_L g14221 ( 
.A(n_14084),
.B(n_1986),
.Y(n_14221)
);

OAI22xp5_ASAP7_75t_L g14222 ( 
.A1(n_14001),
.A2(n_14124),
.B1(n_14104),
.B2(n_14121),
.Y(n_14222)
);

OAI22xp33_ASAP7_75t_L g14223 ( 
.A1(n_14126),
.A2(n_1988),
.B1(n_1986),
.B2(n_1987),
.Y(n_14223)
);

OAI22xp33_ASAP7_75t_SL g14224 ( 
.A1(n_14113),
.A2(n_1989),
.B1(n_1987),
.B2(n_1988),
.Y(n_14224)
);

OAI221xp5_ASAP7_75t_L g14225 ( 
.A1(n_14065),
.A2(n_1991),
.B1(n_1989),
.B2(n_1990),
.C(n_1992),
.Y(n_14225)
);

INVx1_ASAP7_75t_L g14226 ( 
.A(n_14049),
.Y(n_14226)
);

AND2x4_ASAP7_75t_L g14227 ( 
.A(n_14087),
.B(n_1989),
.Y(n_14227)
);

AND2x2_ASAP7_75t_L g14228 ( 
.A(n_14069),
.B(n_1990),
.Y(n_14228)
);

INVx1_ASAP7_75t_L g14229 ( 
.A(n_14059),
.Y(n_14229)
);

AND2x2_ASAP7_75t_L g14230 ( 
.A(n_14078),
.B(n_1990),
.Y(n_14230)
);

AOI22xp33_ASAP7_75t_L g14231 ( 
.A1(n_14108),
.A2(n_1993),
.B1(n_1994),
.B2(n_1992),
.Y(n_14231)
);

INVx1_ASAP7_75t_L g14232 ( 
.A(n_14092),
.Y(n_14232)
);

AND2x4_ASAP7_75t_L g14233 ( 
.A(n_14063),
.B(n_1991),
.Y(n_14233)
);

INVxp33_ASAP7_75t_L g14234 ( 
.A(n_14116),
.Y(n_14234)
);

INVx2_ASAP7_75t_L g14235 ( 
.A(n_14115),
.Y(n_14235)
);

AND2x4_ASAP7_75t_L g14236 ( 
.A(n_14064),
.B(n_1991),
.Y(n_14236)
);

NOR2xp33_ASAP7_75t_L g14237 ( 
.A(n_14117),
.B(n_1992),
.Y(n_14237)
);

INVx3_ASAP7_75t_L g14238 ( 
.A(n_14070),
.Y(n_14238)
);

AND2x2_ASAP7_75t_L g14239 ( 
.A(n_14128),
.B(n_1993),
.Y(n_14239)
);

INVx1_ASAP7_75t_L g14240 ( 
.A(n_14060),
.Y(n_14240)
);

NAND2xp5_ASAP7_75t_L g14241 ( 
.A(n_14080),
.B(n_2412),
.Y(n_14241)
);

OAI21xp5_ASAP7_75t_L g14242 ( 
.A1(n_14120),
.A2(n_1994),
.B(n_1995),
.Y(n_14242)
);

A2O1A1Ixp33_ASAP7_75t_L g14243 ( 
.A1(n_14106),
.A2(n_1997),
.B(n_1995),
.C(n_1996),
.Y(n_14243)
);

INVxp67_ASAP7_75t_L g14244 ( 
.A(n_14103),
.Y(n_14244)
);

AOI21xp33_ASAP7_75t_L g14245 ( 
.A1(n_14097),
.A2(n_2431),
.B(n_2429),
.Y(n_14245)
);

INVx2_ASAP7_75t_L g14246 ( 
.A(n_14119),
.Y(n_14246)
);

A2O1A1Ixp33_ASAP7_75t_L g14247 ( 
.A1(n_14135),
.A2(n_14114),
.B(n_14127),
.C(n_14094),
.Y(n_14247)
);

INVx2_ASAP7_75t_L g14248 ( 
.A(n_14175),
.Y(n_14248)
);

OAI21xp5_ASAP7_75t_L g14249 ( 
.A1(n_14138),
.A2(n_14083),
.B(n_14082),
.Y(n_14249)
);

AOI21xp5_ASAP7_75t_L g14250 ( 
.A1(n_14137),
.A2(n_14090),
.B(n_1996),
.Y(n_14250)
);

INVx2_ASAP7_75t_SL g14251 ( 
.A(n_14196),
.Y(n_14251)
);

INVx1_ASAP7_75t_L g14252 ( 
.A(n_14151),
.Y(n_14252)
);

INVx2_ASAP7_75t_L g14253 ( 
.A(n_14161),
.Y(n_14253)
);

AOI221xp5_ASAP7_75t_L g14254 ( 
.A1(n_14165),
.A2(n_1998),
.B1(n_1996),
.B2(n_1997),
.C(n_1999),
.Y(n_14254)
);

AOI22xp5_ASAP7_75t_L g14255 ( 
.A1(n_14133),
.A2(n_1999),
.B1(n_1997),
.B2(n_1998),
.Y(n_14255)
);

NOR2x1_ASAP7_75t_L g14256 ( 
.A(n_14131),
.B(n_1998),
.Y(n_14256)
);

NAND2x1p5_ASAP7_75t_L g14257 ( 
.A(n_14158),
.B(n_2000),
.Y(n_14257)
);

INVx2_ASAP7_75t_L g14258 ( 
.A(n_14192),
.Y(n_14258)
);

OAI22xp33_ASAP7_75t_SL g14259 ( 
.A1(n_14150),
.A2(n_2007),
.B1(n_2015),
.B2(n_1999),
.Y(n_14259)
);

AND2x4_ASAP7_75t_L g14260 ( 
.A(n_14130),
.B(n_2000),
.Y(n_14260)
);

INVx1_ASAP7_75t_L g14261 ( 
.A(n_14195),
.Y(n_14261)
);

INVx1_ASAP7_75t_L g14262 ( 
.A(n_14152),
.Y(n_14262)
);

INVx1_ASAP7_75t_L g14263 ( 
.A(n_14207),
.Y(n_14263)
);

INVx1_ASAP7_75t_L g14264 ( 
.A(n_14180),
.Y(n_14264)
);

NAND2xp5_ASAP7_75t_L g14265 ( 
.A(n_14206),
.B(n_2401),
.Y(n_14265)
);

AOI21x1_ASAP7_75t_L g14266 ( 
.A1(n_14226),
.A2(n_14181),
.B(n_14218),
.Y(n_14266)
);

O2A1O1Ixp33_ASAP7_75t_L g14267 ( 
.A1(n_14244),
.A2(n_2002),
.B(n_2000),
.C(n_2001),
.Y(n_14267)
);

OAI22xp5_ASAP7_75t_L g14268 ( 
.A1(n_14134),
.A2(n_2003),
.B1(n_2001),
.B2(n_2002),
.Y(n_14268)
);

NOR2xp33_ASAP7_75t_L g14269 ( 
.A(n_14143),
.B(n_2403),
.Y(n_14269)
);

AOI322xp5_ASAP7_75t_L g14270 ( 
.A1(n_14167),
.A2(n_2007),
.A3(n_2006),
.B1(n_2004),
.B2(n_2001),
.C1(n_2003),
.C2(n_2005),
.Y(n_14270)
);

OAI22xp5_ASAP7_75t_L g14271 ( 
.A1(n_14190),
.A2(n_2005),
.B1(n_2003),
.B2(n_2004),
.Y(n_14271)
);

AOI22xp5_ASAP7_75t_L g14272 ( 
.A1(n_14132),
.A2(n_2008),
.B1(n_2004),
.B2(n_2006),
.Y(n_14272)
);

AOI21xp33_ASAP7_75t_SL g14273 ( 
.A1(n_14166),
.A2(n_2411),
.B(n_2410),
.Y(n_14273)
);

INVx1_ASAP7_75t_L g14274 ( 
.A(n_14168),
.Y(n_14274)
);

INVx2_ASAP7_75t_SL g14275 ( 
.A(n_14154),
.Y(n_14275)
);

NAND2xp5_ASAP7_75t_L g14276 ( 
.A(n_14212),
.B(n_2410),
.Y(n_14276)
);

NAND2xp5_ASAP7_75t_L g14277 ( 
.A(n_14156),
.B(n_2411),
.Y(n_14277)
);

INVx2_ASAP7_75t_SL g14278 ( 
.A(n_14227),
.Y(n_14278)
);

O2A1O1Ixp33_ASAP7_75t_L g14279 ( 
.A1(n_14224),
.A2(n_2010),
.B(n_2008),
.C(n_2009),
.Y(n_14279)
);

INVx1_ASAP7_75t_L g14280 ( 
.A(n_14142),
.Y(n_14280)
);

AND2x2_ASAP7_75t_L g14281 ( 
.A(n_14232),
.B(n_2009),
.Y(n_14281)
);

OAI21xp33_ASAP7_75t_L g14282 ( 
.A1(n_14139),
.A2(n_2011),
.B(n_2012),
.Y(n_14282)
);

NOR3xp33_ASAP7_75t_L g14283 ( 
.A(n_14183),
.B(n_2399),
.C(n_2398),
.Y(n_14283)
);

INVx1_ASAP7_75t_L g14284 ( 
.A(n_14174),
.Y(n_14284)
);

HB1xp67_ASAP7_75t_L g14285 ( 
.A(n_14145),
.Y(n_14285)
);

AOI21xp33_ASAP7_75t_L g14286 ( 
.A1(n_14234),
.A2(n_2398),
.B(n_2397),
.Y(n_14286)
);

NAND2xp5_ASAP7_75t_L g14287 ( 
.A(n_14188),
.B(n_2397),
.Y(n_14287)
);

AOI22xp33_ASAP7_75t_SL g14288 ( 
.A1(n_14136),
.A2(n_2014),
.B1(n_2012),
.B2(n_2013),
.Y(n_14288)
);

OAI21xp33_ASAP7_75t_L g14289 ( 
.A1(n_14193),
.A2(n_2012),
.B(n_2014),
.Y(n_14289)
);

NAND2xp5_ASAP7_75t_L g14290 ( 
.A(n_14211),
.B(n_2401),
.Y(n_14290)
);

INVx1_ASAP7_75t_L g14291 ( 
.A(n_14203),
.Y(n_14291)
);

INVx1_ASAP7_75t_L g14292 ( 
.A(n_14169),
.Y(n_14292)
);

INVx1_ASAP7_75t_L g14293 ( 
.A(n_14198),
.Y(n_14293)
);

INVx1_ASAP7_75t_L g14294 ( 
.A(n_14215),
.Y(n_14294)
);

AND2x2_ASAP7_75t_L g14295 ( 
.A(n_14233),
.B(n_2015),
.Y(n_14295)
);

NOR4xp25_ASAP7_75t_L g14296 ( 
.A(n_14162),
.B(n_2019),
.C(n_2016),
.D(n_2017),
.Y(n_14296)
);

OAI21xp33_ASAP7_75t_L g14297 ( 
.A1(n_14171),
.A2(n_2016),
.B(n_2017),
.Y(n_14297)
);

INVx1_ASAP7_75t_L g14298 ( 
.A(n_14221),
.Y(n_14298)
);

AOI22xp33_ASAP7_75t_L g14299 ( 
.A1(n_14202),
.A2(n_2019),
.B1(n_2016),
.B2(n_2017),
.Y(n_14299)
);

NAND2xp5_ASAP7_75t_L g14300 ( 
.A(n_14236),
.B(n_2405),
.Y(n_14300)
);

OAI21xp5_ASAP7_75t_L g14301 ( 
.A1(n_14148),
.A2(n_2019),
.B(n_2020),
.Y(n_14301)
);

AND2x2_ASAP7_75t_L g14302 ( 
.A(n_14228),
.B(n_2020),
.Y(n_14302)
);

NOR2xp33_ASAP7_75t_L g14303 ( 
.A(n_14153),
.B(n_2407),
.Y(n_14303)
);

OAI31xp33_ASAP7_75t_L g14304 ( 
.A1(n_14222),
.A2(n_2022),
.A3(n_2020),
.B(n_2021),
.Y(n_14304)
);

INVx1_ASAP7_75t_L g14305 ( 
.A(n_14164),
.Y(n_14305)
);

NAND2xp5_ASAP7_75t_L g14306 ( 
.A(n_14230),
.B(n_2408),
.Y(n_14306)
);

AND2x2_ASAP7_75t_L g14307 ( 
.A(n_14239),
.B(n_14213),
.Y(n_14307)
);

OAI22xp5_ASAP7_75t_L g14308 ( 
.A1(n_14173),
.A2(n_2023),
.B1(n_2021),
.B2(n_2022),
.Y(n_14308)
);

NOR2xp33_ASAP7_75t_L g14309 ( 
.A(n_14160),
.B(n_2419),
.Y(n_14309)
);

INVx1_ASAP7_75t_L g14310 ( 
.A(n_14159),
.Y(n_14310)
);

OAI21xp33_ASAP7_75t_L g14311 ( 
.A1(n_14177),
.A2(n_2021),
.B(n_2023),
.Y(n_14311)
);

AOI21xp33_ASAP7_75t_SL g14312 ( 
.A1(n_14149),
.A2(n_2443),
.B(n_2023),
.Y(n_14312)
);

INVx1_ASAP7_75t_L g14313 ( 
.A(n_14163),
.Y(n_14313)
);

INVx2_ASAP7_75t_L g14314 ( 
.A(n_14213),
.Y(n_14314)
);

OA21x2_ASAP7_75t_L g14315 ( 
.A1(n_14186),
.A2(n_2024),
.B(n_2025),
.Y(n_14315)
);

INVx1_ASAP7_75t_L g14316 ( 
.A(n_14179),
.Y(n_14316)
);

AOI22xp5_ASAP7_75t_L g14317 ( 
.A1(n_14155),
.A2(n_2026),
.B1(n_2024),
.B2(n_2025),
.Y(n_14317)
);

OAI32xp33_ASAP7_75t_L g14318 ( 
.A1(n_14191),
.A2(n_2028),
.A3(n_2026),
.B1(n_2027),
.B2(n_2029),
.Y(n_14318)
);

INVx1_ASAP7_75t_L g14319 ( 
.A(n_14170),
.Y(n_14319)
);

NAND2xp5_ASAP7_75t_L g14320 ( 
.A(n_14201),
.B(n_2396),
.Y(n_14320)
);

INVx1_ASAP7_75t_L g14321 ( 
.A(n_14145),
.Y(n_14321)
);

OAI322xp33_ASAP7_75t_L g14322 ( 
.A1(n_14204),
.A2(n_2033),
.A3(n_2032),
.B1(n_2030),
.B2(n_2027),
.C1(n_2028),
.C2(n_2031),
.Y(n_14322)
);

NAND2xp33_ASAP7_75t_L g14323 ( 
.A(n_14217),
.B(n_2030),
.Y(n_14323)
);

INVx2_ASAP7_75t_L g14324 ( 
.A(n_14238),
.Y(n_14324)
);

INVxp67_ASAP7_75t_L g14325 ( 
.A(n_14237),
.Y(n_14325)
);

INVx2_ASAP7_75t_L g14326 ( 
.A(n_14199),
.Y(n_14326)
);

AOI22xp5_ASAP7_75t_L g14327 ( 
.A1(n_14205),
.A2(n_2032),
.B1(n_2027),
.B2(n_2031),
.Y(n_14327)
);

AND2x2_ASAP7_75t_L g14328 ( 
.A(n_14208),
.B(n_14209),
.Y(n_14328)
);

NAND2xp5_ASAP7_75t_L g14329 ( 
.A(n_14189),
.B(n_2402),
.Y(n_14329)
);

INVx1_ASAP7_75t_L g14330 ( 
.A(n_14210),
.Y(n_14330)
);

NOR3xp33_ASAP7_75t_L g14331 ( 
.A(n_14172),
.B(n_2404),
.C(n_2403),
.Y(n_14331)
);

INVx1_ASAP7_75t_L g14332 ( 
.A(n_14176),
.Y(n_14332)
);

NAND2xp5_ASAP7_75t_L g14333 ( 
.A(n_14178),
.B(n_2402),
.Y(n_14333)
);

AOI22xp33_ASAP7_75t_L g14334 ( 
.A1(n_14182),
.A2(n_2034),
.B1(n_2031),
.B2(n_2032),
.Y(n_14334)
);

AOI21xp33_ASAP7_75t_SL g14335 ( 
.A1(n_14197),
.A2(n_2408),
.B(n_2407),
.Y(n_14335)
);

AND2x2_ASAP7_75t_L g14336 ( 
.A(n_14231),
.B(n_2034),
.Y(n_14336)
);

NAND2xp5_ASAP7_75t_SL g14337 ( 
.A(n_14157),
.B(n_2036),
.Y(n_14337)
);

INVx2_ASAP7_75t_SL g14338 ( 
.A(n_14216),
.Y(n_14338)
);

AND2x2_ASAP7_75t_L g14339 ( 
.A(n_14146),
.B(n_2035),
.Y(n_14339)
);

INVx2_ASAP7_75t_L g14340 ( 
.A(n_14246),
.Y(n_14340)
);

INVxp67_ASAP7_75t_L g14341 ( 
.A(n_14140),
.Y(n_14341)
);

OR2x2_ASAP7_75t_L g14342 ( 
.A(n_14214),
.B(n_2035),
.Y(n_14342)
);

NAND2xp5_ASAP7_75t_L g14343 ( 
.A(n_14200),
.B(n_2408),
.Y(n_14343)
);

OAI22xp5_ASAP7_75t_L g14344 ( 
.A1(n_14147),
.A2(n_2037),
.B1(n_2035),
.B2(n_2036),
.Y(n_14344)
);

NAND2xp5_ASAP7_75t_L g14345 ( 
.A(n_14184),
.B(n_2443),
.Y(n_14345)
);

NOR2xp33_ASAP7_75t_L g14346 ( 
.A(n_14185),
.B(n_2036),
.Y(n_14346)
);

AOI22xp5_ASAP7_75t_L g14347 ( 
.A1(n_14219),
.A2(n_2039),
.B1(n_2037),
.B2(n_2038),
.Y(n_14347)
);

INVx1_ASAP7_75t_L g14348 ( 
.A(n_14144),
.Y(n_14348)
);

INVx1_ASAP7_75t_L g14349 ( 
.A(n_14235),
.Y(n_14349)
);

OR2x2_ASAP7_75t_L g14350 ( 
.A(n_14241),
.B(n_2038),
.Y(n_14350)
);

NAND2x2_ASAP7_75t_L g14351 ( 
.A(n_14223),
.B(n_2038),
.Y(n_14351)
);

NAND4xp25_ASAP7_75t_L g14352 ( 
.A(n_14242),
.B(n_2041),
.C(n_2039),
.D(n_2040),
.Y(n_14352)
);

AOI21xp5_ASAP7_75t_L g14353 ( 
.A1(n_14252),
.A2(n_14225),
.B(n_14243),
.Y(n_14353)
);

AND2x2_ASAP7_75t_L g14354 ( 
.A(n_14324),
.B(n_14141),
.Y(n_14354)
);

OR2x2_ASAP7_75t_L g14355 ( 
.A(n_14314),
.B(n_14187),
.Y(n_14355)
);

OAI21xp5_ASAP7_75t_L g14356 ( 
.A1(n_14263),
.A2(n_14245),
.B(n_14220),
.Y(n_14356)
);

NAND2xp5_ASAP7_75t_L g14357 ( 
.A(n_14296),
.B(n_14194),
.Y(n_14357)
);

AOI22xp5_ASAP7_75t_L g14358 ( 
.A1(n_14251),
.A2(n_14229),
.B1(n_14240),
.B2(n_2041),
.Y(n_14358)
);

AND2x2_ASAP7_75t_L g14359 ( 
.A(n_14266),
.B(n_2039),
.Y(n_14359)
);

INVx1_ASAP7_75t_SL g14360 ( 
.A(n_14281),
.Y(n_14360)
);

NAND2xp5_ASAP7_75t_L g14361 ( 
.A(n_14291),
.B(n_2040),
.Y(n_14361)
);

AND2x2_ASAP7_75t_L g14362 ( 
.A(n_14313),
.B(n_14249),
.Y(n_14362)
);

AOI222xp33_ASAP7_75t_L g14363 ( 
.A1(n_14321),
.A2(n_2044),
.B1(n_2046),
.B2(n_2042),
.C1(n_2043),
.C2(n_2045),
.Y(n_14363)
);

OAI21xp33_ASAP7_75t_L g14364 ( 
.A1(n_14305),
.A2(n_2051),
.B(n_2043),
.Y(n_14364)
);

AND2x2_ASAP7_75t_L g14365 ( 
.A(n_14310),
.B(n_2043),
.Y(n_14365)
);

AOI322xp5_ASAP7_75t_L g14366 ( 
.A1(n_14256),
.A2(n_2049),
.A3(n_2048),
.B1(n_2046),
.B2(n_2044),
.C1(n_2045),
.C2(n_2047),
.Y(n_14366)
);

AOI22xp33_ASAP7_75t_L g14367 ( 
.A1(n_14280),
.A2(n_2047),
.B1(n_2045),
.B2(n_2046),
.Y(n_14367)
);

NOR2xp33_ASAP7_75t_L g14368 ( 
.A(n_14261),
.B(n_2047),
.Y(n_14368)
);

INVx1_ASAP7_75t_L g14369 ( 
.A(n_14307),
.Y(n_14369)
);

NOR2x1_ASAP7_75t_L g14370 ( 
.A(n_14260),
.B(n_2048),
.Y(n_14370)
);

NAND3xp33_ASAP7_75t_L g14371 ( 
.A(n_14285),
.B(n_2049),
.C(n_2050),
.Y(n_14371)
);

AOI22xp5_ASAP7_75t_SL g14372 ( 
.A1(n_14259),
.A2(n_2052),
.B1(n_2050),
.B2(n_2051),
.Y(n_14372)
);

OAI22xp5_ASAP7_75t_L g14373 ( 
.A1(n_14317),
.A2(n_2052),
.B1(n_2050),
.B2(n_2051),
.Y(n_14373)
);

NAND2xp5_ASAP7_75t_L g14374 ( 
.A(n_14302),
.B(n_2052),
.Y(n_14374)
);

INVx2_ASAP7_75t_L g14375 ( 
.A(n_14257),
.Y(n_14375)
);

NAND2xp5_ASAP7_75t_SL g14376 ( 
.A(n_14273),
.B(n_2053),
.Y(n_14376)
);

NAND4xp25_ASAP7_75t_L g14377 ( 
.A(n_14349),
.B(n_2055),
.C(n_2053),
.D(n_2054),
.Y(n_14377)
);

NAND4xp25_ASAP7_75t_L g14378 ( 
.A(n_14316),
.B(n_2057),
.C(n_2054),
.D(n_2056),
.Y(n_14378)
);

NOR2xp33_ASAP7_75t_L g14379 ( 
.A(n_14248),
.B(n_2056),
.Y(n_14379)
);

XNOR2x1_ASAP7_75t_L g14380 ( 
.A(n_14258),
.B(n_2056),
.Y(n_14380)
);

INVxp67_ASAP7_75t_SL g14381 ( 
.A(n_14276),
.Y(n_14381)
);

INVx1_ASAP7_75t_L g14382 ( 
.A(n_14315),
.Y(n_14382)
);

AOI21xp33_ASAP7_75t_L g14383 ( 
.A1(n_14264),
.A2(n_2057),
.B(n_2058),
.Y(n_14383)
);

INVx1_ASAP7_75t_L g14384 ( 
.A(n_14315),
.Y(n_14384)
);

OR2x2_ASAP7_75t_L g14385 ( 
.A(n_14278),
.B(n_2057),
.Y(n_14385)
);

INVx2_ASAP7_75t_L g14386 ( 
.A(n_14295),
.Y(n_14386)
);

INVx1_ASAP7_75t_L g14387 ( 
.A(n_14326),
.Y(n_14387)
);

INVx2_ASAP7_75t_SL g14388 ( 
.A(n_14275),
.Y(n_14388)
);

AOI22xp33_ASAP7_75t_L g14389 ( 
.A1(n_14338),
.A2(n_2060),
.B1(n_2058),
.B2(n_2059),
.Y(n_14389)
);

INVx1_ASAP7_75t_L g14390 ( 
.A(n_14340),
.Y(n_14390)
);

AOI22xp5_ASAP7_75t_L g14391 ( 
.A1(n_14284),
.A2(n_14332),
.B1(n_14303),
.B2(n_14269),
.Y(n_14391)
);

AOI21xp33_ASAP7_75t_L g14392 ( 
.A1(n_14262),
.A2(n_2059),
.B(n_2060),
.Y(n_14392)
);

AO21x1_ASAP7_75t_L g14393 ( 
.A1(n_14268),
.A2(n_2060),
.B(n_2061),
.Y(n_14393)
);

AOI222xp33_ASAP7_75t_L g14394 ( 
.A1(n_14341),
.A2(n_2063),
.B1(n_2065),
.B2(n_2061),
.C1(n_2062),
.C2(n_2064),
.Y(n_14394)
);

NAND2x1p5_ASAP7_75t_L g14395 ( 
.A(n_14319),
.B(n_2061),
.Y(n_14395)
);

A2O1A1Ixp33_ASAP7_75t_L g14396 ( 
.A1(n_14250),
.A2(n_2064),
.B(n_2062),
.C(n_2063),
.Y(n_14396)
);

AOI21xp5_ASAP7_75t_L g14397 ( 
.A1(n_14300),
.A2(n_2062),
.B(n_2063),
.Y(n_14397)
);

INVx1_ASAP7_75t_L g14398 ( 
.A(n_14274),
.Y(n_14398)
);

INVx2_ASAP7_75t_SL g14399 ( 
.A(n_14351),
.Y(n_14399)
);

AOI32xp33_ASAP7_75t_L g14400 ( 
.A1(n_14323),
.A2(n_2067),
.A3(n_2064),
.B1(n_2066),
.B2(n_2068),
.Y(n_14400)
);

OAI32xp33_ASAP7_75t_L g14401 ( 
.A1(n_14283),
.A2(n_14287),
.A3(n_14277),
.B1(n_14265),
.B2(n_14329),
.Y(n_14401)
);

INVx1_ASAP7_75t_L g14402 ( 
.A(n_14306),
.Y(n_14402)
);

AND2x2_ASAP7_75t_L g14403 ( 
.A(n_14309),
.B(n_2066),
.Y(n_14403)
);

AOI22xp5_ASAP7_75t_L g14404 ( 
.A1(n_14298),
.A2(n_2069),
.B1(n_2067),
.B2(n_2068),
.Y(n_14404)
);

INVxp33_ASAP7_75t_L g14405 ( 
.A(n_14346),
.Y(n_14405)
);

NAND2xp5_ASAP7_75t_L g14406 ( 
.A(n_14312),
.B(n_2067),
.Y(n_14406)
);

AND2x2_ASAP7_75t_L g14407 ( 
.A(n_14301),
.B(n_2068),
.Y(n_14407)
);

OAI322xp33_ASAP7_75t_L g14408 ( 
.A1(n_14337),
.A2(n_2074),
.A3(n_2073),
.B1(n_2071),
.B2(n_2069),
.C1(n_2070),
.C2(n_2072),
.Y(n_14408)
);

OAI21xp5_ASAP7_75t_L g14409 ( 
.A1(n_14247),
.A2(n_2069),
.B(n_2070),
.Y(n_14409)
);

A2O1A1Ixp33_ASAP7_75t_L g14410 ( 
.A1(n_14267),
.A2(n_2072),
.B(n_2070),
.C(n_2071),
.Y(n_14410)
);

INVx1_ASAP7_75t_L g14411 ( 
.A(n_14292),
.Y(n_14411)
);

AOI21xp33_ASAP7_75t_L g14412 ( 
.A1(n_14279),
.A2(n_2071),
.B(n_2073),
.Y(n_14412)
);

INVx2_ASAP7_75t_L g14413 ( 
.A(n_14253),
.Y(n_14413)
);

AOI221xp5_ASAP7_75t_L g14414 ( 
.A1(n_14335),
.A2(n_2075),
.B1(n_2073),
.B2(n_2074),
.C(n_2076),
.Y(n_14414)
);

OAI22xp5_ASAP7_75t_L g14415 ( 
.A1(n_14272),
.A2(n_2076),
.B1(n_2074),
.B2(n_2075),
.Y(n_14415)
);

NAND2xp33_ASAP7_75t_L g14416 ( 
.A(n_14331),
.B(n_2077),
.Y(n_14416)
);

INVx1_ASAP7_75t_L g14417 ( 
.A(n_14293),
.Y(n_14417)
);

INVx1_ASAP7_75t_L g14418 ( 
.A(n_14290),
.Y(n_14418)
);

INVxp67_ASAP7_75t_L g14419 ( 
.A(n_14294),
.Y(n_14419)
);

AO22x1_ASAP7_75t_L g14420 ( 
.A1(n_14271),
.A2(n_14328),
.B1(n_14333),
.B2(n_14320),
.Y(n_14420)
);

OAI321xp33_ASAP7_75t_L g14421 ( 
.A1(n_14348),
.A2(n_2079),
.A3(n_2081),
.B1(n_2077),
.B2(n_2078),
.C(n_2080),
.Y(n_14421)
);

NOR2xp33_ASAP7_75t_L g14422 ( 
.A(n_14322),
.B(n_2077),
.Y(n_14422)
);

OAI322xp33_ASAP7_75t_L g14423 ( 
.A1(n_14325),
.A2(n_14330),
.A3(n_14345),
.B1(n_14343),
.B2(n_14350),
.C1(n_14342),
.C2(n_14255),
.Y(n_14423)
);

OAI332xp33_ASAP7_75t_L g14424 ( 
.A1(n_14308),
.A2(n_2399),
.A3(n_2083),
.B1(n_2080),
.B2(n_2084),
.B3(n_2082),
.C1(n_2078),
.C2(n_2079),
.Y(n_14424)
);

AOI322xp5_ASAP7_75t_L g14425 ( 
.A1(n_14336),
.A2(n_14339),
.A3(n_14282),
.B1(n_14297),
.B2(n_14311),
.C1(n_14289),
.C2(n_14286),
.Y(n_14425)
);

OAI22xp33_ASAP7_75t_SL g14426 ( 
.A1(n_14344),
.A2(n_2080),
.B1(n_2078),
.B2(n_2079),
.Y(n_14426)
);

INVx3_ASAP7_75t_L g14427 ( 
.A(n_14318),
.Y(n_14427)
);

AOI322xp5_ASAP7_75t_L g14428 ( 
.A1(n_14254),
.A2(n_14299),
.A3(n_14334),
.B1(n_14288),
.B2(n_14327),
.C1(n_14347),
.C2(n_14352),
.Y(n_14428)
);

AND2x2_ASAP7_75t_L g14429 ( 
.A(n_14270),
.B(n_2081),
.Y(n_14429)
);

NOR5xp2_ASAP7_75t_L g14430 ( 
.A(n_14304),
.B(n_2083),
.C(n_2081),
.D(n_2082),
.E(n_2084),
.Y(n_14430)
);

NOR2xp33_ASAP7_75t_L g14431 ( 
.A(n_14291),
.B(n_2428),
.Y(n_14431)
);

INVx1_ASAP7_75t_L g14432 ( 
.A(n_14307),
.Y(n_14432)
);

AOI21xp5_ASAP7_75t_L g14433 ( 
.A1(n_14252),
.A2(n_2428),
.B(n_2083),
.Y(n_14433)
);

AOI22xp33_ASAP7_75t_L g14434 ( 
.A1(n_14314),
.A2(n_2407),
.B1(n_2087),
.B2(n_2085),
.Y(n_14434)
);

INVx1_ASAP7_75t_L g14435 ( 
.A(n_14307),
.Y(n_14435)
);

NAND4xp25_ASAP7_75t_L g14436 ( 
.A(n_14252),
.B(n_2087),
.C(n_2085),
.D(n_2086),
.Y(n_14436)
);

AOI211xp5_ASAP7_75t_L g14437 ( 
.A1(n_14252),
.A2(n_2089),
.B(n_2086),
.C(n_2088),
.Y(n_14437)
);

NAND2xp5_ASAP7_75t_L g14438 ( 
.A(n_14314),
.B(n_2088),
.Y(n_14438)
);

AOI21xp5_ASAP7_75t_L g14439 ( 
.A1(n_14252),
.A2(n_2406),
.B(n_2088),
.Y(n_14439)
);

OAI31xp33_ASAP7_75t_L g14440 ( 
.A1(n_14369),
.A2(n_14435),
.A3(n_14432),
.B(n_14359),
.Y(n_14440)
);

OAI21xp33_ASAP7_75t_L g14441 ( 
.A1(n_14387),
.A2(n_2089),
.B(n_2090),
.Y(n_14441)
);

INVx1_ASAP7_75t_L g14442 ( 
.A(n_14382),
.Y(n_14442)
);

AOI222xp33_ASAP7_75t_L g14443 ( 
.A1(n_14384),
.A2(n_2091),
.B1(n_2093),
.B2(n_2089),
.C1(n_2090),
.C2(n_2092),
.Y(n_14443)
);

AOI221xp5_ASAP7_75t_L g14444 ( 
.A1(n_14390),
.A2(n_2092),
.B1(n_2090),
.B2(n_2091),
.C(n_2093),
.Y(n_14444)
);

A2O1A1Ixp33_ASAP7_75t_L g14445 ( 
.A1(n_14355),
.A2(n_2094),
.B(n_2091),
.C(n_2093),
.Y(n_14445)
);

NAND4xp25_ASAP7_75t_SL g14446 ( 
.A(n_14362),
.B(n_2096),
.C(n_2094),
.D(n_2095),
.Y(n_14446)
);

AOI211xp5_ASAP7_75t_L g14447 ( 
.A1(n_14431),
.A2(n_14419),
.B(n_14438),
.C(n_14368),
.Y(n_14447)
);

NAND2xp5_ASAP7_75t_L g14448 ( 
.A(n_14370),
.B(n_2094),
.Y(n_14448)
);

OAI22xp33_ASAP7_75t_L g14449 ( 
.A1(n_14361),
.A2(n_2097),
.B1(n_2095),
.B2(n_2096),
.Y(n_14449)
);

OAI22xp33_ASAP7_75t_L g14450 ( 
.A1(n_14358),
.A2(n_2097),
.B1(n_2095),
.B2(n_2096),
.Y(n_14450)
);

INVx2_ASAP7_75t_L g14451 ( 
.A(n_14395),
.Y(n_14451)
);

AOI221xp5_ASAP7_75t_L g14452 ( 
.A1(n_14398),
.A2(n_2099),
.B1(n_2097),
.B2(n_2098),
.C(n_2100),
.Y(n_14452)
);

INVx2_ASAP7_75t_L g14453 ( 
.A(n_14375),
.Y(n_14453)
);

INVx1_ASAP7_75t_L g14454 ( 
.A(n_14357),
.Y(n_14454)
);

NAND2xp5_ASAP7_75t_L g14455 ( 
.A(n_14360),
.B(n_2098),
.Y(n_14455)
);

AND2x2_ASAP7_75t_L g14456 ( 
.A(n_14388),
.B(n_2098),
.Y(n_14456)
);

AOI22xp5_ASAP7_75t_L g14457 ( 
.A1(n_14399),
.A2(n_2101),
.B1(n_2099),
.B2(n_2100),
.Y(n_14457)
);

INVx2_ASAP7_75t_SL g14458 ( 
.A(n_14385),
.Y(n_14458)
);

NAND2xp5_ASAP7_75t_L g14459 ( 
.A(n_14372),
.B(n_2100),
.Y(n_14459)
);

AND2x2_ASAP7_75t_L g14460 ( 
.A(n_14354),
.B(n_2101),
.Y(n_14460)
);

NAND3xp33_ASAP7_75t_L g14461 ( 
.A(n_14366),
.B(n_2102),
.C(n_2103),
.Y(n_14461)
);

AOI22xp33_ASAP7_75t_L g14462 ( 
.A1(n_14386),
.A2(n_2104),
.B1(n_2102),
.B2(n_2103),
.Y(n_14462)
);

OAI21xp5_ASAP7_75t_SL g14463 ( 
.A1(n_14391),
.A2(n_2102),
.B(n_2104),
.Y(n_14463)
);

O2A1O1Ixp33_ASAP7_75t_L g14464 ( 
.A1(n_14356),
.A2(n_2406),
.B(n_2106),
.C(n_2104),
.Y(n_14464)
);

INVx1_ASAP7_75t_L g14465 ( 
.A(n_14365),
.Y(n_14465)
);

AOI22xp5_ASAP7_75t_L g14466 ( 
.A1(n_14411),
.A2(n_2107),
.B1(n_2105),
.B2(n_2106),
.Y(n_14466)
);

OAI222xp33_ASAP7_75t_L g14467 ( 
.A1(n_14400),
.A2(n_2107),
.B1(n_2109),
.B2(n_2105),
.C1(n_2106),
.C2(n_2108),
.Y(n_14467)
);

O2A1O1Ixp33_ASAP7_75t_L g14468 ( 
.A1(n_14396),
.A2(n_2404),
.B(n_2109),
.C(n_2105),
.Y(n_14468)
);

OAI22xp33_ASAP7_75t_L g14469 ( 
.A1(n_14404),
.A2(n_2111),
.B1(n_2108),
.B2(n_2110),
.Y(n_14469)
);

INVx1_ASAP7_75t_L g14470 ( 
.A(n_14413),
.Y(n_14470)
);

AOI22xp33_ASAP7_75t_SL g14471 ( 
.A1(n_14417),
.A2(n_2111),
.B1(n_2108),
.B2(n_2110),
.Y(n_14471)
);

AOI22xp5_ASAP7_75t_L g14472 ( 
.A1(n_14429),
.A2(n_2113),
.B1(n_2110),
.B2(n_2112),
.Y(n_14472)
);

OAI22xp5_ASAP7_75t_L g14473 ( 
.A1(n_14434),
.A2(n_2114),
.B1(n_2112),
.B2(n_2113),
.Y(n_14473)
);

NAND2xp5_ASAP7_75t_L g14474 ( 
.A(n_14420),
.B(n_2112),
.Y(n_14474)
);

OAI22xp5_ASAP7_75t_L g14475 ( 
.A1(n_14389),
.A2(n_2116),
.B1(n_2114),
.B2(n_2115),
.Y(n_14475)
);

OR2x2_ASAP7_75t_L g14476 ( 
.A(n_14436),
.B(n_2114),
.Y(n_14476)
);

AOI222xp33_ASAP7_75t_L g14477 ( 
.A1(n_14416),
.A2(n_2117),
.B1(n_2119),
.B2(n_2115),
.C1(n_2116),
.C2(n_2118),
.Y(n_14477)
);

AOI21xp5_ASAP7_75t_L g14478 ( 
.A1(n_14353),
.A2(n_2115),
.B(n_2116),
.Y(n_14478)
);

INVx1_ASAP7_75t_L g14479 ( 
.A(n_14374),
.Y(n_14479)
);

INVx1_ASAP7_75t_L g14480 ( 
.A(n_14393),
.Y(n_14480)
);

AND2x2_ASAP7_75t_L g14481 ( 
.A(n_14409),
.B(n_14403),
.Y(n_14481)
);

OAI21xp5_ASAP7_75t_SL g14482 ( 
.A1(n_14422),
.A2(n_14371),
.B(n_14363),
.Y(n_14482)
);

INVxp67_ASAP7_75t_L g14483 ( 
.A(n_14376),
.Y(n_14483)
);

O2A1O1Ixp33_ASAP7_75t_SL g14484 ( 
.A1(n_14410),
.A2(n_2119),
.B(n_2117),
.C(n_2118),
.Y(n_14484)
);

AOI222xp33_ASAP7_75t_L g14485 ( 
.A1(n_14381),
.A2(n_2119),
.B1(n_2121),
.B2(n_2117),
.C1(n_2118),
.C2(n_2120),
.Y(n_14485)
);

AOI22xp5_ASAP7_75t_L g14486 ( 
.A1(n_14407),
.A2(n_2122),
.B1(n_2120),
.B2(n_2121),
.Y(n_14486)
);

AOI22xp33_ASAP7_75t_L g14487 ( 
.A1(n_14405),
.A2(n_2122),
.B1(n_2120),
.B2(n_2121),
.Y(n_14487)
);

INVx2_ASAP7_75t_L g14488 ( 
.A(n_14380),
.Y(n_14488)
);

NAND2xp5_ASAP7_75t_SL g14489 ( 
.A(n_14421),
.B(n_2123),
.Y(n_14489)
);

A2O1A1Ixp33_ASAP7_75t_L g14490 ( 
.A1(n_14364),
.A2(n_2125),
.B(n_2123),
.C(n_2124),
.Y(n_14490)
);

AOI222xp33_ASAP7_75t_L g14491 ( 
.A1(n_14427),
.A2(n_2126),
.B1(n_2128),
.B2(n_2124),
.C1(n_2125),
.C2(n_2127),
.Y(n_14491)
);

OAI21xp5_ASAP7_75t_L g14492 ( 
.A1(n_14433),
.A2(n_2124),
.B(n_2125),
.Y(n_14492)
);

INVx1_ASAP7_75t_L g14493 ( 
.A(n_14427),
.Y(n_14493)
);

OAI221xp5_ASAP7_75t_L g14494 ( 
.A1(n_14437),
.A2(n_2128),
.B1(n_2126),
.B2(n_2127),
.C(n_2129),
.Y(n_14494)
);

OAI221xp5_ASAP7_75t_L g14495 ( 
.A1(n_14377),
.A2(n_2129),
.B1(n_2126),
.B2(n_2128),
.C(n_2130),
.Y(n_14495)
);

AOI221xp5_ASAP7_75t_L g14496 ( 
.A1(n_14401),
.A2(n_2132),
.B1(n_2130),
.B2(n_2131),
.C(n_2133),
.Y(n_14496)
);

INVx1_ASAP7_75t_L g14497 ( 
.A(n_14406),
.Y(n_14497)
);

INVx1_ASAP7_75t_L g14498 ( 
.A(n_14379),
.Y(n_14498)
);

NAND2xp5_ASAP7_75t_L g14499 ( 
.A(n_14402),
.B(n_2130),
.Y(n_14499)
);

AOI211xp5_ASAP7_75t_L g14500 ( 
.A1(n_14373),
.A2(n_2133),
.B(n_2131),
.C(n_2132),
.Y(n_14500)
);

AOI22xp5_ASAP7_75t_L g14501 ( 
.A1(n_14415),
.A2(n_2135),
.B1(n_2131),
.B2(n_2134),
.Y(n_14501)
);

AOI221xp5_ASAP7_75t_L g14502 ( 
.A1(n_14412),
.A2(n_2136),
.B1(n_2134),
.B2(n_2135),
.C(n_2137),
.Y(n_14502)
);

INVx1_ASAP7_75t_L g14503 ( 
.A(n_14378),
.Y(n_14503)
);

NAND2xp5_ASAP7_75t_L g14504 ( 
.A(n_14418),
.B(n_2136),
.Y(n_14504)
);

AOI211xp5_ASAP7_75t_L g14505 ( 
.A1(n_14408),
.A2(n_2139),
.B(n_2137),
.C(n_2138),
.Y(n_14505)
);

NAND2xp5_ASAP7_75t_SL g14506 ( 
.A(n_14493),
.B(n_14394),
.Y(n_14506)
);

AOI32xp33_ASAP7_75t_L g14507 ( 
.A1(n_14454),
.A2(n_14414),
.A3(n_14367),
.B1(n_14428),
.B2(n_14430),
.Y(n_14507)
);

AOI32xp33_ASAP7_75t_L g14508 ( 
.A1(n_14442),
.A2(n_14470),
.A3(n_14503),
.B1(n_14480),
.B2(n_14453),
.Y(n_14508)
);

AND2x2_ASAP7_75t_L g14509 ( 
.A(n_14456),
.B(n_14383),
.Y(n_14509)
);

OAI21xp33_ASAP7_75t_L g14510 ( 
.A1(n_14482),
.A2(n_14463),
.B(n_14455),
.Y(n_14510)
);

O2A1O1Ixp5_ASAP7_75t_L g14511 ( 
.A1(n_14474),
.A2(n_14489),
.B(n_14451),
.C(n_14478),
.Y(n_14511)
);

AND2x2_ASAP7_75t_L g14512 ( 
.A(n_14460),
.B(n_14392),
.Y(n_14512)
);

OAI21xp5_ASAP7_75t_SL g14513 ( 
.A1(n_14440),
.A2(n_14439),
.B(n_14397),
.Y(n_14513)
);

O2A1O1Ixp33_ASAP7_75t_L g14514 ( 
.A1(n_14445),
.A2(n_14423),
.B(n_14426),
.C(n_14424),
.Y(n_14514)
);

OAI211xp5_ASAP7_75t_SL g14515 ( 
.A1(n_14447),
.A2(n_14425),
.B(n_2140),
.C(n_2138),
.Y(n_14515)
);

NAND2xp5_ASAP7_75t_SL g14516 ( 
.A(n_14471),
.B(n_2138),
.Y(n_14516)
);

OAI321xp33_ASAP7_75t_L g14517 ( 
.A1(n_14483),
.A2(n_14461),
.A3(n_14458),
.B1(n_14472),
.B2(n_14488),
.C(n_14465),
.Y(n_14517)
);

AOI221x1_ASAP7_75t_L g14518 ( 
.A1(n_14441),
.A2(n_2141),
.B1(n_2139),
.B2(n_2140),
.C(n_2142),
.Y(n_14518)
);

NAND2xp5_ASAP7_75t_L g14519 ( 
.A(n_14481),
.B(n_2139),
.Y(n_14519)
);

AOI211xp5_ASAP7_75t_SL g14520 ( 
.A1(n_14450),
.A2(n_2142),
.B(n_2140),
.C(n_2141),
.Y(n_14520)
);

AOI221x1_ASAP7_75t_L g14521 ( 
.A1(n_14459),
.A2(n_14499),
.B1(n_14504),
.B2(n_14490),
.C(n_14473),
.Y(n_14521)
);

NAND2xp5_ASAP7_75t_L g14522 ( 
.A(n_14448),
.B(n_2142),
.Y(n_14522)
);

AOI322xp5_ASAP7_75t_L g14523 ( 
.A1(n_14497),
.A2(n_2404),
.A3(n_2148),
.B1(n_2145),
.B2(n_2147),
.C1(n_2143),
.C2(n_2144),
.Y(n_14523)
);

OAI21xp33_ASAP7_75t_L g14524 ( 
.A1(n_14446),
.A2(n_2143),
.B(n_2144),
.Y(n_14524)
);

AOI221xp5_ASAP7_75t_L g14525 ( 
.A1(n_14464),
.A2(n_2146),
.B1(n_2143),
.B2(n_2145),
.C(n_2147),
.Y(n_14525)
);

OAI21xp5_ASAP7_75t_SL g14526 ( 
.A1(n_14491),
.A2(n_14467),
.B(n_14477),
.Y(n_14526)
);

NOR2xp33_ASAP7_75t_L g14527 ( 
.A(n_14476),
.B(n_2145),
.Y(n_14527)
);

AOI21xp5_ASAP7_75t_L g14528 ( 
.A1(n_14484),
.A2(n_2147),
.B(n_2149),
.Y(n_14528)
);

AOI21xp5_ASAP7_75t_L g14529 ( 
.A1(n_14496),
.A2(n_2149),
.B(n_2150),
.Y(n_14529)
);

NAND2xp5_ASAP7_75t_L g14530 ( 
.A(n_14479),
.B(n_2150),
.Y(n_14530)
);

AOI221xp5_ASAP7_75t_L g14531 ( 
.A1(n_14495),
.A2(n_14494),
.B1(n_14469),
.B2(n_14475),
.C(n_14502),
.Y(n_14531)
);

AOI222xp33_ASAP7_75t_L g14532 ( 
.A1(n_14498),
.A2(n_2152),
.B1(n_2154),
.B2(n_2150),
.C1(n_2151),
.C2(n_2153),
.Y(n_14532)
);

AOI211xp5_ASAP7_75t_L g14533 ( 
.A1(n_14449),
.A2(n_2153),
.B(n_2151),
.C(n_2152),
.Y(n_14533)
);

NAND2xp5_ASAP7_75t_L g14534 ( 
.A(n_14505),
.B(n_14443),
.Y(n_14534)
);

INVx2_ASAP7_75t_L g14535 ( 
.A(n_14486),
.Y(n_14535)
);

AOI211xp5_ASAP7_75t_L g14536 ( 
.A1(n_14492),
.A2(n_2153),
.B(n_2151),
.C(n_2152),
.Y(n_14536)
);

NAND2xp5_ASAP7_75t_L g14537 ( 
.A(n_14485),
.B(n_2154),
.Y(n_14537)
);

AOI211xp5_ASAP7_75t_L g14538 ( 
.A1(n_14444),
.A2(n_14452),
.B(n_14468),
.C(n_14500),
.Y(n_14538)
);

AOI21xp5_ASAP7_75t_L g14539 ( 
.A1(n_14462),
.A2(n_2154),
.B(n_2155),
.Y(n_14539)
);

AOI322xp5_ASAP7_75t_L g14540 ( 
.A1(n_14501),
.A2(n_14487),
.A3(n_14466),
.B1(n_14457),
.B2(n_2157),
.C1(n_2160),
.C2(n_2159),
.Y(n_14540)
);

OAI21xp5_ASAP7_75t_SL g14541 ( 
.A1(n_14440),
.A2(n_2155),
.B(n_2156),
.Y(n_14541)
);

AOI21xp5_ASAP7_75t_L g14542 ( 
.A1(n_14440),
.A2(n_2155),
.B(n_2156),
.Y(n_14542)
);

AOI221x1_ASAP7_75t_L g14543 ( 
.A1(n_14442),
.A2(n_2159),
.B1(n_2157),
.B2(n_2158),
.C(n_2160),
.Y(n_14543)
);

AOI211xp5_ASAP7_75t_L g14544 ( 
.A1(n_14454),
.A2(n_2159),
.B(n_2157),
.C(n_2158),
.Y(n_14544)
);

AND2x2_ASAP7_75t_L g14545 ( 
.A(n_14493),
.B(n_2161),
.Y(n_14545)
);

INVx1_ASAP7_75t_L g14546 ( 
.A(n_14460),
.Y(n_14546)
);

NAND2xp5_ASAP7_75t_L g14547 ( 
.A(n_14442),
.B(n_2161),
.Y(n_14547)
);

AOI21xp5_ASAP7_75t_SL g14548 ( 
.A1(n_14454),
.A2(n_2162),
.B(n_2163),
.Y(n_14548)
);

AOI22xp5_ASAP7_75t_L g14549 ( 
.A1(n_14454),
.A2(n_2164),
.B1(n_2162),
.B2(n_2163),
.Y(n_14549)
);

AOI222xp33_ASAP7_75t_L g14550 ( 
.A1(n_14506),
.A2(n_2165),
.B1(n_2167),
.B2(n_2162),
.C1(n_2164),
.C2(n_2166),
.Y(n_14550)
);

AOI221xp5_ASAP7_75t_L g14551 ( 
.A1(n_14508),
.A2(n_2167),
.B1(n_2165),
.B2(n_2166),
.C(n_2168),
.Y(n_14551)
);

OAI21xp5_ASAP7_75t_L g14552 ( 
.A1(n_14511),
.A2(n_2165),
.B(n_2166),
.Y(n_14552)
);

OAI21xp33_ASAP7_75t_L g14553 ( 
.A1(n_14510),
.A2(n_2167),
.B(n_2168),
.Y(n_14553)
);

NAND4xp25_ASAP7_75t_L g14554 ( 
.A(n_14514),
.B(n_2172),
.C(n_2169),
.D(n_2171),
.Y(n_14554)
);

O2A1O1Ixp33_ASAP7_75t_L g14555 ( 
.A1(n_14541),
.A2(n_2173),
.B(n_2169),
.C(n_2171),
.Y(n_14555)
);

OAI211xp5_ASAP7_75t_SL g14556 ( 
.A1(n_14507),
.A2(n_2174),
.B(n_2171),
.C(n_2173),
.Y(n_14556)
);

AOI21xp5_ASAP7_75t_L g14557 ( 
.A1(n_14547),
.A2(n_2174),
.B(n_2175),
.Y(n_14557)
);

AOI21xp33_ASAP7_75t_L g14558 ( 
.A1(n_14546),
.A2(n_2174),
.B(n_2176),
.Y(n_14558)
);

AOI211xp5_ASAP7_75t_SL g14559 ( 
.A1(n_14517),
.A2(n_2178),
.B(n_2176),
.C(n_2177),
.Y(n_14559)
);

AOI21xp5_ASAP7_75t_L g14560 ( 
.A1(n_14548),
.A2(n_14519),
.B(n_14537),
.Y(n_14560)
);

OAI211xp5_ASAP7_75t_L g14561 ( 
.A1(n_14513),
.A2(n_2400),
.B(n_2179),
.C(n_2177),
.Y(n_14561)
);

NAND3xp33_ASAP7_75t_L g14562 ( 
.A(n_14542),
.B(n_2178),
.C(n_2179),
.Y(n_14562)
);

AOI22xp5_ASAP7_75t_L g14563 ( 
.A1(n_14515),
.A2(n_2182),
.B1(n_2180),
.B2(n_2181),
.Y(n_14563)
);

INVx1_ASAP7_75t_L g14564 ( 
.A(n_14545),
.Y(n_14564)
);

NOR3xp33_ASAP7_75t_L g14565 ( 
.A(n_14530),
.B(n_2180),
.C(n_2181),
.Y(n_14565)
);

OAI21xp5_ASAP7_75t_L g14566 ( 
.A1(n_14528),
.A2(n_2180),
.B(n_2181),
.Y(n_14566)
);

AOI322xp5_ASAP7_75t_L g14567 ( 
.A1(n_14527),
.A2(n_2187),
.A3(n_2186),
.B1(n_2184),
.B2(n_2182),
.C1(n_2183),
.C2(n_2185),
.Y(n_14567)
);

INVx1_ASAP7_75t_L g14568 ( 
.A(n_14543),
.Y(n_14568)
);

AOI21xp5_ASAP7_75t_L g14569 ( 
.A1(n_14522),
.A2(n_14516),
.B(n_14526),
.Y(n_14569)
);

NAND2xp5_ASAP7_75t_L g14570 ( 
.A(n_14512),
.B(n_2182),
.Y(n_14570)
);

AOI21xp5_ASAP7_75t_L g14571 ( 
.A1(n_14524),
.A2(n_2184),
.B(n_2185),
.Y(n_14571)
);

NAND2xp5_ASAP7_75t_L g14572 ( 
.A(n_14509),
.B(n_2184),
.Y(n_14572)
);

AOI211xp5_ASAP7_75t_L g14573 ( 
.A1(n_14525),
.A2(n_2187),
.B(n_2185),
.C(n_2186),
.Y(n_14573)
);

OAI221xp5_ASAP7_75t_L g14574 ( 
.A1(n_14544),
.A2(n_2188),
.B1(n_2186),
.B2(n_2187),
.C(n_2189),
.Y(n_14574)
);

NOR2xp33_ASAP7_75t_L g14575 ( 
.A(n_14534),
.B(n_2188),
.Y(n_14575)
);

AOI22xp5_ASAP7_75t_L g14576 ( 
.A1(n_14549),
.A2(n_2190),
.B1(n_2188),
.B2(n_2189),
.Y(n_14576)
);

AND2x2_ASAP7_75t_L g14577 ( 
.A(n_14520),
.B(n_2189),
.Y(n_14577)
);

OAI21xp33_ASAP7_75t_SL g14578 ( 
.A1(n_14540),
.A2(n_2191),
.B(n_2192),
.Y(n_14578)
);

AOI22xp5_ASAP7_75t_L g14579 ( 
.A1(n_14531),
.A2(n_2194),
.B1(n_2191),
.B2(n_2193),
.Y(n_14579)
);

NAND4xp75_ASAP7_75t_L g14580 ( 
.A(n_14521),
.B(n_2194),
.C(n_2191),
.D(n_2193),
.Y(n_14580)
);

AND2x2_ASAP7_75t_L g14581 ( 
.A(n_14577),
.B(n_14536),
.Y(n_14581)
);

NAND2xp5_ASAP7_75t_L g14582 ( 
.A(n_14568),
.B(n_14535),
.Y(n_14582)
);

NAND4xp25_ASAP7_75t_L g14583 ( 
.A(n_14559),
.B(n_14533),
.C(n_14518),
.D(n_14538),
.Y(n_14583)
);

NOR2x1_ASAP7_75t_L g14584 ( 
.A(n_14572),
.B(n_14529),
.Y(n_14584)
);

INVx1_ASAP7_75t_L g14585 ( 
.A(n_14580),
.Y(n_14585)
);

HB1xp67_ASAP7_75t_L g14586 ( 
.A(n_14564),
.Y(n_14586)
);

NOR2x1_ASAP7_75t_L g14587 ( 
.A(n_14570),
.B(n_14539),
.Y(n_14587)
);

NAND2xp5_ASAP7_75t_L g14588 ( 
.A(n_14560),
.B(n_14532),
.Y(n_14588)
);

NAND2xp5_ASAP7_75t_L g14589 ( 
.A(n_14569),
.B(n_14523),
.Y(n_14589)
);

AOI21xp33_ASAP7_75t_L g14590 ( 
.A1(n_14575),
.A2(n_2193),
.B(n_2194),
.Y(n_14590)
);

XNOR2x2_ASAP7_75t_L g14591 ( 
.A(n_14554),
.B(n_2195),
.Y(n_14591)
);

NAND3xp33_ASAP7_75t_L g14592 ( 
.A(n_14551),
.B(n_2195),
.C(n_2196),
.Y(n_14592)
);

OA211x2_ASAP7_75t_L g14593 ( 
.A1(n_14553),
.A2(n_2198),
.B(n_2196),
.C(n_2197),
.Y(n_14593)
);

OR2x2_ASAP7_75t_L g14594 ( 
.A(n_14563),
.B(n_2197),
.Y(n_14594)
);

NAND2xp5_ASAP7_75t_L g14595 ( 
.A(n_14565),
.B(n_2198),
.Y(n_14595)
);

OAI211xp5_ASAP7_75t_L g14596 ( 
.A1(n_14550),
.A2(n_2200),
.B(n_2198),
.C(n_2199),
.Y(n_14596)
);

NAND2xp5_ASAP7_75t_L g14597 ( 
.A(n_14557),
.B(n_2199),
.Y(n_14597)
);

AND2x2_ASAP7_75t_L g14598 ( 
.A(n_14552),
.B(n_2200),
.Y(n_14598)
);

NOR2x1_ASAP7_75t_L g14599 ( 
.A(n_14556),
.B(n_2201),
.Y(n_14599)
);

INVx2_ASAP7_75t_SL g14600 ( 
.A(n_14562),
.Y(n_14600)
);

NAND2xp5_ASAP7_75t_SL g14601 ( 
.A(n_14578),
.B(n_2201),
.Y(n_14601)
);

HB1xp67_ASAP7_75t_L g14602 ( 
.A(n_14566),
.Y(n_14602)
);

INVx1_ASAP7_75t_L g14603 ( 
.A(n_14561),
.Y(n_14603)
);

NOR2xp33_ASAP7_75t_L g14604 ( 
.A(n_14582),
.B(n_14558),
.Y(n_14604)
);

NOR3xp33_ASAP7_75t_L g14605 ( 
.A(n_14586),
.B(n_14588),
.C(n_14589),
.Y(n_14605)
);

NAND5xp2_ASAP7_75t_L g14606 ( 
.A(n_14585),
.B(n_14571),
.C(n_14555),
.D(n_14573),
.E(n_14574),
.Y(n_14606)
);

NOR2x1p5_ASAP7_75t_L g14607 ( 
.A(n_14583),
.B(n_14579),
.Y(n_14607)
);

AOI211xp5_ASAP7_75t_L g14608 ( 
.A1(n_14590),
.A2(n_14576),
.B(n_14567),
.C(n_2203),
.Y(n_14608)
);

NOR3xp33_ASAP7_75t_L g14609 ( 
.A(n_14587),
.B(n_2201),
.C(n_2202),
.Y(n_14609)
);

NOR3xp33_ASAP7_75t_L g14610 ( 
.A(n_14603),
.B(n_2202),
.C(n_2204),
.Y(n_14610)
);

INVx2_ASAP7_75t_L g14611 ( 
.A(n_14591),
.Y(n_14611)
);

NOR2xp67_ASAP7_75t_SL g14612 ( 
.A(n_14602),
.B(n_14581),
.Y(n_14612)
);

AOI211xp5_ASAP7_75t_L g14613 ( 
.A1(n_14596),
.A2(n_2205),
.B(n_2202),
.C(n_2204),
.Y(n_14613)
);

AOI21xp5_ASAP7_75t_L g14614 ( 
.A1(n_14601),
.A2(n_2205),
.B(n_2206),
.Y(n_14614)
);

NAND2xp5_ASAP7_75t_L g14615 ( 
.A(n_14584),
.B(n_2206),
.Y(n_14615)
);

A2O1A1Ixp33_ASAP7_75t_L g14616 ( 
.A1(n_14592),
.A2(n_2208),
.B(n_2206),
.C(n_2207),
.Y(n_14616)
);

NOR3xp33_ASAP7_75t_L g14617 ( 
.A(n_14600),
.B(n_2207),
.C(n_2208),
.Y(n_14617)
);

NOR3xp33_ASAP7_75t_L g14618 ( 
.A(n_14597),
.B(n_2207),
.C(n_2208),
.Y(n_14618)
);

NOR4xp25_ASAP7_75t_L g14619 ( 
.A(n_14598),
.B(n_2211),
.C(n_2209),
.D(n_2210),
.Y(n_14619)
);

NOR3xp33_ASAP7_75t_L g14620 ( 
.A(n_14595),
.B(n_2209),
.C(n_2210),
.Y(n_14620)
);

NAND3xp33_ASAP7_75t_L g14621 ( 
.A(n_14599),
.B(n_2209),
.C(n_2211),
.Y(n_14621)
);

OAI211xp5_ASAP7_75t_L g14622 ( 
.A1(n_14594),
.A2(n_2213),
.B(n_2211),
.C(n_2212),
.Y(n_14622)
);

NAND3xp33_ASAP7_75t_SL g14623 ( 
.A(n_14593),
.B(n_2212),
.C(n_2213),
.Y(n_14623)
);

NAND2xp5_ASAP7_75t_L g14624 ( 
.A(n_14586),
.B(n_2213),
.Y(n_14624)
);

INVx1_ASAP7_75t_L g14625 ( 
.A(n_14612),
.Y(n_14625)
);

OA21x2_ASAP7_75t_L g14626 ( 
.A1(n_14615),
.A2(n_2214),
.B(n_2215),
.Y(n_14626)
);

NOR2xp33_ASAP7_75t_L g14627 ( 
.A(n_14623),
.B(n_14611),
.Y(n_14627)
);

OAI21xp33_ASAP7_75t_SL g14628 ( 
.A1(n_14607),
.A2(n_14604),
.B(n_14619),
.Y(n_14628)
);

INVx1_ASAP7_75t_L g14629 ( 
.A(n_14621),
.Y(n_14629)
);

INVx1_ASAP7_75t_SL g14630 ( 
.A(n_14624),
.Y(n_14630)
);

INVxp67_ASAP7_75t_L g14631 ( 
.A(n_14605),
.Y(n_14631)
);

XNOR2x1_ASAP7_75t_SL g14632 ( 
.A(n_14606),
.B(n_2214),
.Y(n_14632)
);

INVx1_ASAP7_75t_L g14633 ( 
.A(n_14609),
.Y(n_14633)
);

INVx1_ASAP7_75t_L g14634 ( 
.A(n_14622),
.Y(n_14634)
);

AND2x2_ASAP7_75t_L g14635 ( 
.A(n_14618),
.B(n_2215),
.Y(n_14635)
);

INVx1_ASAP7_75t_SL g14636 ( 
.A(n_14614),
.Y(n_14636)
);

NOR2x1_ASAP7_75t_L g14637 ( 
.A(n_14616),
.B(n_2215),
.Y(n_14637)
);

NAND2xp5_ASAP7_75t_L g14638 ( 
.A(n_14620),
.B(n_2216),
.Y(n_14638)
);

INVxp67_ASAP7_75t_SL g14639 ( 
.A(n_14610),
.Y(n_14639)
);

INVx1_ASAP7_75t_L g14640 ( 
.A(n_14617),
.Y(n_14640)
);

NOR2x1_ASAP7_75t_L g14641 ( 
.A(n_14613),
.B(n_2216),
.Y(n_14641)
);

NAND2xp5_ASAP7_75t_L g14642 ( 
.A(n_14608),
.B(n_2217),
.Y(n_14642)
);

INVx1_ASAP7_75t_L g14643 ( 
.A(n_14612),
.Y(n_14643)
);

AND2x4_ASAP7_75t_L g14644 ( 
.A(n_14643),
.B(n_2217),
.Y(n_14644)
);

INVx1_ASAP7_75t_L g14645 ( 
.A(n_14632),
.Y(n_14645)
);

NAND3xp33_ASAP7_75t_L g14646 ( 
.A(n_14625),
.B(n_2217),
.C(n_2218),
.Y(n_14646)
);

NOR3xp33_ASAP7_75t_L g14647 ( 
.A(n_14631),
.B(n_2218),
.C(n_2219),
.Y(n_14647)
);

NOR2x1_ASAP7_75t_L g14648 ( 
.A(n_14627),
.B(n_2219),
.Y(n_14648)
);

NOR2xp33_ASAP7_75t_L g14649 ( 
.A(n_14628),
.B(n_2220),
.Y(n_14649)
);

BUFx2_ASAP7_75t_L g14650 ( 
.A(n_14626),
.Y(n_14650)
);

NAND4xp25_ASAP7_75t_L g14651 ( 
.A(n_14641),
.B(n_2222),
.C(n_2220),
.D(n_2221),
.Y(n_14651)
);

NOR3x1_ASAP7_75t_L g14652 ( 
.A(n_14642),
.B(n_2221),
.C(n_2222),
.Y(n_14652)
);

NAND2xp5_ASAP7_75t_L g14653 ( 
.A(n_14630),
.B(n_14639),
.Y(n_14653)
);

NOR2x1_ASAP7_75t_L g14654 ( 
.A(n_14634),
.B(n_2222),
.Y(n_14654)
);

NAND2x1p5_ASAP7_75t_L g14655 ( 
.A(n_14636),
.B(n_2223),
.Y(n_14655)
);

AND5x1_ASAP7_75t_L g14656 ( 
.A(n_14637),
.B(n_14633),
.C(n_14629),
.D(n_14640),
.E(n_14638),
.Y(n_14656)
);

NOR2x1_ASAP7_75t_L g14657 ( 
.A(n_14650),
.B(n_14626),
.Y(n_14657)
);

INVx1_ASAP7_75t_L g14658 ( 
.A(n_14655),
.Y(n_14658)
);

INVx1_ASAP7_75t_L g14659 ( 
.A(n_14648),
.Y(n_14659)
);

AOI22xp5_ASAP7_75t_L g14660 ( 
.A1(n_14645),
.A2(n_14635),
.B1(n_2225),
.B2(n_2223),
.Y(n_14660)
);

AO22x2_ASAP7_75t_L g14661 ( 
.A1(n_14653),
.A2(n_2225),
.B1(n_2223),
.B2(n_2224),
.Y(n_14661)
);

AOI22xp5_ASAP7_75t_L g14662 ( 
.A1(n_14649),
.A2(n_14647),
.B1(n_14651),
.B2(n_14646),
.Y(n_14662)
);

AND2x2_ASAP7_75t_L g14663 ( 
.A(n_14654),
.B(n_14652),
.Y(n_14663)
);

INVx2_ASAP7_75t_L g14664 ( 
.A(n_14644),
.Y(n_14664)
);

AND2x4_ASAP7_75t_L g14665 ( 
.A(n_14664),
.B(n_14656),
.Y(n_14665)
);

NAND2xp5_ASAP7_75t_SL g14666 ( 
.A(n_14657),
.B(n_14644),
.Y(n_14666)
);

NAND4xp75_ASAP7_75t_L g14667 ( 
.A(n_14659),
.B(n_2227),
.C(n_2224),
.D(n_2226),
.Y(n_14667)
);

AOI21xp5_ASAP7_75t_L g14668 ( 
.A1(n_14663),
.A2(n_2224),
.B(n_2226),
.Y(n_14668)
);

NAND2xp5_ASAP7_75t_L g14669 ( 
.A(n_14658),
.B(n_2227),
.Y(n_14669)
);

NAND4xp75_ASAP7_75t_L g14670 ( 
.A(n_14666),
.B(n_14660),
.C(n_14662),
.D(n_14661),
.Y(n_14670)
);

OR4x1_ASAP7_75t_L g14671 ( 
.A(n_14665),
.B(n_2398),
.C(n_2230),
.D(n_2228),
.Y(n_14671)
);

AND3x2_ASAP7_75t_L g14672 ( 
.A(n_14669),
.B(n_2229),
.C(n_2230),
.Y(n_14672)
);

NOR2x1_ASAP7_75t_L g14673 ( 
.A(n_14667),
.B(n_2229),
.Y(n_14673)
);

INVx1_ASAP7_75t_L g14674 ( 
.A(n_14670),
.Y(n_14674)
);

NOR3xp33_ASAP7_75t_L g14675 ( 
.A(n_14673),
.B(n_14668),
.C(n_2230),
.Y(n_14675)
);

A2O1A1Ixp33_ASAP7_75t_L g14676 ( 
.A1(n_14674),
.A2(n_14671),
.B(n_14672),
.C(n_2233),
.Y(n_14676)
);

OAI221xp5_ASAP7_75t_L g14677 ( 
.A1(n_14675),
.A2(n_2233),
.B1(n_2231),
.B2(n_2232),
.C(n_2234),
.Y(n_14677)
);

INVx1_ASAP7_75t_L g14678 ( 
.A(n_14674),
.Y(n_14678)
);

INVx1_ASAP7_75t_L g14679 ( 
.A(n_14678),
.Y(n_14679)
);

INVx2_ASAP7_75t_L g14680 ( 
.A(n_14677),
.Y(n_14680)
);

INVx1_ASAP7_75t_L g14681 ( 
.A(n_14676),
.Y(n_14681)
);

AND2x2_ASAP7_75t_SL g14682 ( 
.A(n_14679),
.B(n_2231),
.Y(n_14682)
);

INVx2_ASAP7_75t_L g14683 ( 
.A(n_14681),
.Y(n_14683)
);

INVx2_ASAP7_75t_L g14684 ( 
.A(n_14680),
.Y(n_14684)
);

XNOR2x2_ASAP7_75t_L g14685 ( 
.A(n_14683),
.B(n_2231),
.Y(n_14685)
);

INVxp67_ASAP7_75t_SL g14686 ( 
.A(n_14684),
.Y(n_14686)
);

NOR2xp33_ASAP7_75t_L g14687 ( 
.A(n_14682),
.B(n_2232),
.Y(n_14687)
);

INVx1_ASAP7_75t_L g14688 ( 
.A(n_14686),
.Y(n_14688)
);

NAND2xp33_ASAP7_75t_SL g14689 ( 
.A(n_14685),
.B(n_2232),
.Y(n_14689)
);

AOI22xp5_ASAP7_75t_L g14690 ( 
.A1(n_14687),
.A2(n_2235),
.B1(n_2233),
.B2(n_2234),
.Y(n_14690)
);

OAI22xp5_ASAP7_75t_L g14691 ( 
.A1(n_14688),
.A2(n_2236),
.B1(n_2234),
.B2(n_2235),
.Y(n_14691)
);

NOR2xp67_ASAP7_75t_L g14692 ( 
.A(n_14690),
.B(n_2235),
.Y(n_14692)
);

XNOR2xp5_ASAP7_75t_L g14693 ( 
.A(n_14692),
.B(n_14689),
.Y(n_14693)
);

AOI221xp5_ASAP7_75t_L g14694 ( 
.A1(n_14693),
.A2(n_14691),
.B1(n_2238),
.B2(n_2236),
.C(n_2237),
.Y(n_14694)
);

AOI22x1_ASAP7_75t_L g14695 ( 
.A1(n_14694),
.A2(n_2238),
.B1(n_2236),
.B2(n_2237),
.Y(n_14695)
);

AOI221xp5_ASAP7_75t_L g14696 ( 
.A1(n_14695),
.A2(n_2240),
.B1(n_2238),
.B2(n_2239),
.C(n_2242),
.Y(n_14696)
);

NAND2xp5_ASAP7_75t_SL g14697 ( 
.A(n_14695),
.B(n_2239),
.Y(n_14697)
);

INVx4_ASAP7_75t_L g14698 ( 
.A(n_14697),
.Y(n_14698)
);

BUFx3_ASAP7_75t_L g14699 ( 
.A(n_14696),
.Y(n_14699)
);

OA21x2_ASAP7_75t_L g14700 ( 
.A1(n_14698),
.A2(n_2240),
.B(n_2242),
.Y(n_14700)
);

OR2x6_ASAP7_75t_L g14701 ( 
.A(n_14699),
.B(n_2240),
.Y(n_14701)
);

AOI221xp5_ASAP7_75t_L g14702 ( 
.A1(n_14701),
.A2(n_2244),
.B1(n_2242),
.B2(n_2243),
.C(n_2245),
.Y(n_14702)
);

AOI22xp5_ASAP7_75t_L g14703 ( 
.A1(n_14700),
.A2(n_2245),
.B1(n_2243),
.B2(n_2244),
.Y(n_14703)
);

AOI21xp33_ASAP7_75t_L g14704 ( 
.A1(n_14703),
.A2(n_2243),
.B(n_2244),
.Y(n_14704)
);

AOI211xp5_ASAP7_75t_L g14705 ( 
.A1(n_14704),
.A2(n_14702),
.B(n_2246),
.C(n_2245),
.Y(n_14705)
);


endmodule