module fake_jpeg_11504_n_139 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_7),
.B(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_13),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_1),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_3),
.Y(n_39)
);

AO22x1_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_24),
.B1(n_18),
.B2(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_45),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_24),
.B(n_18),
.C(n_23),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_22),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_38),
.A3(n_24),
.B1(n_15),
.B2(n_28),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_18),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_3),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_15),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_25),
.B1(n_22),
.B2(n_19),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_19),
.B1(n_21),
.B2(n_20),
.Y(n_62)
);

OA21x2_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_40),
.B(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_73),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_68),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_28),
.B1(n_21),
.B2(n_20),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_66),
.B1(n_14),
.B2(n_40),
.Y(n_86)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_3),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_11),
.C(n_7),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_41),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_5),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_26),
.Y(n_73)
);

A2O1A1O1Ixp25_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_53),
.B(n_45),
.C(n_44),
.D(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_80),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_14),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_87),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_61),
.B1(n_42),
.B2(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_46),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_55),
.B(n_66),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_72),
.C(n_64),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_92),
.C(n_79),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_72),
.C(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_84),
.B(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_99),
.Y(n_107)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_55),
.B(n_71),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_78),
.B(n_88),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_89),
.B1(n_78),
.B2(n_85),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_109),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_106),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_83),
.A3(n_76),
.B1(n_10),
.B2(n_12),
.C1(n_9),
.C2(n_86),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_65),
.C(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_94),
.B1(n_100),
.B2(n_101),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_98),
.B1(n_92),
.B2(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_121),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_125),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_104),
.C(n_111),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_127),
.B(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_90),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_130),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_120),
.B1(n_121),
.B2(n_117),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_115),
.A3(n_114),
.B1(n_110),
.B2(n_113),
.C1(n_103),
.C2(n_93),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_125),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_135),
.C(n_133),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_95),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_133),
.C(n_56),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_136),
.Y(n_139)
);


endmodule