module fake_netlist_1_7148_n_25 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_25);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_13), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_17) );
NOR2xp33_ASAP7_75t_SL g18 ( .A(n_14), .B(n_7), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_17), .B(n_15), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_18), .B1(n_16), .B2(n_2), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_16), .B(n_4), .Y(n_21) );
NAND4xp25_ASAP7_75t_L g22 ( .A(n_21), .B(n_16), .C(n_5), .D(n_9), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_3), .Y(n_23) );
BUFx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_25) );
endmodule