module fake_netlist_1_4042_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_8), .B(n_6), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_0), .B(n_4), .Y(n_15) );
AOI22xp33_ASAP7_75t_L g16 ( .A1(n_12), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_13), .B(n_15), .Y(n_20) );
INVx2_ASAP7_75t_SL g21 ( .A(n_20), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_19), .B(n_14), .Y(n_22) );
INVx5_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_19), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_23), .A2(n_16), .B1(n_13), .B2(n_4), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
AOI221xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_23), .B1(n_3), .B2(n_5), .C(n_2), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
NAND2x1_ASAP7_75t_SL g30 ( .A(n_27), .B(n_23), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
NOR4xp75_ASAP7_75t_L g32 ( .A(n_28), .B(n_5), .C(n_9), .D(n_10), .Y(n_32) );
OAI21xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_23), .B(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
AOI22xp5_ASAP7_75t_SL g36 ( .A1(n_35), .A2(n_34), .B1(n_33), .B2(n_32), .Y(n_36) );
endmodule