module fake_jpeg_30356_n_503 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_13),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_0),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_53),
.B(n_55),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_54),
.A2(n_25),
.B1(n_46),
.B2(n_45),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_58),
.Y(n_105)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_61),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_26),
.B(n_50),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_65),
.B(n_75),
.Y(n_156)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_40),
.B(n_12),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_69),
.B(n_74),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_30),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_26),
.B(n_0),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx4f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_35),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_94),
.B(n_96),
.Y(n_155)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_16),
.B(n_0),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_48),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_0),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_45),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_115),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g169 ( 
.A(n_107),
.Y(n_169)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_53),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_150),
.Y(n_163)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_63),
.A2(n_39),
.B(n_35),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_132),
.B(n_137),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_60),
.A2(n_36),
.B1(n_42),
.B2(n_33),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_136),
.A2(n_139),
.B1(n_46),
.B2(n_22),
.Y(n_194)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_78),
.B(n_25),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_48),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_79),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_71),
.A2(n_36),
.B1(n_38),
.B2(n_31),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_73),
.B1(n_31),
.B2(n_70),
.Y(n_166)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_82),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_162),
.B(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_165),
.B(n_168),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_166),
.A2(n_180),
.B1(n_181),
.B2(n_107),
.Y(n_234)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_84),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_105),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_176),
.Y(n_209)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_106),
.Y(n_176)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_85),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_178),
.B(n_37),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_88),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_186),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_73),
.B1(n_95),
.B2(n_93),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_110),
.A2(n_112),
.B1(n_64),
.B2(n_43),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_117),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_128),
.Y(n_187)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

CKINVDCx12_ASAP7_75t_R g189 ( 
.A(n_116),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

CKINVDCx9p33_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

BUFx8_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_127),
.A2(n_97),
.B1(n_91),
.B2(n_81),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_192),
.A2(n_194),
.B1(n_20),
.B2(n_80),
.Y(n_249)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_126),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_197),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_156),
.Y(n_197)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_90),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_199),
.B(n_200),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

BUFx16f_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_203),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_51),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_206),
.Y(n_229)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_101),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_144),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_151),
.C(n_113),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_211),
.B(n_87),
.C(n_148),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_163),
.A2(n_142),
.B1(n_127),
.B2(n_122),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_213),
.A2(n_249),
.B1(n_144),
.B2(n_103),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_161),
.B(n_102),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g258 ( 
.A1(n_215),
.A2(n_234),
.B(n_247),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_201),
.B(n_23),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_220),
.B(n_107),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_166),
.A2(n_180),
.B(n_200),
.C(n_181),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_239),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_37),
.B(n_23),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_224),
.A2(n_236),
.B(n_248),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_159),
.B(n_111),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_232),
.B(n_235),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_142),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_177),
.A2(n_103),
.B(n_39),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_240),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_57),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_145),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_192),
.A2(n_66),
.B1(n_92),
.B2(n_52),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_169),
.A2(n_22),
.B(n_20),
.Y(n_248)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_203),
.Y(n_252)
);

A2O1A1O1Ixp25_ASAP7_75t_L g315 ( 
.A1(n_252),
.A2(n_257),
.B(n_264),
.C(n_169),
.D(n_245),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_222),
.A2(n_112),
.B1(n_158),
.B2(n_167),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_254),
.A2(n_278),
.B1(n_286),
.B2(n_268),
.Y(n_320)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

AND2x6_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_262),
.B(n_268),
.Y(n_304)
);

CKINVDCx12_ASAP7_75t_R g263 ( 
.A(n_221),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_263),
.Y(n_294)
);

OR2x4_ASAP7_75t_L g264 ( 
.A(n_215),
.B(n_236),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_241),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_205),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_269),
.B(n_270),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_210),
.B(n_185),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_214),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_271),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_209),
.B(n_198),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_272),
.B(n_273),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_215),
.A2(n_145),
.B1(n_122),
.B2(n_135),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_288),
.B1(n_230),
.B2(n_243),
.Y(n_295)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_275),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_276),
.B(n_169),
.Y(n_321)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_212),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_279),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_223),
.B(n_123),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_280),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_239),
.B1(n_225),
.B2(n_229),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_237),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_216),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_241),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_289),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_249),
.A2(n_135),
.B1(n_207),
.B2(n_171),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_225),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_290),
.A2(n_295),
.B1(n_301),
.B2(n_313),
.Y(n_336)
);

AO22x1_ASAP7_75t_SL g291 ( 
.A1(n_259),
.A2(n_247),
.B1(n_243),
.B2(n_238),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_318),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_255),
.A2(n_248),
.B(n_224),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_293),
.A2(n_310),
.B(n_315),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_218),
.C(n_267),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_319),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_250),
.C(n_218),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_321),
.C(n_289),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_273),
.A2(n_247),
.B1(n_242),
.B2(n_226),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_255),
.A2(n_230),
.B(n_245),
.Y(n_310)
);

OAI32xp33_ASAP7_75t_L g311 ( 
.A1(n_285),
.A2(n_250),
.A3(n_247),
.B1(n_238),
.B2(n_219),
.Y(n_311)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_285),
.A2(n_187),
.B1(n_160),
.B2(n_242),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_264),
.A2(n_219),
.B(n_227),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_317),
.A2(n_231),
.B(n_278),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_260),
.B(n_253),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_121),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_253),
.B(n_227),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_279),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_288),
.A2(n_266),
.B1(n_258),
.B2(n_274),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_325),
.A2(n_258),
.B1(n_281),
.B2(n_257),
.Y(n_344)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_316),
.Y(n_327)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_327),
.Y(n_369)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_328),
.Y(n_372)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_252),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_329),
.A2(n_358),
.B(n_307),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_262),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_330),
.B(n_333),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_331),
.B(n_355),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_296),
.B(n_284),
.Y(n_333)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_334),
.Y(n_384)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_338),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_318),
.B(n_283),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_340),
.B(n_342),
.Y(n_376)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_341),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_343),
.B(n_346),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_344),
.A2(n_357),
.B1(n_323),
.B2(n_307),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_348),
.Y(n_360)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_265),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_349),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_305),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_308),
.B(n_277),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_352),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_287),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_354),
.Y(n_367)
);

NOR4xp25_ASAP7_75t_SL g352 ( 
.A(n_311),
.B(n_271),
.C(n_251),
.D(n_275),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_353),
.A2(n_309),
.B(n_291),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

XNOR2x1_ASAP7_75t_L g355 ( 
.A(n_298),
.B(n_286),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_322),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_246),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_295),
.A2(n_246),
.B1(n_208),
.B2(n_256),
.Y(n_357)
);

AOI22x1_ASAP7_75t_SL g358 ( 
.A1(n_293),
.A2(n_226),
.B1(n_208),
.B2(n_231),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_361),
.A2(n_326),
.B1(n_353),
.B2(n_341),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_331),
.B(n_321),
.C(n_319),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_370),
.C(n_381),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_317),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_364),
.B(n_368),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_351),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_366),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_345),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_292),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_355),
.B(n_292),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_314),
.Y(n_371)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_354),
.A2(n_309),
.B(n_299),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_374),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_313),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_378),
.B(n_190),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_291),
.Y(n_380)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_380),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_332),
.B(n_306),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_335),
.A2(n_303),
.B(n_302),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_385),
.B(n_126),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_297),
.Y(n_388)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_388),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_389),
.A2(n_391),
.B1(n_395),
.B2(n_410),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_375),
.A2(n_326),
.B1(n_337),
.B2(n_338),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_332),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_392),
.B(n_407),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_375),
.A2(n_337),
.B1(n_344),
.B2(n_336),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_382),
.A2(n_336),
.B1(n_357),
.B2(n_329),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_397),
.A2(n_406),
.B1(n_414),
.B2(n_404),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_328),
.C(n_334),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_409),
.C(n_364),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_402),
.B(n_378),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_403),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_359),
.A2(n_42),
.B1(n_297),
.B2(n_38),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_148),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_373),
.B(n_182),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_413),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_175),
.C(n_172),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_361),
.A2(n_108),
.B1(n_172),
.B2(n_157),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_365),
.A2(n_190),
.B1(n_42),
.B2(n_157),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_412),
.A2(n_387),
.B1(n_371),
.B2(n_360),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_1),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_368),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_415),
.B(n_417),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_381),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_419),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_377),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_420),
.B(n_421),
.Y(n_448)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_367),
.C(n_370),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_367),
.C(n_374),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_431),
.C(n_432),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_411),
.A2(n_380),
.B1(n_366),
.B2(n_369),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_423),
.B(n_424),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_395),
.A2(n_369),
.B1(n_383),
.B2(n_360),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_433),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_427),
.A2(n_428),
.B1(n_410),
.B2(n_389),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_398),
.A2(n_383),
.B1(n_372),
.B2(n_384),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_399),
.B(n_385),
.Y(n_429)
);

XNOR2x1_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_2),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_68),
.C(n_43),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_393),
.B(n_43),
.C(n_41),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_390),
.A2(n_41),
.B(n_3),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_41),
.C(n_27),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_400),
.C(n_412),
.Y(n_444)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_436),
.Y(n_453)
);

BUFx12_ASAP7_75t_L g438 ( 
.A(n_434),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_445),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_430),
.A2(n_391),
.B1(n_405),
.B2(n_394),
.Y(n_440)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_440),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_430),
.A2(n_405),
.B(n_390),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_441),
.A2(n_435),
.B(n_431),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_450),
.Y(n_454)
);

INVx13_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_400),
.C(n_414),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_429),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_418),
.B(n_2),
.Y(n_449)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_449),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_417),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_451),
.B(n_420),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_452),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_446),
.B(n_421),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_455),
.B(n_458),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_416),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_438),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_462),
.B(n_463),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_437),
.A2(n_432),
.B1(n_415),
.B2(n_5),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_465),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_444),
.A2(n_452),
.B1(n_441),
.B2(n_439),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_467),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_443),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_453),
.A2(n_456),
.B1(n_461),
.B2(n_459),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_7),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_467),
.B(n_443),
.C(n_439),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_471),
.C(n_454),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_448),
.C(n_450),
.Y(n_471)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_472),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_457),
.A2(n_438),
.B1(n_445),
.B2(n_448),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_473),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_2),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_477),
.Y(n_484)
);

XNOR2x1_ASAP7_75t_L g477 ( 
.A(n_454),
.B(n_4),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_460),
.A2(n_5),
.B(n_7),
.Y(n_478)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_478),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_485),
.C(n_476),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_482),
.B(n_483),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_472),
.B(n_8),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_8),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_486),
.B(n_487),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_9),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_492),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_475),
.C(n_470),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_480),
.B(n_479),
.Y(n_493)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_493),
.Y(n_495)
);

NOR2x1_ASAP7_75t_L g494 ( 
.A(n_491),
.B(n_488),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_490),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_497),
.A2(n_498),
.B(n_495),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_471),
.B(n_477),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_499),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_500),
.B(n_485),
.C(n_484),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_501),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_502),
.B(n_484),
.Y(n_503)
);


endmodule