module fake_jpeg_7695_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_2),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_22),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_17)
);

AO21x2_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_24),
.B(n_25),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_5),
.B(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_16),
.B1(n_21),
.B2(n_9),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_37),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_27),
.B1(n_33),
.B2(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_30),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.C(n_16),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_34),
.B(n_26),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_9),
.Y(n_43)
);


endmodule