module real_jpeg_1098_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_1),
.A2(n_31),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_1),
.A2(n_37),
.B1(n_43),
.B2(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_1),
.A2(n_37),
.B1(n_65),
.B2(n_67),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_1),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_2),
.A2(n_43),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_52),
.B1(n_65),
.B2(n_67),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_31),
.B1(n_38),
.B2(n_52),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_2),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_3),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_3),
.A2(n_65),
.B1(n_67),
.B2(n_69),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_3),
.A2(n_43),
.B1(n_45),
.B2(n_69),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_31),
.B1(n_38),
.B2(n_69),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_5),
.A2(n_65),
.B1(n_67),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_77),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_5),
.A2(n_43),
.B1(n_45),
.B2(n_77),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_31),
.B1(n_38),
.B2(n_77),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_6),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_6),
.A2(n_65),
.B1(n_67),
.B2(n_127),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_6),
.A2(n_43),
.B1(n_45),
.B2(n_127),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_6),
.A2(n_31),
.B1(n_38),
.B2(n_127),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_7),
.B(n_59),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_7),
.B(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_7),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_7),
.A2(n_59),
.B(n_171),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_7),
.B(n_80),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_7),
.A2(n_67),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_7),
.B(n_31),
.C(n_48),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_7),
.A2(n_43),
.B1(n_45),
.B2(n_207),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_7),
.B(n_34),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_7),
.B(n_53),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_12),
.A2(n_42),
.B1(n_65),
.B2(n_67),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_12),
.A2(n_42),
.B1(n_59),
.B2(n_60),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_12),
.A2(n_31),
.B1(n_38),
.B2(n_42),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_13),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_13),
.A2(n_65),
.B1(n_67),
.B2(n_161),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_13),
.A2(n_43),
.B1(n_45),
.B2(n_161),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_13),
.A2(n_31),
.B1(n_38),
.B2(n_161),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_14),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_14),
.A2(n_65),
.B1(n_67),
.B2(n_181),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_14),
.A2(n_43),
.B1(n_45),
.B2(n_181),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_14),
.A2(n_31),
.B1(n_38),
.B2(n_181),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_15),
.A2(n_65),
.B1(n_67),
.B2(n_71),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_15),
.A2(n_43),
.B1(n_45),
.B2(n_71),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g198 ( 
.A1(n_15),
.A2(n_31),
.B1(n_38),
.B2(n_71),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_315),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_302),
.B(n_314),
.Y(n_20)
);

AO21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_141),
.B(n_299),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_128),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_101),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_24),
.B(n_101),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_72),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_25),
.B(n_87),
.C(n_99),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_54),
.B(n_55),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_26),
.A2(n_27),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_28),
.A2(n_54),
.B1(n_55),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_28),
.A2(n_39),
.B1(n_40),
.B2(n_54),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B(n_35),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_29),
.A2(n_33),
.B1(n_115),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_29),
.A2(n_33),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_29),
.A2(n_33),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_30),
.A2(n_34),
.B1(n_36),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_30),
.A2(n_34),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_30),
.A2(n_34),
.B1(n_174),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_30),
.A2(n_34),
.B1(n_211),
.B2(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_30),
.A2(n_34),
.B1(n_207),
.B2(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_30),
.A2(n_34),
.B1(n_261),
.B2(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_31),
.B(n_259),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_41),
.A2(n_46),
.B1(n_53),
.B2(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_45),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_43),
.A2(n_67),
.A3(n_81),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_43),
.B(n_249),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_45),
.B(n_82),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_51),
.B1(n_53),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_53),
.B(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_46),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_46),
.A2(n_53),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_46),
.A2(n_53),
.B1(n_203),
.B2(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_46),
.A2(n_53),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_46),
.A2(n_53),
.B1(n_231),
.B2(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_50),
.A2(n_119),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_50),
.A2(n_154),
.B1(n_202),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_64),
.B1(n_68),
.B2(n_70),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_64),
.B1(n_70),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_56),
.A2(n_64),
.B1(n_68),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_56),
.A2(n_64),
.B1(n_90),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_56),
.A2(n_64),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_56),
.A2(n_64),
.B1(n_180),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_57),
.A2(n_126),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_57),
.A2(n_162),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_57),
.A2(n_162),
.B1(n_310),
.B2(n_318),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_64),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_60),
.A2(n_63),
.A3(n_67),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_62),
.B(n_65),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_64),
.Y(n_162)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_67),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_65),
.B(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_87),
.B1(n_99),
.B2(n_100),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_74),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_85),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_80),
.B2(n_84),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_79),
.B1(n_121),
.B2(n_123),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_80),
.B1(n_84),
.B2(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_78),
.A2(n_80),
.B1(n_122),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_78),
.A2(n_80),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_79),
.A2(n_97),
.B1(n_123),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_79),
.A2(n_123),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_79),
.A2(n_123),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_79),
.A2(n_123),
.B1(n_177),
.B2(n_193),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_79),
.A2(n_123),
.B1(n_192),
.B2(n_240),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_89),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_93),
.C(n_95),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_89),
.B(n_132),
.C(n_139),
.Y(n_303)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_98),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_98),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_93),
.B(n_135),
.C(n_137),
.Y(n_313)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_109),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_120),
.C(n_124),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_111),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_124),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_128),
.A2(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_140),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_129),
.B(n_140),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_136),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_138),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_163),
.B(n_298),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_143),
.B(n_145),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_149),
.Y(n_185)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_157),
.C(n_159),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_152),
.B(n_155),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_153),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_159),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_186),
.B(n_297),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_184),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_165),
.B(n_184),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.C(n_183),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_166),
.B(n_183),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_168),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.C(n_179),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_169),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_173),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_176),
.B(n_179),
.Y(n_287)
);

AOI31xp33_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_281),
.A3(n_290),
.B(n_294),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_226),
.B(n_280),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_213),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_189),
.B(n_213),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_200),
.C(n_204),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_190),
.B(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_195),
.C(n_199),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_199),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_200),
.B(n_204),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_215),
.B(n_216),
.C(n_217),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_221),
.C(n_225),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_275),
.B(n_279),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_244),
.B(n_274),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_236),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.C(n_234),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_233),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_239),
.C(n_242),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_255),
.B(n_273),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_267),
.B(n_272),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_262),
.B(n_266),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_271),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_278),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_285),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.C(n_289),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_289),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_313),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_308),
.B1(n_311),
.B2(n_312),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_306),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_308),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_311),
.C(n_313),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_320),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);


endmodule