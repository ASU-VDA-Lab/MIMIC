module fake_jpeg_21243_n_184 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_28),
.Y(n_41)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_6),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_23),
.C(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_43),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_28),
.B(n_24),
.C(n_29),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_16),
.B(n_17),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_15),
.B1(n_17),
.B2(n_16),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_18),
.B1(n_23),
.B2(n_12),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_13),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_34),
.B1(n_39),
.B2(n_35),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_31),
.B1(n_27),
.B2(n_16),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_59),
.B1(n_35),
.B2(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_27),
.B1(n_17),
.B2(n_13),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_54),
.B1(n_42),
.B2(n_36),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_55),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_27),
.B1(n_18),
.B2(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_21),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_30),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_67),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_68),
.B1(n_72),
.B2(n_51),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_25),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_71),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_39),
.B1(n_44),
.B2(n_33),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_36),
.B1(n_30),
.B2(n_32),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_58),
.B1(n_48),
.B2(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_23),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_59),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_59),
.B(n_60),
.C(n_45),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_82),
.B(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_90),
.B1(n_66),
.B2(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_50),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_78),
.B1(n_69),
.B2(n_67),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_25),
.Y(n_100)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_46),
.B1(n_12),
.B2(n_22),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_22),
.A3(n_63),
.B1(n_70),
.B2(n_23),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_32),
.B1(n_25),
.B2(n_12),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_23),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_56),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_105),
.B1(n_113),
.B2(n_94),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_77),
.B1(n_62),
.B2(n_76),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_99),
.B1(n_108),
.B2(n_110),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_112),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_103),
.C(n_104),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_87),
.C(n_90),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_77),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_32),
.B1(n_12),
.B2(n_22),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_32),
.B1(n_70),
.B2(n_10),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_32),
.B1(n_70),
.B2(n_10),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_81),
.B(n_82),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_22),
.B1(n_19),
.B2(n_47),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_20),
.B(n_2),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_113),
.B1(n_107),
.B2(n_104),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_92),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_95),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_127),
.B1(n_99),
.B2(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_126),
.B(n_105),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_83),
.B1(n_80),
.B2(n_93),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_80),
.C(n_63),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_56),
.C(n_47),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_134),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_103),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_142),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_111),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

OAI322xp33_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_20),
.A3(n_8),
.B1(n_10),
.B2(n_7),
.C1(n_9),
.C2(n_19),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_129),
.C(n_120),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_140),
.C(n_136),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_126),
.B1(n_127),
.B2(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_121),
.C(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_152),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_151),
.B(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_141),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_119),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_146),
.C(n_143),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_130),
.C(n_118),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_20),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_114),
.B1(n_128),
.B2(n_118),
.Y(n_159)
);

OAI221xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_143),
.B1(n_146),
.B2(n_149),
.C(n_119),
.Y(n_162)
);

XOR2x1_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_132),
.Y(n_160)
);

AOI31xp33_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_142),
.A3(n_7),
.B(n_8),
.Y(n_167)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_164),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_168),
.B(n_153),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_170),
.B(n_173),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_0),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_166),
.B(n_156),
.C(n_164),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_9),
.B(n_2),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_166),
.A2(n_7),
.B1(n_9),
.B2(n_3),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_177),
.C(n_178),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_174),
.A2(n_0),
.B(n_2),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_170),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_179),
.A2(n_3),
.B(n_4),
.Y(n_182)
);

AOI321xp33_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_169),
.C(n_174),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_182),
.C(n_4),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_5),
.Y(n_184)
);


endmodule