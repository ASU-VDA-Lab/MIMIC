module fake_jpeg_12139_n_468 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_468);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_468;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_8),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_76),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_56),
.B(n_65),
.Y(n_143)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_6),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_20),
.B(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_69),
.B(n_74),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_73),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_9),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g114 ( 
.A(n_75),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_28),
.B(n_9),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_24),
.B(n_9),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_82),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_24),
.B(n_5),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_95),
.Y(n_120)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_96),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_93),
.B(n_94),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_43),
.B(n_5),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_37),
.B1(n_27),
.B2(n_26),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_102),
.A2(n_124),
.B1(n_138),
.B2(n_54),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_48),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_116),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_52),
.B(n_35),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_31),
.B1(n_27),
.B2(n_37),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_122),
.A2(n_126),
.B1(n_136),
.B2(n_150),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_47),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_123),
.B(n_142),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_77),
.A2(n_37),
.B1(n_27),
.B2(n_31),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_43),
.B1(n_42),
.B2(n_29),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_70),
.A2(n_46),
.B1(n_45),
.B2(n_34),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_49),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_53),
.B(n_44),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_94),
.C(n_93),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_72),
.B(n_96),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_60),
.B(n_40),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_0),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_79),
.A2(n_34),
.B1(n_29),
.B2(n_38),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_59),
.B1(n_67),
.B2(n_66),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_84),
.A2(n_40),
.B1(n_38),
.B2(n_33),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_61),
.B(n_44),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_61),
.Y(n_189)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_152),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_83),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_153),
.B(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_154),
.B(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_89),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_158),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_128),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g223 ( 
.A(n_159),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_92),
.C(n_78),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_160),
.B(n_189),
.C(n_195),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_62),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_162),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_110),
.A2(n_88),
.B1(n_87),
.B2(n_86),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_164),
.A2(n_168),
.B1(n_196),
.B2(n_159),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_115),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_170),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_191),
.Y(n_209)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_116),
.B(n_90),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_173),
.B(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_0),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_177),
.B(n_190),
.Y(n_237)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_184),
.B(n_188),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_122),
.A2(n_58),
.B1(n_73),
.B2(n_71),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_186),
.Y(n_224)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_125),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_75),
.B(n_55),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_128),
.B(n_1),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_1),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_104),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_139),
.B(n_1),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_193),
.B(n_200),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_199),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_114),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_148),
.A2(n_51),
.B1(n_44),
.B2(n_4),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_101),
.B(n_44),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_137),
.C(n_133),
.Y(n_201)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_198),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_201),
.B(n_208),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_127),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_199),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_168),
.A2(n_117),
.B1(n_107),
.B2(n_131),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_220),
.B1(n_239),
.B2(n_134),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_167),
.A2(n_145),
.B1(n_131),
.B2(n_107),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_229),
.B1(n_175),
.B2(n_176),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_167),
.A2(n_145),
.B1(n_117),
.B2(n_135),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_188),
.A2(n_108),
.B(n_119),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_240),
.B(n_132),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_171),
.B(n_141),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_232),
.B(n_178),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_174),
.A2(n_135),
.B1(n_134),
.B2(n_127),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_190),
.A2(n_108),
.B(n_133),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_211),
.A2(n_170),
.B1(n_132),
.B2(n_169),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_177),
.C(n_193),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_265),
.C(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_191),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_247),
.Y(n_281)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_245),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_179),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_246),
.B(n_248),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_156),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_155),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_202),
.Y(n_249)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_251),
.A2(n_254),
.B1(n_255),
.B2(n_261),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_187),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_174),
.B1(n_197),
.B2(n_172),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_197),
.B1(n_185),
.B2(n_162),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_258),
.A2(n_271),
.B1(n_218),
.B2(n_207),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_203),
.B(n_235),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_259),
.A2(n_205),
.B(n_218),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_262),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_219),
.A2(n_186),
.B1(n_192),
.B2(n_141),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_163),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_214),
.Y(n_263)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_235),
.B(n_106),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_264),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_208),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_267),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_208),
.B(n_146),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_270),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_209),
.B(n_146),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_226),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_109),
.B1(n_125),
.B2(n_118),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_201),
.A2(n_208),
.B1(n_213),
.B2(n_230),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_208),
.A2(n_109),
.B1(n_180),
.B2(n_194),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_213),
.A2(n_152),
.B1(n_198),
.B2(n_182),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_106),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_214),
.Y(n_276)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_225),
.A3(n_226),
.B1(n_203),
.B2(n_224),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_295),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_268),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_240),
.C(n_223),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_296),
.C(n_300),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_254),
.A2(n_223),
.B1(n_205),
.B2(n_207),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_289),
.A2(n_305),
.B1(n_271),
.B2(n_256),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_248),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_291),
.B(n_292),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_294),
.A2(n_303),
.B1(n_261),
.B2(n_221),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_245),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_253),
.B(n_223),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_245),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_297),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_272),
.A2(n_267),
.B(n_253),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_270),
.B(n_253),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_233),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_258),
.A2(n_222),
.B1(n_234),
.B2(n_206),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_243),
.B(n_231),
.C(n_212),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_275),
.C(n_259),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_252),
.A2(n_222),
.B1(n_234),
.B2(n_212),
.Y(n_305)
);

AOI21x1_ASAP7_75t_SL g358 ( 
.A1(n_312),
.A2(n_314),
.B(n_316),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_243),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_319),
.C(n_322),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_307),
.A2(n_268),
.B(n_264),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_268),
.B(n_262),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_283),
.A2(n_251),
.B1(n_260),
.B2(n_269),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_317),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_342)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_244),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_323),
.Y(n_347)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_326),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_250),
.C(n_242),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_307),
.A2(n_273),
.B(n_246),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_327),
.A2(n_340),
.B(n_292),
.Y(n_356)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_330),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_281),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_331),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_249),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_302),
.A2(n_276),
.B1(n_263),
.B2(n_255),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_333),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_284),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_236),
.C(n_231),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_339),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_294),
.A2(n_234),
.B1(n_236),
.B2(n_221),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_303),
.A2(n_228),
.B1(n_238),
.B2(n_200),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_281),
.B(n_278),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_282),
.A2(n_228),
.B(n_238),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_317),
.A2(n_298),
.B1(n_289),
.B2(n_305),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_344),
.A2(n_360),
.B1(n_362),
.B2(n_314),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_335),
.B(n_301),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_346),
.A2(n_351),
.B1(n_361),
.B2(n_328),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_357),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_338),
.A2(n_279),
.B1(n_337),
.B2(n_308),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_308),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_354),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_356),
.A2(n_140),
.B(n_111),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_332),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_312),
.A2(n_288),
.B1(n_310),
.B2(n_279),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_324),
.B(n_310),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_316),
.A2(n_282),
.B1(n_299),
.B2(n_287),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_333),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_365),
.Y(n_375)
);

OA21x2_ASAP7_75t_L g365 ( 
.A1(n_330),
.A2(n_306),
.B(n_309),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_340),
.Y(n_366)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_366),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_318),
.A2(n_306),
.B(n_277),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_367),
.A2(n_327),
.B(n_334),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_331),
.C(n_318),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_373),
.C(n_374),
.Y(n_403)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_371),
.A2(n_386),
.B(n_356),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_322),
.C(n_313),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_329),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_341),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_357),
.A2(n_359),
.B1(n_353),
.B2(n_366),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_376),
.A2(n_384),
.B1(n_343),
.B2(n_355),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_377),
.A2(n_360),
.B(n_358),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_344),
.A2(n_306),
.B1(n_287),
.B2(n_285),
.Y(n_378)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_378),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_342),
.A2(n_319),
.B1(n_325),
.B2(n_290),
.Y(n_379)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_379),
.Y(n_395)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_380),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_309),
.B1(n_285),
.B2(n_290),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_342),
.A2(n_339),
.B1(n_140),
.B2(n_4),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_385),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_365),
.A2(n_359),
.B1(n_353),
.B2(n_364),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_347),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_111),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_350),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_2),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_390),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_362),
.A2(n_111),
.B1(n_12),
.B2(n_4),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g391 ( 
.A(n_373),
.B(n_358),
.CI(n_367),
.CON(n_391),
.SN(n_391)
);

FAx1_ASAP7_75t_SL g415 ( 
.A(n_391),
.B(n_400),
.CI(n_371),
.CON(n_415),
.SN(n_415)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_398),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_404),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_375),
.A2(n_361),
.B(n_365),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_406),
.Y(n_411)
);

FAx1_ASAP7_75t_SL g400 ( 
.A(n_377),
.B(n_363),
.CI(n_341),
.CON(n_400),
.SN(n_400)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_402),
.A2(n_345),
.B1(n_347),
.B2(n_5),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_403),
.B(n_387),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_343),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_379),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_408),
.B(n_388),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_409),
.B(n_412),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_401),
.A2(n_376),
.B1(n_372),
.B2(n_384),
.Y(n_410)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_403),
.B(n_383),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_422),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_370),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_414),
.B(n_416),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_393),
.C(n_395),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_370),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_392),
.A2(n_372),
.B1(n_375),
.B2(n_389),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_421),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_378),
.C(n_382),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_423),
.C(n_405),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_402),
.A2(n_390),
.B1(n_386),
.B2(n_355),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_345),
.C(n_63),
.Y(n_423)
);

FAx1_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_415),
.CI(n_400),
.CON(n_443),
.SN(n_443)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_395),
.C(n_396),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_431),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_433),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_392),
.C(n_398),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_411),
.A2(n_410),
.B(n_423),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_415),
.B(n_397),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_399),
.C(n_405),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_406),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_434),
.B(n_435),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_422),
.C(n_417),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_394),
.Y(n_437)
);

AO21x1_ASAP7_75t_L g450 ( 
.A1(n_437),
.A2(n_443),
.B(n_444),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_430),
.B(n_391),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_440),
.B(n_12),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_431),
.B(n_391),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_442),
.A2(n_447),
.B(n_12),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_394),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_421),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_436),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_446),
.B(n_424),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_427),
.A2(n_400),
.B(n_397),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_438),
.B(n_426),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_448),
.B(n_452),
.Y(n_458)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_449),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_SL g451 ( 
.A(n_441),
.B(n_436),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_451),
.A2(n_454),
.B(n_455),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_453),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_444),
.Y(n_454)
);

NAND4xp25_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_439),
.C(n_437),
.D(n_443),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_460),
.B(n_12),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_461),
.A2(n_463),
.B(n_457),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_458),
.B(n_5),
.C(n_11),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_462),
.A2(n_456),
.B(n_13),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_459),
.A2(n_11),
.B(n_13),
.Y(n_463)
);

OAI321xp33_ASAP7_75t_L g466 ( 
.A1(n_464),
.A2(n_465),
.A3(n_14),
.B1(n_15),
.B2(n_2),
.C(n_3),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_466),
.A2(n_15),
.B(n_3),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_467),
.A2(n_3),
.B(n_321),
.Y(n_468)
);


endmodule