module real_jpeg_21038_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_0),
.A2(n_35),
.B1(n_38),
.B2(n_56),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_56),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_24),
.B1(n_32),
.B2(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_2),
.A2(n_35),
.B1(n_38),
.B2(n_72),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_37),
.B(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_3),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_3),
.A2(n_12),
.B(n_23),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_28),
.B1(n_111),
.B2(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_3),
.B(n_65),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_25),
.Y(n_26)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_11),
.A2(n_35),
.B1(n_38),
.B2(n_48),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_48),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_12),
.A2(n_32),
.B(n_52),
.C(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_12),
.B(n_32),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_12),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_13),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_88),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_87),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_59),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_18),
.B(n_59),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.C(n_49),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_19),
.A2(n_20),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_31),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_27),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_22),
.B(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_25),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_26),
.B(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_26),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_28),
.B(n_101),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.A3(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_33),
.B1(n_36),
.B2(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_33),
.A2(n_54),
.B(n_101),
.C(n_102),
.Y(n_100)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_40),
.B(n_44),
.C(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_41),
.A2(n_42),
.B1(n_49),
.B2(n_50),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_57),
.B(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_53),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_51),
.A2(n_53),
.B1(n_55),
.B2(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_101),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_80),
.B2(n_81),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B(n_78),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_94),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_131),
.B(n_136),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_119),
.B(n_130),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_107),
.B(n_118),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_112),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_103),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_113),
.B(n_117),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_126),
.C(n_127),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.Y(n_136)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);


endmodule