module fake_jpeg_29875_n_528 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_528);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_55),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_1),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_70),
.Y(n_112)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_2),
.Y(n_70)
);

CKINVDCx9p33_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_2),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_74),
.B(n_89),
.Y(n_149)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_100),
.Y(n_138)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_28),
.B(n_3),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_22),
.A2(n_26),
.B(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_99),
.B(n_102),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_30),
.B(n_4),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_30),
.B(n_4),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_43),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_47),
.B1(n_40),
.B2(n_39),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_47),
.B1(n_40),
.B2(n_39),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_124),
.B(n_153),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_85),
.A2(n_40),
.B1(n_49),
.B2(n_29),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_126),
.A2(n_129),
.B1(n_156),
.B2(n_81),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_70),
.A2(n_37),
.B1(n_51),
.B2(n_22),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_74),
.B(n_37),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_157),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_54),
.A2(n_40),
.B1(n_49),
.B2(n_21),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_58),
.A2(n_51),
.B1(n_26),
.B2(n_33),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_161),
.A2(n_95),
.B1(n_38),
.B2(n_23),
.Y(n_214)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_112),
.A2(n_29),
.B1(n_27),
.B2(n_24),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_174),
.Y(n_257)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_166),
.A2(n_77),
.B1(n_29),
.B2(n_27),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_177),
.A2(n_188),
.B1(n_212),
.B2(n_217),
.Y(n_242)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_178),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_112),
.B(n_27),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_185),
.Y(n_237)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_21),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_181),
.B(n_183),
.Y(n_265)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_21),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_49),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_24),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_187),
.B(n_195),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_116),
.A2(n_24),
.B1(n_78),
.B2(n_94),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_189),
.Y(n_228)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_190),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_191),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_126),
.A2(n_42),
.B1(n_43),
.B2(n_38),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_192),
.B(n_218),
.Y(n_241)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_194),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_156),
.A2(n_82),
.B1(n_63),
.B2(n_92),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_205),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_131),
.B(n_87),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_197),
.B(n_165),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_199),
.Y(n_260)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_200),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_147),
.B(n_43),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_201),
.B(n_204),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_141),
.B(n_61),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_203),
.B(n_220),
.C(n_151),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_142),
.B(n_43),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_159),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_140),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_206),
.Y(n_259)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_208),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_151),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_211),
.Y(n_230)
);

BUFx8_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

INVx6_ASAP7_75t_SL g270 ( 
.A(n_210),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_144),
.B(n_43),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_123),
.A2(n_72),
.B1(n_68),
.B2(n_105),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_215),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_221),
.B1(n_132),
.B2(n_125),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_143),
.B(n_38),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_222),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_139),
.A2(n_42),
.B1(n_5),
.B2(n_6),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_113),
.B(n_4),
.C(n_5),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_118),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_133),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_225),
.Y(n_249)
);

INVx3_ASAP7_75t_SL g224 ( 
.A(n_122),
.Y(n_224)
);

INVx2_ASAP7_75t_R g271 ( 
.A(n_224),
.Y(n_271)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_107),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_132),
.Y(n_253)
);

OR2x2_ASAP7_75t_SL g232 ( 
.A(n_179),
.B(n_109),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_232),
.Y(n_282)
);

AND2x6_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_108),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_239),
.B(n_263),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_245),
.A2(n_224),
.B1(n_130),
.B2(n_165),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_266),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_258),
.Y(n_284)
);

NOR4xp25_ASAP7_75t_SL g256 ( 
.A(n_169),
.B(n_120),
.C(n_9),
.D(n_10),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_220),
.B(n_157),
.C(n_199),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_202),
.B(n_173),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_189),
.B(n_118),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_197),
.B(n_135),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_267),
.B(n_203),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_168),
.B(n_182),
.C(n_184),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_186),
.C(n_208),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_237),
.B(n_198),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_274),
.B(n_278),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_228),
.A2(n_195),
.B1(n_192),
.B2(n_203),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_275),
.A2(n_287),
.B1(n_288),
.B2(n_297),
.Y(n_315)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_277),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_243),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_281),
.B(n_283),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_249),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_234),
.Y(n_285)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_270),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_293),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_240),
.B1(n_242),
.B2(n_267),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_230),
.B(n_210),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_296),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_242),
.A2(n_170),
.B1(n_178),
.B2(n_193),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_290),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_269),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_291),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_271),
.A2(n_171),
.B1(n_191),
.B2(n_176),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_292),
.A2(n_268),
.B1(n_254),
.B2(n_190),
.Y(n_346)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_252),
.A2(n_175),
.B1(n_194),
.B2(n_135),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_252),
.A2(n_233),
.B(n_263),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_298),
.A2(n_312),
.B(n_314),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_237),
.B(n_200),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_302),
.Y(n_330)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_264),
.Y(n_300)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_300),
.Y(n_341)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_301),
.Y(n_349)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_305),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_269),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_304),
.Y(n_347)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_248),
.B(n_210),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_307),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_174),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_308),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_239),
.A2(n_125),
.B1(n_134),
.B2(n_130),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_265),
.B1(n_247),
.B2(n_259),
.Y(n_317)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_250),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_310),
.Y(n_345)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_218),
.B1(n_261),
.B2(n_246),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_256),
.A2(n_206),
.B1(n_213),
.B2(n_180),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_273),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_271),
.A2(n_207),
.B(n_222),
.Y(n_314)
);

AO21x2_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_271),
.B(n_241),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_316),
.A2(n_268),
.B(n_262),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_317),
.A2(n_322),
.B1(n_344),
.B2(n_297),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_240),
.B1(n_232),
.B2(n_247),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_323),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_272),
.C(n_257),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_331),
.C(n_337),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_257),
.C(n_246),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_312),
.B(n_307),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_335),
.A2(n_342),
.B(n_255),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_270),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_282),
.A2(n_259),
.B(n_262),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_338),
.A2(n_342),
.B(n_330),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_343),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_282),
.A2(n_259),
.B(n_262),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_299),
.B(n_273),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_274),
.A2(n_255),
.B1(n_225),
.B2(n_119),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_346),
.A2(n_286),
.B1(n_288),
.B2(n_275),
.Y(n_356)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_351),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_319),
.B(n_280),
.Y(n_354)
);

AOI21xp33_ASAP7_75t_L g391 ( 
.A1(n_354),
.A2(n_343),
.B(n_338),
.Y(n_391)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_355),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_356),
.A2(n_361),
.B1(n_381),
.B2(n_328),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_321),
.A2(n_311),
.B1(n_283),
.B2(n_296),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_357),
.A2(n_359),
.B1(n_368),
.B2(n_369),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_348),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_358),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_321),
.A2(n_280),
.B1(n_281),
.B2(n_309),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_326),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_360),
.Y(n_404)
);

OAI22x1_ASAP7_75t_SL g361 ( 
.A1(n_316),
.A2(n_293),
.B1(n_284),
.B2(n_292),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_362),
.A2(n_367),
.B1(n_370),
.B2(n_376),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_289),
.Y(n_363)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_363),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_284),
.Y(n_364)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_320),
.Y(n_365)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_365),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_329),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_380),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_322),
.A2(n_293),
.B1(n_278),
.B2(n_313),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_335),
.A2(n_306),
.B1(n_305),
.B2(n_303),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_336),
.A2(n_286),
.B1(n_291),
.B2(n_304),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_315),
.A2(n_294),
.B1(n_302),
.B2(n_300),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_319),
.B(n_261),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_373),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_317),
.B(n_301),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_324),
.B(n_279),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_378),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_315),
.A2(n_295),
.B1(n_285),
.B2(n_255),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_377),
.A2(n_382),
.B(n_383),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_329),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_336),
.A2(n_310),
.B1(n_308),
.B2(n_254),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_379),
.A2(n_345),
.B1(n_334),
.B2(n_341),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_330),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_332),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_327),
.C(n_339),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_398),
.C(n_399),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_386),
.A2(n_400),
.B1(n_403),
.B2(n_371),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_331),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_390),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_337),
.Y(n_390)
);

OAI21xp33_ASAP7_75t_SL g423 ( 
.A1(n_391),
.A2(n_379),
.B(n_374),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_383),
.A2(n_316),
.B(n_328),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_392),
.A2(n_397),
.B(n_369),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_362),
.A2(n_346),
.B1(n_316),
.B2(n_347),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_393),
.A2(n_394),
.B1(n_406),
.B2(n_356),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_370),
.A2(n_316),
.B1(n_344),
.B2(n_350),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_341),
.B(n_332),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_357),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_367),
.B(n_359),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_368),
.B(n_364),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_402),
.C(n_398),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_334),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_361),
.A2(n_345),
.B1(n_333),
.B2(n_349),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_376),
.A2(n_345),
.B1(n_333),
.B2(n_349),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_358),
.A2(n_340),
.B1(n_134),
.B2(n_119),
.Y(n_408)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

A2O1A1Ixp33_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_354),
.B(n_380),
.C(n_363),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_414),
.A2(n_392),
.B(n_409),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_412),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_421),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_419),
.Y(n_445)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_412),
.Y(n_418)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

XNOR2x1_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_363),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_432),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_360),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_351),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_430),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_423),
.A2(n_388),
.B1(n_384),
.B2(n_400),
.Y(n_443)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_410),
.Y(n_424)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_424),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_385),
.B(n_366),
.C(n_378),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_427),
.C(n_431),
.Y(n_458)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_389),
.B(n_381),
.C(n_365),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_428),
.A2(n_434),
.B1(n_393),
.B2(n_406),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_355),
.Y(n_429)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_397),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_401),
.C(n_402),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_413),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_433),
.A2(n_387),
.B1(n_397),
.B2(n_411),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_403),
.A2(n_375),
.B1(n_235),
.B2(n_244),
.Y(n_434)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_407),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_436),
.B(n_437),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_413),
.Y(n_437)
);

OAI21xp33_ASAP7_75t_L g439 ( 
.A1(n_405),
.A2(n_375),
.B(n_235),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_394),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_428),
.Y(n_464)
);

XNOR2x1_ASAP7_75t_L g468 ( 
.A(n_446),
.B(n_431),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_388),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_453),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_450),
.A2(n_429),
.B1(n_236),
.B2(n_107),
.Y(n_474)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_452),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_396),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_396),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_457),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_418),
.A2(n_426),
.B1(n_424),
.B2(n_387),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_455),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_415),
.B(n_409),
.Y(n_457)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_459),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_425),
.B(n_244),
.C(n_236),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_417),
.C(n_419),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_457),
.B(n_447),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_463),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_427),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_468),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_448),
.B(n_436),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_466),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_456),
.A2(n_438),
.B1(n_432),
.B2(n_437),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_440),
.Y(n_467)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_441),
.A2(n_444),
.B1(n_451),
.B2(n_446),
.Y(n_471)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_471),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_475),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_443),
.A2(n_434),
.B1(n_420),
.B2(n_414),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_473),
.A2(n_470),
.B(n_440),
.Y(n_478)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_474),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_236),
.C(n_9),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_477),
.B(n_442),
.C(n_468),
.Y(n_479)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_478),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_479),
.B(n_484),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_461),
.A2(n_449),
.B1(n_453),
.B2(n_452),
.Y(n_480)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_461),
.A2(n_455),
.B1(n_459),
.B2(n_445),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_488),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_477),
.A2(n_460),
.B(n_458),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_486),
.B(n_16),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_445),
.C(n_442),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_491),
.C(n_472),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_476),
.A2(n_236),
.B(n_11),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_16),
.C(n_11),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_490),
.A2(n_469),
.B1(n_464),
.B2(n_473),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_495),
.A2(n_498),
.B1(n_480),
.B2(n_482),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_496),
.B(n_504),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_489),
.A2(n_474),
.B1(n_12),
.B2(n_13),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_481),
.B(n_7),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_500),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_7),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_492),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_12),
.C(n_13),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_491),
.C(n_487),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_479),
.B(n_12),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_483),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_506),
.Y(n_514)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_494),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_507),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.Y(n_513)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_502),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_512),
.A2(n_493),
.B(n_497),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_515),
.B(n_511),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_SL g516 ( 
.A(n_508),
.B(n_496),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_516),
.A2(n_514),
.B(n_513),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_510),
.A2(n_503),
.B(n_483),
.Y(n_517)
);

AOI21xp33_ASAP7_75t_L g518 ( 
.A1(n_517),
.A2(n_506),
.B(n_509),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_518),
.A2(n_520),
.B(n_505),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_519),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_498),
.C(n_14),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_522),
.C(n_14),
.Y(n_524)
);

OAI21xp33_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_13),
.B(n_14),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_13),
.B1(n_15),
.B2(n_209),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_15),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_15),
.Y(n_528)
);


endmodule