module fake_netlist_1_1110_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_0), .B(n_7), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
BUFx8_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_4), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
INVxp67_ASAP7_75t_SL g20 ( .A(n_16), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_15), .B(n_2), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_15), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_12), .B(n_5), .Y(n_24) );
BUFx6f_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_19), .A2(n_13), .B1(n_11), .B2(n_16), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_20), .A2(n_17), .B1(n_5), .B2(n_10), .Y(n_27) );
AND2x2_ASAP7_75t_SL g28 ( .A(n_21), .B(n_17), .Y(n_28) );
NAND4xp25_ASAP7_75t_L g29 ( .A(n_26), .B(n_24), .C(n_22), .D(n_23), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_23), .Y(n_30) );
BUFx3_ASAP7_75t_L g31 ( .A(n_25), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_28), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_29), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_32), .B(n_23), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_34), .B(n_32), .Y(n_36) );
AOI321xp33_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_33), .A3(n_23), .B1(n_31), .B2(n_8), .C(n_25), .Y(n_37) );
INVx2_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_37), .B(n_25), .Y(n_39) );
NAND2xp5_ASAP7_75t_L g40 ( .A(n_38), .B(n_39), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_40), .Y(n_41) );
endmodule