module fake_ibex_1938_n_3796 (n_151, n_85, n_599, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_421, n_738, n_475, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_768, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_762, n_410, n_308, n_675, n_463, n_624, n_706, n_411, n_135, n_520, n_684, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_728, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_3796);

input n_151;
input n_85;
input n_599;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_738;
input n_475;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_768;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_684;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_3796;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_3750;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3395;
wire n_3242;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_2924;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_784;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_1969;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_3317;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_3416;
wire n_1031;
wire n_2962;
wire n_2879;
wire n_2958;
wire n_3694;
wire n_3147;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3660;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_3626;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_2252;
wire n_1982;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_2294;
wire n_1977;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2991;
wire n_2234;
wire n_847;
wire n_2699;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1395;
wire n_998;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2654;
wire n_2463;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_2974;
wire n_871;
wire n_2990;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2923;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_991;
wire n_1331;
wire n_1223;
wire n_961;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1946;
wire n_1726;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3333;
wire n_3096;
wire n_839;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2251;
wire n_2012;
wire n_3512;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_1455;
wire n_804;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3619;
wire n_3349;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2675;
wire n_786;
wire n_2348;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_3465;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_3066;
wire n_2714;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_1542;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1547;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3561;
wire n_2381;
wire n_2313;
wire n_3368;
wire n_956;
wire n_3586;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3360;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_3227;
wire n_2938;
wire n_1438;
wire n_3774;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_3380;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3557;
wire n_3596;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3483;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3622;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_2148;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3189;
wire n_3052;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2673;
wire n_2676;
wire n_921;
wire n_2430;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_3180;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

INVx1_ASAP7_75t_L g769 ( 
.A(n_623),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_341),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_712),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_630),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_214),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_8),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_327),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_314),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_284),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_298),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_646),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_312),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_436),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_358),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_738),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_389),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_19),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_137),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_528),
.Y(n_787)
);

BUFx8_ASAP7_75t_SL g788 ( 
.A(n_14),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_487),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_381),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_431),
.Y(n_791)
);

BUFx5_ASAP7_75t_L g792 ( 
.A(n_583),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_288),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_258),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_225),
.Y(n_795)
);

NOR2xp67_ASAP7_75t_L g796 ( 
.A(n_391),
.B(n_60),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_476),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_614),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_710),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_546),
.Y(n_800)
);

BUFx10_ASAP7_75t_L g801 ( 
.A(n_95),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_102),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_15),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_327),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_356),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_146),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_525),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_241),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_50),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_293),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_266),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_569),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_15),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_438),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_324),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_672),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_450),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_22),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_740),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_200),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_266),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_588),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_199),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_411),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_669),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_729),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_57),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_740),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_547),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_117),
.Y(n_830)
);

CKINVDCx14_ASAP7_75t_R g831 ( 
.A(n_104),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_7),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_92),
.Y(n_833)
);

BUFx8_ASAP7_75t_SL g834 ( 
.A(n_743),
.Y(n_834)
);

XOR2xp5_ASAP7_75t_L g835 ( 
.A(n_51),
.B(n_571),
.Y(n_835)
);

CKINVDCx14_ASAP7_75t_R g836 ( 
.A(n_491),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_403),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_508),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_689),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_249),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_219),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_77),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_264),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_368),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_243),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_755),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_283),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_505),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_515),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_18),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_663),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_510),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_160),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_498),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_390),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_350),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_137),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_399),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_344),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_697),
.Y(n_860)
);

BUFx10_ASAP7_75t_L g861 ( 
.A(n_240),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_414),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_L g863 ( 
.A(n_730),
.B(n_602),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_608),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_661),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_269),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_218),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_642),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_572),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_165),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_768),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_759),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_357),
.Y(n_873)
);

CKINVDCx16_ASAP7_75t_R g874 ( 
.A(n_372),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_87),
.Y(n_875)
);

INVx1_ASAP7_75t_SL g876 ( 
.A(n_556),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_173),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_370),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_447),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_208),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_523),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_396),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_718),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_428),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_50),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_573),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_473),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_763),
.Y(n_888)
);

INVxp33_ASAP7_75t_SL g889 ( 
.A(n_227),
.Y(n_889)
);

BUFx5_ASAP7_75t_L g890 ( 
.A(n_422),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_681),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_319),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_105),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_9),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_564),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_120),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_230),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_685),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_16),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_101),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_258),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_213),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_238),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_298),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_485),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_641),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_697),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_92),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_350),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_186),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_353),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_607),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_730),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_3),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_738),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_453),
.Y(n_916)
);

INVxp67_ASAP7_75t_SL g917 ( 
.A(n_3),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_590),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_270),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_180),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_273),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_480),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_145),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_191),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_675),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_33),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_600),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_472),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_680),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_270),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_54),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_68),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_180),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_254),
.Y(n_934)
);

CKINVDCx16_ASAP7_75t_R g935 ( 
.A(n_545),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_408),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_361),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_178),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_698),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_677),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_121),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_565),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_491),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_362),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_115),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_651),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_477),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_293),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_705),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_156),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_304),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_23),
.Y(n_952)
);

NOR2xp67_ASAP7_75t_L g953 ( 
.A(n_310),
.B(n_76),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_177),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_94),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_528),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_239),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_760),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_171),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_331),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_401),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_69),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_186),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_360),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_456),
.Y(n_965)
);

CKINVDCx16_ASAP7_75t_R g966 ( 
.A(n_607),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_107),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_619),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_750),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_105),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_317),
.Y(n_971)
);

BUFx8_ASAP7_75t_SL g972 ( 
.A(n_96),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_524),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_222),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_369),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_223),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_272),
.Y(n_977)
);

BUFx8_ASAP7_75t_SL g978 ( 
.A(n_499),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_393),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_118),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_685),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_359),
.Y(n_982)
);

NOR2xp67_ASAP7_75t_L g983 ( 
.A(n_505),
.B(n_160),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_280),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_69),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_353),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_478),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_236),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_242),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_278),
.Y(n_990)
);

BUFx5_ASAP7_75t_L g991 ( 
.A(n_382),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_322),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_572),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_378),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_242),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_68),
.B(n_704),
.Y(n_996)
);

CKINVDCx16_ASAP7_75t_R g997 ( 
.A(n_9),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_296),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_378),
.Y(n_999)
);

BUFx8_ASAP7_75t_SL g1000 ( 
.A(n_384),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_38),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_451),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_382),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_723),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_38),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_111),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_518),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_511),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_500),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_640),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_486),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_537),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_536),
.B(n_303),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_714),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_337),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_578),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_532),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_739),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_19),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_187),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_184),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_29),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_442),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_74),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_82),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_446),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_650),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_489),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_108),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_116),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_713),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_404),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_495),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_597),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_174),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_72),
.Y(n_1036)
);

CKINVDCx16_ASAP7_75t_R g1037 ( 
.A(n_558),
.Y(n_1037)
);

INVxp33_ASAP7_75t_SL g1038 ( 
.A(n_564),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_762),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_218),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_486),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_688),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_676),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_273),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_533),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_732),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_43),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_635),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_192),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_676),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_479),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_21),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_724),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_254),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_765),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_448),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_169),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_L g1058 ( 
.A(n_488),
.B(n_395),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_720),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_367),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_498),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_467),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_745),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_220),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_648),
.Y(n_1065)
);

BUFx5_ASAP7_75t_L g1066 ( 
.A(n_597),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_115),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_703),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_540),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_271),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_26),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_368),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_250),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_229),
.Y(n_1074)
);

BUFx10_ASAP7_75t_L g1075 ( 
.A(n_244),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_269),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_93),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_548),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_130),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_508),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_415),
.B(n_323),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_544),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_331),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_496),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_406),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_724),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_513),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_318),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_277),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_672),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_519),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_537),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_683),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_150),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_543),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_358),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_260),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_548),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_526),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_11),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_557),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_253),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_577),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_157),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_340),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_727),
.Y(n_1106)
);

CKINVDCx16_ASAP7_75t_R g1107 ( 
.A(n_312),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_294),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_451),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_438),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_392),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_406),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_428),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_699),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_409),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_453),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_340),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_601),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_404),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_557),
.Y(n_1120)
);

INVxp67_ASAP7_75t_SL g1121 ( 
.A(n_124),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_550),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_370),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_104),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_444),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_305),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_226),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_133),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_629),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_164),
.Y(n_1130)
);

BUFx10_ASAP7_75t_L g1131 ( 
.A(n_464),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_163),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_263),
.Y(n_1133)
);

INVxp33_ASAP7_75t_SL g1134 ( 
.A(n_52),
.Y(n_1134)
);

XNOR2xp5_ASAP7_75t_L g1135 ( 
.A(n_278),
.B(n_535),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_256),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_10),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_197),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_11),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_401),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_29),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_764),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_113),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_461),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_420),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_387),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_244),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_17),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_247),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_155),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_460),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_512),
.Y(n_1152)
);

CKINVDCx16_ASAP7_75t_R g1153 ( 
.A(n_169),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_656),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_58),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_281),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_262),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_543),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_302),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_355),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_587),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_419),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_345),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_189),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_464),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_121),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_253),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_680),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_656),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_177),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_59),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_566),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_544),
.Y(n_1173)
);

NOR2xp67_ASAP7_75t_L g1174 ( 
.A(n_496),
.B(n_755),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_364),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_398),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_326),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_752),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_658),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_658),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_471),
.Y(n_1181)
);

CKINVDCx16_ASAP7_75t_R g1182 ( 
.A(n_25),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_666),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_230),
.B(n_700),
.Y(n_1184)
);

NOR2xp67_ASAP7_75t_L g1185 ( 
.A(n_112),
.B(n_67),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_772),
.A2(n_0),
.B(n_1),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_831),
.Y(n_1187)
);

BUFx8_ASAP7_75t_L g1188 ( 
.A(n_906),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_831),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_783),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_836),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_792),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_792),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_801),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_792),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_783),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_770),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_836),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_783),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_849),
.Y(n_1200)
);

BUFx8_ASAP7_75t_L g1201 ( 
.A(n_922),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_788),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_792),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_770),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_849),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_963),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_963),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_963),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_849),
.Y(n_1209)
);

BUFx12f_ASAP7_75t_L g1210 ( 
.A(n_801),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_792),
.Y(n_1211)
);

INVxp33_ASAP7_75t_SL g1212 ( 
.A(n_799),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_792),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1046),
.B(n_2),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_788),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_849),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_990),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_792),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1055),
.B(n_3),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_990),
.A2(n_4),
.B(n_5),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_890),
.Y(n_1221)
);

OAI22x1_ASAP7_75t_R g1222 ( 
.A1(n_781),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_990),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_772),
.A2(n_784),
.B(n_773),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1173),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1173),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_914),
.A2(n_935),
.B1(n_966),
.B2(n_874),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1173),
.B(n_4),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_858),
.Y(n_1229)
);

AND2x6_ASAP7_75t_L g1230 ( 
.A(n_782),
.B(n_5),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_970),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1065),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_773),
.A2(n_6),
.B(n_761),
.Y(n_1233)
);

AOI22x1_ASAP7_75t_SL g1234 ( 
.A1(n_781),
.A2(n_6),
.B1(n_8),
.B2(n_7),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_786),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_970),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_890),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_858),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1015),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_782),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1015),
.B(n_12),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1167),
.B(n_12),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1073),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_858),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_890),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_890),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_890),
.Y(n_1247)
);

AND2x6_ASAP7_75t_L g1248 ( 
.A(n_828),
.B(n_13),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1073),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_817),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_828),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_829),
.Y(n_1252)
);

INVx5_ASAP7_75t_L g1253 ( 
.A(n_858),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_784),
.A2(n_13),
.B(n_14),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_889),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_870),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_829),
.Y(n_1257)
);

AOI22x1_ASAP7_75t_SL g1258 ( 
.A1(n_786),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_834),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_869),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_889),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_997),
.A2(n_760),
.B1(n_761),
.B2(n_758),
.Y(n_1262)
);

INVx5_ASAP7_75t_L g1263 ( 
.A(n_870),
.Y(n_1263)
);

CKINVDCx6p67_ASAP7_75t_R g1264 ( 
.A(n_801),
.Y(n_1264)
);

AOI22x1_ASAP7_75t_SL g1265 ( 
.A1(n_830),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_869),
.B(n_27),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1038),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_939),
.Y(n_1268)
);

INVx6_ASAP7_75t_L g1269 ( 
.A(n_851),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1172),
.B(n_30),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_939),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_834),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_913),
.Y(n_1273)
);

BUFx8_ASAP7_75t_SL g1274 ( 
.A(n_972),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_956),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_890),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_890),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_991),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_870),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_991),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_SL g1281 ( 
.A1(n_830),
.A2(n_32),
.B1(n_28),
.B2(n_31),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_991),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_991),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_967),
.B(n_32),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_952),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_952),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_991),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_851),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_964),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_964),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_870),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_851),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1002),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1208),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1224),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1214),
.B(n_1103),
.C(n_947),
.Y(n_1296)
);

NAND3xp33_ASAP7_75t_L g1297 ( 
.A(n_1219),
.B(n_1270),
.C(n_1242),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1228),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1208),
.B(n_1038),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1228),
.B(n_991),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1230),
.A2(n_917),
.B1(n_777),
.B2(n_778),
.Y(n_1301)
);

NOR3xp33_ASAP7_75t_L g1302 ( 
.A(n_1262),
.B(n_1107),
.C(n_1037),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1224),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1197),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1192),
.B(n_991),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1200),
.Y(n_1306)
);

AND2x2_ASAP7_75t_SL g1307 ( 
.A(n_1266),
.B(n_1013),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1226),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1226),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1187),
.B(n_1182),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1197),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1204),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1192),
.B(n_1066),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1224),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1269),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1241),
.Y(n_1316)
);

NAND2xp33_ASAP7_75t_L g1317 ( 
.A(n_1230),
.B(n_1066),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1241),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1288),
.B(n_1134),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1217),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1288),
.B(n_806),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1204),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1266),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1200),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1240),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1193),
.B(n_1066),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1212),
.A2(n_1232),
.B1(n_1227),
.B2(n_1275),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1269),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1212),
.A2(n_1134),
.B1(n_1153),
.B2(n_807),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1231),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1273),
.B(n_861),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1193),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1195),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1195),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1269),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1203),
.B(n_1066),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1292),
.B(n_806),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1264),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1257),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1200),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1236),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1239),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1194),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1243),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1200),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_L g1346 ( 
.A(n_1232),
.B(n_1139),
.C(n_1062),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1203),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1211),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1198),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1257),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1211),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1249),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1213),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1194),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1274),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1273),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1218),
.B(n_1066),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1210),
.B(n_796),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1218),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1230),
.A2(n_779),
.B1(n_780),
.B2(n_769),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1221),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_SL g1362 ( 
.A(n_1230),
.B(n_1210),
.Y(n_1362)
);

OR2x6_ASAP7_75t_L g1363 ( 
.A(n_1281),
.B(n_863),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1189),
.A2(n_850),
.B1(n_852),
.B2(n_832),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1221),
.B(n_1066),
.Y(n_1365)
);

INVx8_ASAP7_75t_L g1366 ( 
.A(n_1198),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1271),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1289),
.Y(n_1368)
);

INVx5_ASAP7_75t_L g1369 ( 
.A(n_1248),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1289),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1293),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1196),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1196),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_SL g1374 ( 
.A(n_1250),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1207),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1207),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1223),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1223),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1190),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1199),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_SL g1381 ( 
.A(n_1250),
.Y(n_1381)
);

NOR2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1215),
.B(n_807),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1237),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1206),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1225),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1253),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1251),
.Y(n_1387)
);

INVxp67_ASAP7_75t_SL g1388 ( 
.A(n_1186),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1292),
.B(n_808),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1252),
.B(n_1290),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1260),
.Y(n_1391)
);

CKINVDCx6p67_ASAP7_75t_R g1392 ( 
.A(n_1259),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1268),
.B(n_771),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1253),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1237),
.B(n_1066),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1215),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1285),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1286),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1253),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1284),
.B(n_809),
.C(n_808),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1245),
.B(n_775),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1188),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1248),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1254),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1263),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1222),
.B(n_1220),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1188),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1245),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1274),
.Y(n_1409)
);

NAND3xp33_ASAP7_75t_L g1410 ( 
.A(n_1186),
.B(n_1191),
.C(n_1233),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1246),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1247),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1247),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1276),
.B(n_809),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1276),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1277),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1278),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1278),
.B(n_810),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1280),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1272),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1282),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1282),
.B(n_776),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1283),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1248),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1283),
.B(n_940),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1287),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1272),
.B(n_861),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1287),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1205),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1205),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1209),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1209),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1209),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1233),
.Y(n_1434)
);

OAI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1255),
.A2(n_850),
.B1(n_852),
.B2(n_832),
.Y(n_1435)
);

INVxp33_ASAP7_75t_L g1436 ( 
.A(n_1235),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1201),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1216),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1216),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1291),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1229),
.B(n_785),
.Y(n_1441)
);

NAND2xp33_ASAP7_75t_L g1442 ( 
.A(n_1229),
.B(n_1118),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1229),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1238),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1238),
.B(n_812),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1202),
.B(n_861),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1259),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1238),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1238),
.B(n_787),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1244),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1235),
.B(n_955),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1201),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1244),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1261),
.B(n_955),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1267),
.Y(n_1455)
);

INVxp33_ASAP7_75t_SL g1456 ( 
.A(n_1234),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1244),
.B(n_955),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1256),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1291),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1256),
.B(n_1118),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1256),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1256),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1279),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1279),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1350),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1294),
.B(n_813),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1308),
.B(n_816),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1315),
.B(n_789),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1309),
.B(n_819),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1350),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1298),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1298),
.B(n_819),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1356),
.A2(n_1081),
.B(n_1184),
.C(n_790),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1373),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1373),
.B(n_821),
.Y(n_1475)
);

NAND2xp33_ASAP7_75t_L g1476 ( 
.A(n_1369),
.B(n_1130),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1316),
.B(n_1002),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1410),
.B(n_996),
.C(n_822),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1362),
.B(n_1130),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1377),
.B(n_821),
.Y(n_1480)
);

NOR2x1_ASAP7_75t_L g1481 ( 
.A(n_1400),
.B(n_1007),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1320),
.B(n_822),
.Y(n_1482)
);

AND2x2_ASAP7_75t_SL g1483 ( 
.A(n_1437),
.B(n_1356),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1330),
.Y(n_1484)
);

NAND2xp33_ASAP7_75t_L g1485 ( 
.A(n_1369),
.B(n_1142),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1341),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1424),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1342),
.Y(n_1488)
);

O2A1O1Ixp5_ASAP7_75t_L g1489 ( 
.A1(n_1388),
.A2(n_844),
.B(n_848),
.C(n_811),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1318),
.B(n_824),
.Y(n_1490)
);

O2A1O1Ixp5_ASAP7_75t_L g1491 ( 
.A1(n_1388),
.A2(n_848),
.B(n_886),
.C(n_844),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1344),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1331),
.B(n_825),
.Y(n_1493)
);

AOI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1364),
.A2(n_827),
.B1(n_833),
.B2(n_826),
.C(n_825),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1321),
.B(n_826),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1406),
.A2(n_1121),
.B1(n_833),
.B2(n_976),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_SL g1497 ( 
.A(n_1403),
.B(n_972),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1337),
.B(n_827),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1352),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1389),
.B(n_976),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1372),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1304),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1299),
.B(n_980),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1311),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1299),
.B(n_1323),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1307),
.A2(n_1024),
.B1(n_1128),
.B2(n_1007),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1406),
.A2(n_1101),
.B1(n_1136),
.B2(n_980),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1328),
.B(n_953),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1307),
.A2(n_1128),
.B1(n_1148),
.B2(n_1024),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1375),
.Y(n_1510)
);

CKINVDCx11_ASAP7_75t_R g1511 ( 
.A(n_1392),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1319),
.B(n_791),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1376),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1414),
.B(n_1418),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1319),
.B(n_793),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1378),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1406),
.B(n_1258),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1301),
.A2(n_884),
.B1(n_907),
.B2(n_897),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1457),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1312),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1343),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1401),
.B(n_1101),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1401),
.B(n_1136),
.Y(n_1523)
);

CKINVDCx14_ASAP7_75t_R g1524 ( 
.A(n_1355),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1422),
.B(n_1137),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1328),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1354),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1322),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1338),
.B(n_835),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1379),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1335),
.B(n_983),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1380),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1325),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1385),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1310),
.B(n_1075),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1422),
.B(n_1137),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1297),
.B(n_797),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1301),
.A2(n_1455),
.B1(n_1302),
.B2(n_1360),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1384),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1374),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1339),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1387),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1397),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1335),
.B(n_800),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1368),
.Y(n_1545)
);

OR2x6_ASAP7_75t_L g1546 ( 
.A(n_1402),
.B(n_1407),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1391),
.B(n_1141),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1393),
.B(n_1141),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1393),
.B(n_1143),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1300),
.B(n_1143),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1300),
.B(n_1144),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1398),
.B(n_1144),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1390),
.B(n_1145),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1445),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1367),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1452),
.B(n_1145),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1370),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1390),
.B(n_1148),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1371),
.B(n_1162),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1296),
.B(n_892),
.Y(n_1560)
);

NAND2xp33_ASAP7_75t_L g1561 ( 
.A(n_1434),
.B(n_804),
.Y(n_1561)
);

AOI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1302),
.A2(n_794),
.B1(n_798),
.B2(n_795),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1404),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1346),
.B(n_1349),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1441),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1295),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1441),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1449),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1295),
.Y(n_1569)
);

NOR3xp33_ASAP7_75t_L g1570 ( 
.A(n_1435),
.B(n_846),
.C(n_774),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1454),
.A2(n_803),
.B1(n_805),
.B2(n_802),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1374),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1381),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1449),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1303),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1303),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1366),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1423),
.B(n_1314),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1363),
.A2(n_815),
.B(n_818),
.C(n_814),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1317),
.A2(n_1279),
.B(n_950),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1366),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1423),
.B(n_837),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1317),
.A2(n_823),
.B1(n_838),
.B2(n_820),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1427),
.B(n_899),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1446),
.B(n_950),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1366),
.B(n_1265),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1464),
.Y(n_1587)
);

NOR3xp33_ASAP7_75t_L g1588 ( 
.A(n_1435),
.B(n_912),
.C(n_876),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1329),
.B(n_840),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1408),
.B(n_961),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1464),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1412),
.B(n_841),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1327),
.B(n_961),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1415),
.B(n_842),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1386),
.Y(n_1595)
);

OR2x6_ASAP7_75t_L g1596 ( 
.A(n_1451),
.B(n_978),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1396),
.B(n_982),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1416),
.B(n_982),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1358),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1382),
.B(n_1058),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1394),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1358),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1305),
.A2(n_1279),
.B(n_1008),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1417),
.B(n_843),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1420),
.B(n_1436),
.Y(n_1605)
);

OAI22x1_ASAP7_75t_SL g1606 ( 
.A1(n_1456),
.A2(n_897),
.B1(n_907),
.B2(n_884),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1436),
.B(n_1364),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1381),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1332),
.B(n_845),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1358),
.B(n_1174),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1399),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1333),
.B(n_1006),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1334),
.B(n_1008),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1405),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1347),
.A2(n_847),
.B1(n_855),
.B2(n_839),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1348),
.B(n_862),
.C(n_859),
.Y(n_1616)
);

O2A1O1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1363),
.A2(n_867),
.B(n_871),
.C(n_864),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1351),
.A2(n_1359),
.B1(n_1361),
.B2(n_1353),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1458),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1351),
.B(n_1020),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1447),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1363),
.B(n_1075),
.Y(n_1622)
);

O2A1O1Ixp5_ASAP7_75t_L g1623 ( 
.A1(n_1305),
.A2(n_1022),
.B(n_1029),
.C(n_1020),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1353),
.B(n_1022),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1313),
.A2(n_875),
.B1(n_877),
.B2(n_872),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1359),
.B(n_853),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1313),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_SL g1628 ( 
.A(n_1361),
.B(n_1029),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1383),
.A2(n_879),
.B1(n_881),
.B2(n_878),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1326),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1383),
.Y(n_1631)
);

INVx8_ASAP7_75t_L g1632 ( 
.A(n_1409),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1411),
.B(n_854),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1411),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1413),
.B(n_856),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1326),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1413),
.B(n_1032),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1336),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1419),
.B(n_857),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1357),
.A2(n_885),
.B1(n_888),
.B2(n_882),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1419),
.B(n_860),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1421),
.Y(n_1642)
);

OR2x2_ASAP7_75t_SL g1643 ( 
.A(n_1421),
.B(n_978),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1426),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1365),
.B(n_865),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1428),
.Y(n_1646)
);

NOR2xp67_ASAP7_75t_L g1647 ( 
.A(n_1395),
.B(n_35),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1428),
.B(n_866),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1395),
.A2(n_943),
.B1(n_965),
.B2(n_929),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1425),
.B(n_868),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1425),
.A2(n_894),
.B(n_893),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1461),
.B(n_873),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1458),
.Y(n_1653)
);

BUFx5_ASAP7_75t_L g1654 ( 
.A(n_1463),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1463),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1460),
.B(n_880),
.Y(n_1656)
);

INVx8_ASAP7_75t_L g1657 ( 
.A(n_1306),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1306),
.Y(n_1658)
);

O2A1O1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1460),
.A2(n_900),
.B(n_901),
.C(n_896),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1442),
.A2(n_903),
.B1(n_904),
.B2(n_902),
.Y(n_1660)
);

INVx8_ASAP7_75t_L g1661 ( 
.A(n_1306),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1306),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1442),
.B(n_883),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1440),
.B(n_887),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1448),
.B(n_891),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1459),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1438),
.B(n_895),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1324),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1439),
.B(n_898),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1450),
.B(n_911),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1453),
.A2(n_908),
.B1(n_909),
.B2(n_905),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1462),
.B(n_915),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1429),
.Y(n_1673)
);

INVx8_ASAP7_75t_L g1674 ( 
.A(n_1324),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1430),
.B(n_921),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1324),
.B(n_923),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1340),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1430),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1345),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1431),
.B(n_924),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1432),
.B(n_925),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1432),
.B(n_926),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1345),
.B(n_928),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1433),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1433),
.B(n_931),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1345),
.B(n_932),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1443),
.Y(n_1687)
);

NOR3xp33_ASAP7_75t_L g1688 ( 
.A(n_1443),
.B(n_1098),
.C(n_1005),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1563),
.A2(n_1444),
.B(n_1111),
.Y(n_1689)
);

OR2x6_ASAP7_75t_L g1690 ( 
.A(n_1632),
.B(n_1185),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1505),
.B(n_936),
.Y(n_1691)
);

A2O1A1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1514),
.A2(n_916),
.B(n_918),
.C(n_910),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1471),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1484),
.B(n_938),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1577),
.B(n_919),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1576),
.Y(n_1696)
);

OAI321xp33_ASAP7_75t_L g1697 ( 
.A1(n_1506),
.A2(n_930),
.A3(n_927),
.B1(n_934),
.B2(n_933),
.C(n_920),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1489),
.A2(n_944),
.B(n_937),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1491),
.A2(n_948),
.B(n_945),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1486),
.B(n_941),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1488),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1538),
.A2(n_942),
.B1(n_949),
.B2(n_946),
.Y(n_1702)
);

BUFx2_ASAP7_75t_L g1703 ( 
.A(n_1581),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1492),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1556),
.B(n_1000),
.Y(n_1705)
);

NAND2x1p5_ASAP7_75t_L g1706 ( 
.A(n_1605),
.B(n_1159),
.Y(n_1706)
);

CKINVDCx20_ASAP7_75t_R g1707 ( 
.A(n_1511),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1538),
.A2(n_943),
.B1(n_965),
.B2(n_929),
.Y(n_1708)
);

AOI21xp33_ASAP7_75t_L g1709 ( 
.A1(n_1564),
.A2(n_1135),
.B(n_954),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1566),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1483),
.B(n_969),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1535),
.B(n_1000),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1569),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1546),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1546),
.B(n_973),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1518),
.B(n_969),
.Y(n_1716)
);

NOR2x1p5_ASAP7_75t_L g1717 ( 
.A(n_1529),
.B(n_986),
.Y(n_1717)
);

AOI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1580),
.A2(n_975),
.B(n_974),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1499),
.B(n_951),
.Y(n_1719)
);

BUFx6f_ASAP7_75t_L g1720 ( 
.A(n_1575),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1509),
.A2(n_1012),
.B1(n_1028),
.B2(n_986),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1546),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1473),
.A2(n_979),
.B(n_981),
.C(n_977),
.Y(n_1723)
);

A2O1A1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1583),
.A2(n_988),
.B(n_993),
.C(n_987),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1599),
.B(n_1012),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1646),
.B(n_957),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1497),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1623),
.A2(n_999),
.B(n_998),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1583),
.A2(n_1031),
.B1(n_1044),
.B2(n_1028),
.Y(n_1729)
);

AO21x1_ASAP7_75t_L g1730 ( 
.A1(n_1603),
.A2(n_1004),
.B(n_1001),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1512),
.B(n_958),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1518),
.B(n_1031),
.Y(n_1732)
);

O2A1O1Ixp33_ASAP7_75t_SL g1733 ( 
.A1(n_1479),
.A2(n_1181),
.B(n_1180),
.C(n_1010),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_L g1734 ( 
.A1(n_1589),
.A2(n_960),
.B(n_959),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1593),
.A2(n_1011),
.B(n_1014),
.C(n_1009),
.Y(n_1735)
);

A2O1A1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1539),
.A2(n_1019),
.B(n_1021),
.C(n_1016),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1497),
.A2(n_968),
.B1(n_971),
.B2(n_962),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1521),
.B(n_1023),
.Y(n_1738)
);

BUFx12f_ASAP7_75t_L g1739 ( 
.A(n_1596),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1515),
.B(n_984),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1575),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1527),
.B(n_1026),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1542),
.A2(n_1035),
.B(n_1036),
.C(n_1033),
.Y(n_1743)
);

A2O1A1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1543),
.A2(n_1041),
.B(n_1042),
.C(n_1039),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1575),
.Y(n_1745)
);

AO32x2_ASAP7_75t_L g1746 ( 
.A1(n_1478),
.A2(n_1131),
.A3(n_1075),
.B1(n_1116),
.B2(n_1111),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1503),
.B(n_985),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1519),
.B(n_989),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1493),
.B(n_992),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1561),
.A2(n_1047),
.B(n_1043),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1688),
.B(n_995),
.C(n_994),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1587),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1522),
.B(n_1003),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1602),
.B(n_1044),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1627),
.A2(n_1051),
.B(n_1048),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1523),
.B(n_1525),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1590),
.Y(n_1757)
);

AO21x1_ASAP7_75t_L g1758 ( 
.A1(n_1565),
.A2(n_1060),
.B(n_1054),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1584),
.B(n_1061),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1591),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1490),
.A2(n_1049),
.B1(n_1069),
.B2(n_1045),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1630),
.A2(n_1064),
.B(n_1063),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1636),
.A2(n_1074),
.B(n_1068),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1638),
.A2(n_1078),
.B(n_1076),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1478),
.A2(n_1080),
.B(n_1079),
.Y(n_1765)
);

O2A1O1Ixp33_ASAP7_75t_L g1766 ( 
.A1(n_1570),
.A2(n_1086),
.B(n_1089),
.C(n_1083),
.Y(n_1766)
);

AO21x1_ASAP7_75t_L g1767 ( 
.A1(n_1567),
.A2(n_1091),
.B(n_1090),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1536),
.B(n_1017),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1596),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1590),
.Y(n_1770)
);

OR2x6_ASAP7_75t_L g1771 ( 
.A(n_1632),
.B(n_1116),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1585),
.B(n_1045),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1477),
.A2(n_1096),
.B(n_1093),
.Y(n_1773)
);

NOR3xp33_ASAP7_75t_L g1774 ( 
.A(n_1494),
.B(n_1179),
.C(n_1025),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1553),
.B(n_1018),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1466),
.B(n_1027),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1467),
.B(n_1030),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1469),
.B(n_1034),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1495),
.B(n_1040),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1507),
.B(n_1049),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1477),
.A2(n_1100),
.B(n_1097),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1498),
.B(n_1050),
.Y(n_1782)
);

AND2x2_ASAP7_75t_SL g1783 ( 
.A(n_1507),
.B(n_1069),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1537),
.B(n_1070),
.Y(n_1784)
);

INVx4_ASAP7_75t_L g1785 ( 
.A(n_1526),
.Y(n_1785)
);

O2A1O1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1588),
.A2(n_1106),
.B(n_1108),
.C(n_1104),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1500),
.B(n_1052),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1552),
.B(n_1053),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1482),
.A2(n_1115),
.B(n_1112),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1550),
.A2(n_1124),
.B(n_1122),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1551),
.A2(n_1554),
.B(n_1568),
.Y(n_1791)
);

O2A1O1Ixp33_ASAP7_75t_L g1792 ( 
.A1(n_1579),
.A2(n_1129),
.B(n_1132),
.C(n_1127),
.Y(n_1792)
);

AO21x1_ASAP7_75t_L g1793 ( 
.A1(n_1574),
.A2(n_1140),
.B(n_1138),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1530),
.B(n_1056),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1592),
.A2(n_1604),
.B(n_1594),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1532),
.B(n_1057),
.Y(n_1796)
);

NOR2x1_ASAP7_75t_L g1797 ( 
.A(n_1596),
.B(n_1070),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1664),
.A2(n_1150),
.B(n_1149),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1631),
.A2(n_1152),
.B(n_1151),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1534),
.B(n_1059),
.Y(n_1800)
);

O2A1O1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1617),
.A2(n_1155),
.B(n_1156),
.C(n_1154),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1571),
.A2(n_1085),
.B1(n_1113),
.B2(n_1071),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1634),
.A2(n_1158),
.B(n_1157),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1548),
.B(n_1071),
.Y(n_1804)
);

NOR2xp67_ASAP7_75t_L g1805 ( 
.A(n_1616),
.B(n_34),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1642),
.A2(n_1163),
.B(n_1161),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1598),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_L g1808 ( 
.A(n_1586),
.B(n_1085),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1549),
.B(n_1113),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1472),
.B(n_1067),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1571),
.A2(n_1165),
.B1(n_1169),
.B2(n_1164),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1598),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1597),
.B(n_1547),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1644),
.A2(n_1170),
.B(n_1166),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1555),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1513),
.Y(n_1816)
);

OA22x2_ASAP7_75t_L g1817 ( 
.A1(n_1496),
.A2(n_1165),
.B1(n_1169),
.B2(n_1164),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1609),
.A2(n_1177),
.B(n_1176),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1508),
.Y(n_1819)
);

OAI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1496),
.A2(n_1168),
.B(n_1160),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1622),
.B(n_1175),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1475),
.B(n_1480),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1626),
.A2(n_1171),
.B(n_1146),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1468),
.B(n_1175),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1562),
.A2(n_1077),
.B1(n_1082),
.B2(n_1072),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1633),
.A2(n_1171),
.B(n_1087),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1618),
.A2(n_1088),
.B(n_1084),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1625),
.A2(n_1094),
.B(n_1095),
.C(n_1092),
.Y(n_1828)
);

NAND2x1p5_ASAP7_75t_L g1829 ( 
.A(n_1610),
.B(n_1178),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1516),
.B(n_1099),
.Y(n_1830)
);

INVx6_ASAP7_75t_L g1831 ( 
.A(n_1632),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1559),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1607),
.B(n_1102),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1560),
.B(n_1105),
.Y(n_1834)
);

O2A1O1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1649),
.A2(n_1131),
.B(n_1110),
.C(n_1114),
.Y(n_1835)
);

NOR2x1_ASAP7_75t_L g1836 ( 
.A(n_1586),
.B(n_1109),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1635),
.B(n_1117),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1639),
.A2(n_1120),
.B(n_1119),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1641),
.A2(n_1125),
.B(n_1123),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1648),
.A2(n_1133),
.B(n_1126),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1582),
.B(n_1147),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1619),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1502),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1501),
.Y(n_1844)
);

BUFx12f_ASAP7_75t_L g1845 ( 
.A(n_1643),
.Y(n_1845)
);

BUFx8_ASAP7_75t_SL g1846 ( 
.A(n_1586),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1619),
.Y(n_1847)
);

AND2x6_ASAP7_75t_SL g1848 ( 
.A(n_1517),
.B(n_1183),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1562),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1544),
.B(n_36),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1558),
.A2(n_40),
.B(n_37),
.C(n_39),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1668),
.A2(n_1474),
.B(n_1675),
.Y(n_1852)
);

NOR2x1_ASAP7_75t_L g1853 ( 
.A(n_1616),
.B(n_1517),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1640),
.B(n_39),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1680),
.A2(n_40),
.B(n_41),
.Y(n_1855)
);

OAI321xp33_ASAP7_75t_L g1856 ( 
.A1(n_1615),
.A2(n_1629),
.A3(n_1640),
.B1(n_1671),
.B2(n_1651),
.C(n_1517),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1606),
.Y(n_1857)
);

NOR2xp67_ASAP7_75t_L g1858 ( 
.A(n_1540),
.B(n_41),
.Y(n_1858)
);

AO32x1_ASAP7_75t_L g1859 ( 
.A1(n_1465),
.A2(n_44),
.A3(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1510),
.B(n_42),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1572),
.B(n_46),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1681),
.A2(n_46),
.B(n_47),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1573),
.B(n_1608),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_SL g1864 ( 
.A(n_1645),
.B(n_47),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1682),
.A2(n_48),
.B(n_49),
.Y(n_1865)
);

A2O1A1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1659),
.A2(n_51),
.B(n_48),
.C(n_49),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1504),
.Y(n_1867)
);

NOR2x1_ASAP7_75t_L g1868 ( 
.A(n_1610),
.B(n_52),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1481),
.B(n_53),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1685),
.A2(n_53),
.B(n_54),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1520),
.Y(n_1871)
);

OR2x6_ASAP7_75t_L g1872 ( 
.A(n_1621),
.B(n_55),
.Y(n_1872)
);

NOR2xp67_ASAP7_75t_SL g1873 ( 
.A(n_1619),
.B(n_56),
.Y(n_1873)
);

O2A1O1Ixp33_ASAP7_75t_L g1874 ( 
.A1(n_1612),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1874)
);

OAI321xp33_ASAP7_75t_L g1875 ( 
.A1(n_1651),
.A2(n_1660),
.A3(n_1624),
.B1(n_1620),
.B2(n_1637),
.C(n_1628),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1600),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1876)
);

NAND3xp33_ASAP7_75t_L g1877 ( 
.A(n_1600),
.B(n_61),
.C(n_62),
.Y(n_1877)
);

INVx11_ASAP7_75t_L g1878 ( 
.A(n_1524),
.Y(n_1878)
);

O2A1O1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1613),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_1879)
);

BUFx8_ASAP7_75t_L g1880 ( 
.A(n_1531),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1528),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1531),
.B(n_66),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1533),
.B(n_752),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1650),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1470),
.A2(n_70),
.B(n_71),
.Y(n_1885)
);

BUFx6f_ASAP7_75t_L g1886 ( 
.A(n_1657),
.Y(n_1886)
);

AND2x2_ASAP7_75t_SL g1887 ( 
.A(n_1476),
.B(n_71),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1541),
.A2(n_1557),
.B(n_1545),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1656),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1667),
.A2(n_73),
.B(n_74),
.Y(n_1890)
);

AOI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1669),
.A2(n_73),
.B(n_75),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1595),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1660),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1601),
.A2(n_78),
.B(n_79),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1652),
.B(n_80),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1611),
.B(n_81),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1614),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1670),
.A2(n_83),
.B(n_84),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1672),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1665),
.B(n_85),
.Y(n_1900)
);

NOR2xp67_ASAP7_75t_L g1901 ( 
.A(n_1676),
.B(n_86),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1683),
.B(n_87),
.Y(n_1902)
);

OAI22xp5_ASAP7_75t_L g1903 ( 
.A1(n_1647),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1663),
.B(n_88),
.Y(n_1904)
);

AOI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1686),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1657),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1653),
.B(n_1655),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1485),
.A2(n_97),
.B(n_98),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1654),
.B(n_1666),
.Y(n_1909)
);

CKINVDCx6p67_ASAP7_75t_R g1910 ( 
.A(n_1657),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1661),
.Y(n_1911)
);

INVx5_ASAP7_75t_L g1912 ( 
.A(n_1661),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1661),
.B(n_99),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1674),
.Y(n_1914)
);

OAI21xp33_ASAP7_75t_L g1915 ( 
.A1(n_1678),
.A2(n_100),
.B(n_101),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1684),
.B(n_102),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1687),
.A2(n_103),
.B(n_106),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1674),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1674),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1658),
.B(n_103),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1673),
.Y(n_1921)
);

OAI21xp33_ASAP7_75t_L g1922 ( 
.A1(n_1679),
.A2(n_106),
.B(n_107),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1662),
.B(n_109),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1677),
.B(n_110),
.Y(n_1924)
);

AO32x2_ASAP7_75t_L g1925 ( 
.A1(n_1677),
.A2(n_112),
.A3(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_SL g1926 ( 
.A1(n_1518),
.A2(n_117),
.B1(n_114),
.B2(n_116),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1578),
.A2(n_118),
.B(n_119),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1487),
.B(n_119),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1505),
.B(n_120),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1575),
.Y(n_1930)
);

A2O1A1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1514),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_1931)
);

AOI21xp33_ASAP7_75t_L g1932 ( 
.A1(n_1564),
.A2(n_123),
.B(n_125),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1505),
.B(n_125),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1505),
.B(n_126),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1578),
.A2(n_126),
.B(n_127),
.Y(n_1935)
);

OAI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1538),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1483),
.B(n_767),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1538),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_1938)
);

A2O1A1Ixp33_ASAP7_75t_L g1939 ( 
.A1(n_1514),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1578),
.A2(n_131),
.B(n_132),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1578),
.A2(n_134),
.B(n_135),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1471),
.Y(n_1942)
);

OAI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1538),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1556),
.B(n_136),
.Y(n_1944)
);

HB1xp67_ASAP7_75t_L g1945 ( 
.A(n_1577),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1605),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1576),
.Y(n_1947)
);

AND2x6_ASAP7_75t_L g1948 ( 
.A(n_1886),
.B(n_138),
.Y(n_1948)
);

BUFx6f_ASAP7_75t_L g1949 ( 
.A(n_1720),
.Y(n_1949)
);

OAI21x1_ASAP7_75t_L g1950 ( 
.A1(n_1689),
.A2(n_138),
.B(n_139),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1757),
.B(n_139),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1791),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_1952)
);

INVxp67_ASAP7_75t_L g1953 ( 
.A(n_1946),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1701),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1770),
.B(n_1807),
.Y(n_1955)
);

AO31x2_ASAP7_75t_L g1956 ( 
.A1(n_1730),
.A2(n_1767),
.A3(n_1793),
.B(n_1758),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1795),
.A2(n_140),
.B(n_141),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1716),
.B(n_142),
.Y(n_1958)
);

NOR2xp67_ASAP7_75t_L g1959 ( 
.A(n_1739),
.B(n_143),
.Y(n_1959)
);

OAI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1765),
.A2(n_143),
.B(n_144),
.Y(n_1960)
);

NOR3xp33_ASAP7_75t_L g1961 ( 
.A(n_1856),
.B(n_144),
.C(n_145),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1802),
.B(n_1811),
.Y(n_1962)
);

INVxp67_ASAP7_75t_L g1963 ( 
.A(n_1706),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1722),
.B(n_1704),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1816),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1696),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1812),
.B(n_147),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1756),
.B(n_147),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1815),
.B(n_148),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1707),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1720),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1947),
.B(n_149),
.Y(n_1972)
);

OAI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1698),
.A2(n_150),
.B(n_151),
.Y(n_1973)
);

A2O1A1Ixp33_ASAP7_75t_L g1974 ( 
.A1(n_1813),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_1974)
);

AO21x1_ASAP7_75t_L g1975 ( 
.A1(n_1894),
.A2(n_152),
.B(n_153),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1710),
.Y(n_1976)
);

AOI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1822),
.A2(n_154),
.B(n_155),
.Y(n_1977)
);

INVx1_ASAP7_75t_SL g1978 ( 
.A(n_1910),
.Y(n_1978)
);

OAI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1699),
.A2(n_154),
.B(n_156),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1833),
.B(n_158),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1893),
.A2(n_162),
.B1(n_159),
.B2(n_161),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1852),
.A2(n_161),
.B(n_162),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1784),
.B(n_748),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1761),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1899),
.B(n_166),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1832),
.B(n_167),
.Y(n_1986)
);

AO31x2_ASAP7_75t_L g1987 ( 
.A1(n_1931),
.A2(n_171),
.A3(n_168),
.B(n_170),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1732),
.B(n_168),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1912),
.B(n_172),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1752),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1912),
.B(n_175),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1713),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_L g1993 ( 
.A(n_1824),
.B(n_176),
.C(n_179),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1692),
.B(n_181),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1912),
.B(n_182),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1886),
.Y(n_1996)
);

AO32x2_ASAP7_75t_L g1997 ( 
.A1(n_1936),
.A2(n_185),
.A3(n_183),
.B1(n_184),
.B2(n_187),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1783),
.B(n_188),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1760),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1773),
.B(n_1781),
.Y(n_2000)
);

AO31x2_ASAP7_75t_L g2001 ( 
.A1(n_1939),
.A2(n_190),
.A3(n_188),
.B(n_189),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1843),
.Y(n_2002)
);

O2A1O1Ixp5_ASAP7_75t_L g2003 ( 
.A1(n_1850),
.A2(n_193),
.B(n_191),
.C(n_192),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1780),
.B(n_1937),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1790),
.B(n_193),
.Y(n_2005)
);

AO31x2_ASAP7_75t_L g2006 ( 
.A1(n_1866),
.A2(n_196),
.A3(n_194),
.B(n_195),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1789),
.B(n_198),
.Y(n_2007)
);

NAND2xp33_ASAP7_75t_SL g2008 ( 
.A(n_1918),
.B(n_749),
.Y(n_2008)
);

AO31x2_ASAP7_75t_L g2009 ( 
.A1(n_1943),
.A2(n_200),
.A3(n_198),
.B(n_199),
.Y(n_2009)
);

NOR2x1_ASAP7_75t_L g2010 ( 
.A(n_1836),
.B(n_1872),
.Y(n_2010)
);

AO32x2_ASAP7_75t_L g2011 ( 
.A1(n_1903),
.A2(n_203),
.A3(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_2011)
);

O2A1O1Ixp5_ASAP7_75t_L g2012 ( 
.A1(n_1864),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_2012)
);

AOI21xp5_ASAP7_75t_L g2013 ( 
.A1(n_1888),
.A2(n_205),
.B(n_206),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1831),
.Y(n_2014)
);

O2A1O1Ixp5_ASAP7_75t_L g2015 ( 
.A1(n_1902),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_2015)
);

NOR2x1_ASAP7_75t_L g2016 ( 
.A(n_1872),
.B(n_209),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1844),
.Y(n_2017)
);

BUFx3_ASAP7_75t_L g2018 ( 
.A(n_1831),
.Y(n_2018)
);

OAI21x1_ASAP7_75t_L g2019 ( 
.A1(n_1718),
.A2(n_210),
.B(n_211),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1929),
.A2(n_212),
.B(n_213),
.Y(n_2020)
);

OAI21x1_ASAP7_75t_L g2021 ( 
.A1(n_1923),
.A2(n_212),
.B(n_214),
.Y(n_2021)
);

INVx5_ASAP7_75t_L g2022 ( 
.A(n_1918),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1906),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1933),
.B(n_215),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_1934),
.A2(n_1745),
.B(n_1741),
.Y(n_2025)
);

OAI21x1_ASAP7_75t_L g2026 ( 
.A1(n_1924),
.A2(n_216),
.B(n_217),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_1705),
.B(n_217),
.C(n_219),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1906),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1711),
.B(n_220),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1821),
.B(n_1712),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1818),
.B(n_221),
.Y(n_2031)
);

OAI21xp33_ASAP7_75t_L g2032 ( 
.A1(n_1804),
.A2(n_224),
.B(n_225),
.Y(n_2032)
);

AOI221xp5_ASAP7_75t_SL g2033 ( 
.A1(n_1736),
.A2(n_231),
.B1(n_228),
.B2(n_229),
.C(n_232),
.Y(n_2033)
);

A2O1A1Ixp33_ASAP7_75t_L g2034 ( 
.A1(n_1900),
.A2(n_233),
.B(n_228),
.C(n_232),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1714),
.B(n_1889),
.Y(n_2035)
);

NAND3xp33_ASAP7_75t_SL g2036 ( 
.A(n_1926),
.B(n_233),
.C(n_234),
.Y(n_2036)
);

OAI21x1_ASAP7_75t_L g2037 ( 
.A1(n_1920),
.A2(n_234),
.B(n_235),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1693),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1846),
.Y(n_2039)
);

A2O1A1Ixp33_ASAP7_75t_L g2040 ( 
.A1(n_1904),
.A2(n_1895),
.B(n_1750),
.C(n_1798),
.Y(n_2040)
);

AOI21x1_ASAP7_75t_L g2041 ( 
.A1(n_1901),
.A2(n_237),
.B(n_239),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1755),
.B(n_240),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1853),
.B(n_241),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1938),
.A2(n_246),
.B1(n_243),
.B2(n_245),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1762),
.B(n_245),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1708),
.B(n_1729),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1867),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1763),
.B(n_248),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1871),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1764),
.B(n_249),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1702),
.B(n_250),
.Y(n_2051)
);

OAI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1724),
.A2(n_1828),
.B(n_1823),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1774),
.B(n_251),
.Y(n_2053)
);

AO21x1_ASAP7_75t_L g2054 ( 
.A1(n_1927),
.A2(n_251),
.B(n_252),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1942),
.B(n_252),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1715),
.B(n_255),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_1703),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1809),
.B(n_1721),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1860),
.Y(n_2059)
);

OAI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1728),
.A2(n_1940),
.B(n_1935),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1892),
.Y(n_2061)
);

INVx8_ASAP7_75t_L g2062 ( 
.A(n_1771),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1759),
.Y(n_2063)
);

AO31x2_ASAP7_75t_L g2064 ( 
.A1(n_1743),
.A2(n_260),
.A3(n_257),
.B(n_259),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1825),
.B(n_261),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_1829),
.B(n_262),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1723),
.B(n_265),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1715),
.B(n_267),
.Y(n_2068)
);

AO31x2_ASAP7_75t_L g2069 ( 
.A1(n_1744),
.A2(n_274),
.A3(n_268),
.B(n_272),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1878),
.Y(n_2070)
);

A2O1A1Ixp33_ASAP7_75t_L g2071 ( 
.A1(n_1735),
.A2(n_279),
.B(n_275),
.C(n_276),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_SL g2072 ( 
.A1(n_1930),
.A2(n_275),
.B(n_276),
.Y(n_2072)
);

BUFx10_ASAP7_75t_L g2073 ( 
.A(n_1771),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1691),
.B(n_279),
.Y(n_2074)
);

OAI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_1941),
.A2(n_282),
.B(n_283),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1737),
.B(n_282),
.Y(n_2076)
);

BUFx2_ASAP7_75t_L g2077 ( 
.A(n_1880),
.Y(n_2077)
);

AO21x2_ASAP7_75t_L g2078 ( 
.A1(n_1869),
.A2(n_284),
.B(n_285),
.Y(n_2078)
);

AOI221xp5_ASAP7_75t_SL g2079 ( 
.A1(n_1766),
.A2(n_288),
.B1(n_286),
.B2(n_287),
.C(n_289),
.Y(n_2079)
);

NAND3xp33_ASAP7_75t_L g2080 ( 
.A(n_1944),
.B(n_289),
.C(n_290),
.Y(n_2080)
);

AOI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_1930),
.A2(n_1837),
.B(n_1788),
.Y(n_2081)
);

AO31x2_ASAP7_75t_L g2082 ( 
.A1(n_1885),
.A2(n_292),
.A3(n_290),
.B(n_291),
.Y(n_2082)
);

AO31x2_ASAP7_75t_L g2083 ( 
.A1(n_1855),
.A2(n_295),
.A3(n_292),
.B(n_294),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_1909),
.A2(n_297),
.B(n_299),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1759),
.Y(n_2085)
);

AO21x1_ASAP7_75t_L g2086 ( 
.A1(n_1851),
.A2(n_300),
.B(n_301),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1883),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_1725),
.B(n_304),
.Y(n_2088)
);

AO21x1_ASAP7_75t_L g2089 ( 
.A1(n_1916),
.A2(n_306),
.B(n_307),
.Y(n_2089)
);

AOI221x1_ASAP7_75t_L g2090 ( 
.A1(n_1915),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.C(n_310),
.Y(n_2090)
);

BUFx3_ASAP7_75t_L g2091 ( 
.A(n_1880),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1826),
.B(n_311),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1842),
.Y(n_2093)
);

AOI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_1779),
.A2(n_311),
.B(n_313),
.Y(n_2094)
);

NOR2xp67_ASAP7_75t_L g2095 ( 
.A(n_1857),
.B(n_313),
.Y(n_2095)
);

A2O1A1Ixp33_ASAP7_75t_L g2096 ( 
.A1(n_1862),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_2096)
);

NOR2x1_ASAP7_75t_SL g2097 ( 
.A(n_1842),
.B(n_315),
.Y(n_2097)
);

INVx3_ASAP7_75t_L g2098 ( 
.A(n_1785),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_1887),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1817),
.B(n_319),
.Y(n_2100)
);

BUFx2_ASAP7_75t_L g2101 ( 
.A(n_1945),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1884),
.B(n_320),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1847),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_1738),
.B(n_320),
.Y(n_2104)
);

A2O1A1Ixp33_ASAP7_75t_L g2105 ( 
.A1(n_1865),
.A2(n_323),
.B(n_321),
.C(n_322),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_1754),
.B(n_321),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1738),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1921),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1799),
.B(n_325),
.Y(n_2109)
);

OAI21x1_ASAP7_75t_L g2110 ( 
.A1(n_1896),
.A2(n_325),
.B(n_328),
.Y(n_2110)
);

BUFx6f_ASAP7_75t_L g2111 ( 
.A(n_1847),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1803),
.B(n_328),
.Y(n_2112)
);

AOI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_1782),
.A2(n_329),
.B(n_330),
.Y(n_2113)
);

NOR2xp67_ASAP7_75t_L g2114 ( 
.A(n_1845),
.B(n_1727),
.Y(n_2114)
);

A2O1A1Ixp33_ASAP7_75t_L g2115 ( 
.A1(n_1870),
.A2(n_332),
.B(n_329),
.C(n_330),
.Y(n_2115)
);

NOR2x1_ASAP7_75t_SL g2116 ( 
.A(n_1847),
.B(n_1690),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1911),
.Y(n_2117)
);

O2A1O1Ixp5_ASAP7_75t_L g2118 ( 
.A1(n_1873),
.A2(n_1928),
.B(n_1854),
.C(n_1913),
.Y(n_2118)
);

AND2x6_ASAP7_75t_L g2119 ( 
.A(n_1914),
.B(n_333),
.Y(n_2119)
);

A2O1A1Ixp33_ASAP7_75t_L g2120 ( 
.A1(n_1890),
.A2(n_336),
.B(n_334),
.C(n_335),
.Y(n_2120)
);

AOI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_1787),
.A2(n_334),
.B(n_335),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1806),
.B(n_336),
.Y(n_2122)
);

AOI211x1_ASAP7_75t_L g2123 ( 
.A1(n_1932),
.A2(n_339),
.B(n_337),
.C(n_338),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1861),
.B(n_338),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1814),
.B(n_339),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1742),
.B(n_341),
.Y(n_2126)
);

INVx1_ASAP7_75t_SL g2127 ( 
.A(n_1695),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1694),
.A2(n_1719),
.B(n_1700),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1742),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1775),
.B(n_342),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1748),
.Y(n_2131)
);

NOR3xp33_ASAP7_75t_L g2132 ( 
.A(n_1734),
.B(n_343),
.C(n_344),
.Y(n_2132)
);

CKINVDCx11_ASAP7_75t_R g2133 ( 
.A(n_1848),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1907),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1794),
.Y(n_2135)
);

OAI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_1697),
.A2(n_346),
.B(n_347),
.Y(n_2136)
);

OR2x6_ASAP7_75t_L g2137 ( 
.A(n_1769),
.B(n_347),
.Y(n_2137)
);

AO31x2_ASAP7_75t_L g2138 ( 
.A1(n_1891),
.A2(n_351),
.A3(n_348),
.B(n_349),
.Y(n_2138)
);

INVx1_ASAP7_75t_SL g2139 ( 
.A(n_1695),
.Y(n_2139)
);

OAI22xp5_ASAP7_75t_L g2140 ( 
.A1(n_1849),
.A2(n_351),
.B1(n_348),
.B2(n_349),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1772),
.B(n_352),
.Y(n_2141)
);

OA21x2_ASAP7_75t_L g2142 ( 
.A1(n_1922),
.A2(n_352),
.B(n_354),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_SL g2143 ( 
.A1(n_1874),
.A2(n_354),
.B(n_355),
.Y(n_2143)
);

AO22x2_ASAP7_75t_L g2144 ( 
.A1(n_1877),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1796),
.Y(n_2145)
);

AO31x2_ASAP7_75t_L g2146 ( 
.A1(n_1898),
.A2(n_365),
.A3(n_363),
.B(n_364),
.Y(n_2146)
);

OAI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_1875),
.A2(n_365),
.B(n_366),
.Y(n_2147)
);

BUFx6f_ASAP7_75t_L g2148 ( 
.A(n_1919),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_1776),
.A2(n_366),
.B(n_367),
.Y(n_2149)
);

AOI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_1777),
.A2(n_369),
.B(n_371),
.Y(n_2150)
);

BUFx3_ASAP7_75t_L g2151 ( 
.A(n_1785),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_1907),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_1726),
.B(n_373),
.Y(n_2153)
);

OA22x2_ASAP7_75t_L g2154 ( 
.A1(n_1876),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1747),
.B(n_374),
.Y(n_2155)
);

OAI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_1905),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_2156)
);

OAI21xp33_ASAP7_75t_L g2157 ( 
.A1(n_1749),
.A2(n_376),
.B(n_379),
.Y(n_2157)
);

OR2x2_ASAP7_75t_L g2158 ( 
.A(n_1717),
.B(n_379),
.Y(n_2158)
);

AOI21xp33_ASAP7_75t_L g2159 ( 
.A1(n_1879),
.A2(n_380),
.B(n_381),
.Y(n_2159)
);

OAI21xp5_ASAP7_75t_L g2160 ( 
.A1(n_1792),
.A2(n_380),
.B(n_383),
.Y(n_2160)
);

AOI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_1778),
.A2(n_383),
.B(n_384),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1753),
.B(n_1768),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_1820),
.A2(n_388),
.B1(n_385),
.B2(n_386),
.Y(n_2163)
);

OAI21xp33_ASAP7_75t_L g2164 ( 
.A1(n_1731),
.A2(n_385),
.B(n_386),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1801),
.B(n_388),
.Y(n_2165)
);

NOR2x1_ASAP7_75t_SL g2166 ( 
.A(n_1690),
.B(n_389),
.Y(n_2166)
);

AO31x2_ASAP7_75t_L g2167 ( 
.A1(n_1908),
.A2(n_394),
.A3(n_391),
.B(n_392),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1740),
.B(n_396),
.Y(n_2168)
);

OAI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_1881),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_1827),
.B(n_397),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1830),
.B(n_400),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_1838),
.B(n_1839),
.Y(n_2172)
);

OAI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_1786),
.A2(n_400),
.B(n_402),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1897),
.Y(n_2174)
);

NAND2x1p5_ASAP7_75t_L g2175 ( 
.A(n_1868),
.B(n_402),
.Y(n_2175)
);

A2O1A1Ixp33_ASAP7_75t_L g2176 ( 
.A1(n_1805),
.A2(n_407),
.B(n_403),
.C(n_405),
.Y(n_2176)
);

OAI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_1840),
.A2(n_408),
.B(n_409),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_1709),
.B(n_410),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_1805),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1810),
.B(n_412),
.Y(n_2180)
);

OAI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_1882),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1800),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1841),
.B(n_1835),
.Y(n_2183)
);

OAI211xp5_ASAP7_75t_L g2184 ( 
.A1(n_1797),
.A2(n_418),
.B(n_416),
.C(n_417),
.Y(n_2184)
);

AOI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_1834),
.A2(n_417),
.B(n_418),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_1863),
.Y(n_2186)
);

INVx2_ASAP7_75t_SL g2187 ( 
.A(n_1819),
.Y(n_2187)
);

CKINVDCx12_ASAP7_75t_R g2188 ( 
.A(n_1808),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1746),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1751),
.B(n_420),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_1858),
.B(n_421),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_1925),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_1746),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_2193)
);

AOI31xp67_ASAP7_75t_L g2194 ( 
.A1(n_1746),
.A2(n_1859),
.A3(n_1925),
.B(n_1733),
.Y(n_2194)
);

A2O1A1Ixp33_ASAP7_75t_L g2195 ( 
.A1(n_1859),
.A2(n_429),
.B(n_426),
.C(n_427),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1757),
.B(n_429),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1701),
.Y(n_2197)
);

AOI221x1_ASAP7_75t_L g2198 ( 
.A1(n_1915),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.C(n_433),
.Y(n_2198)
);

OAI21xp33_ASAP7_75t_L g2199 ( 
.A1(n_1833),
.A2(n_430),
.B(n_432),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1757),
.B(n_434),
.Y(n_2200)
);

A2O1A1Ixp33_ASAP7_75t_L g2201 ( 
.A1(n_1791),
.A2(n_437),
.B(n_435),
.C(n_436),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_1720),
.Y(n_2202)
);

AOI21xp5_ASAP7_75t_L g2203 ( 
.A1(n_1795),
.A2(n_435),
.B(n_439),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1757),
.B(n_440),
.Y(n_2204)
);

INVx5_ASAP7_75t_L g2205 ( 
.A(n_1886),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1701),
.Y(n_2206)
);

OAI21x1_ASAP7_75t_L g2207 ( 
.A1(n_1689),
.A2(n_440),
.B(n_441),
.Y(n_2207)
);

OAI21x1_ASAP7_75t_L g2208 ( 
.A1(n_1689),
.A2(n_443),
.B(n_444),
.Y(n_2208)
);

BUFx12f_ASAP7_75t_L g2209 ( 
.A(n_1739),
.Y(n_2209)
);

OAI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1757),
.A2(n_446),
.B1(n_443),
.B2(n_445),
.Y(n_2210)
);

INVx4_ASAP7_75t_L g2211 ( 
.A(n_1912),
.Y(n_2211)
);

INVx2_ASAP7_75t_SL g2212 ( 
.A(n_1831),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_1716),
.B(n_445),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1757),
.B(n_447),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1757),
.B(n_448),
.Y(n_2215)
);

BUFx3_ASAP7_75t_L g2216 ( 
.A(n_1831),
.Y(n_2216)
);

AO21x2_ASAP7_75t_L g2217 ( 
.A1(n_1765),
.A2(n_449),
.B(n_452),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1716),
.B(n_452),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1757),
.B(n_454),
.Y(n_2219)
);

OAI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_1757),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1757),
.B(n_455),
.Y(n_2221)
);

NAND2x1p5_ASAP7_75t_L g2222 ( 
.A(n_1912),
.B(n_457),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_SL g2223 ( 
.A(n_1912),
.B(n_457),
.Y(n_2223)
);

NAND2xp33_ASAP7_75t_L g2224 ( 
.A(n_1720),
.B(n_458),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1757),
.B(n_458),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_1946),
.Y(n_2226)
);

AO31x2_ASAP7_75t_L g2227 ( 
.A1(n_1730),
.A2(n_461),
.A3(n_459),
.B(n_460),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_1912),
.B(n_462),
.Y(n_2228)
);

OAI21x1_ASAP7_75t_L g2229 ( 
.A1(n_1689),
.A2(n_463),
.B(n_465),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1716),
.B(n_465),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1701),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1757),
.B(n_466),
.Y(n_2232)
);

BUFx8_ASAP7_75t_L g2233 ( 
.A(n_1739),
.Y(n_2233)
);

AOI21xp33_ASAP7_75t_L g2234 ( 
.A1(n_1902),
.A2(n_468),
.B(n_469),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_1757),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1701),
.Y(n_2236)
);

OAI21xp5_ASAP7_75t_L g2237 ( 
.A1(n_1791),
.A2(n_474),
.B(n_475),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_1707),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1757),
.B(n_474),
.Y(n_2239)
);

INVx1_ASAP7_75t_SL g2240 ( 
.A(n_1946),
.Y(n_2240)
);

OAI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_1757),
.A2(n_479),
.B1(n_477),
.B2(n_478),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1696),
.Y(n_2242)
);

A2O1A1Ixp33_ASAP7_75t_L g2243 ( 
.A1(n_1791),
.A2(n_482),
.B(n_480),
.C(n_481),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1716),
.B(n_481),
.Y(n_2244)
);

AOI21xp5_ASAP7_75t_L g2245 ( 
.A1(n_1795),
.A2(n_482),
.B(n_483),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_1757),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.Y(n_2246)
);

AOI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_1795),
.A2(n_484),
.B(n_487),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1757),
.B(n_488),
.Y(n_2248)
);

AND2x4_ASAP7_75t_L g2249 ( 
.A(n_1722),
.B(n_490),
.Y(n_2249)
);

OAI21x1_ASAP7_75t_L g2250 ( 
.A1(n_1689),
.A2(n_492),
.B(n_493),
.Y(n_2250)
);

OAI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_1757),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_2251)
);

AOI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_1795),
.A2(n_494),
.B(n_497),
.Y(n_2252)
);

AO31x2_ASAP7_75t_L g2253 ( 
.A1(n_1730),
.A2(n_500),
.A3(n_497),
.B(n_499),
.Y(n_2253)
);

AOI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_1795),
.A2(n_501),
.B(n_502),
.Y(n_2254)
);

OAI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_1791),
.A2(n_501),
.B(n_502),
.Y(n_2255)
);

AO21x1_ASAP7_75t_L g2256 ( 
.A1(n_1894),
.A2(n_503),
.B(n_504),
.Y(n_2256)
);

A2O1A1Ixp33_ASAP7_75t_L g2257 ( 
.A1(n_1791),
.A2(n_506),
.B(n_503),
.C(n_504),
.Y(n_2257)
);

OA22x2_ASAP7_75t_L g2258 ( 
.A1(n_1716),
.A2(n_510),
.B1(n_507),
.B2(n_509),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1701),
.Y(n_2259)
);

A2O1A1Ixp33_ASAP7_75t_L g2260 ( 
.A1(n_1791),
.A2(n_512),
.B(n_509),
.C(n_511),
.Y(n_2260)
);

INVx1_ASAP7_75t_SL g2261 ( 
.A(n_1946),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_1946),
.B(n_514),
.Y(n_2262)
);

CKINVDCx20_ASAP7_75t_R g2263 ( 
.A(n_1707),
.Y(n_2263)
);

OAI21x1_ASAP7_75t_SL g2264 ( 
.A1(n_1917),
.A2(n_515),
.B(n_516),
.Y(n_2264)
);

OAI21x1_ASAP7_75t_L g2265 ( 
.A1(n_1689),
.A2(n_516),
.B(n_517),
.Y(n_2265)
);

AND2x4_ASAP7_75t_L g2266 ( 
.A(n_1722),
.B(n_517),
.Y(n_2266)
);

A2O1A1Ixp33_ASAP7_75t_L g2267 ( 
.A1(n_1791),
.A2(n_520),
.B(n_518),
.C(n_519),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1757),
.B(n_521),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1946),
.B(n_521),
.Y(n_2269)
);

AOI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_1795),
.A2(n_522),
.B(n_523),
.Y(n_2270)
);

AOI21xp5_ASAP7_75t_L g2271 ( 
.A1(n_1795),
.A2(n_522),
.B(n_524),
.Y(n_2271)
);

AOI21xp5_ASAP7_75t_L g2272 ( 
.A1(n_1795),
.A2(n_525),
.B(n_527),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1757),
.B(n_527),
.Y(n_2273)
);

INVxp67_ASAP7_75t_SL g2274 ( 
.A(n_1729),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_1757),
.B(n_529),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1757),
.B(n_529),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_1757),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.Y(n_2277)
);

BUFx4f_ASAP7_75t_SL g2278 ( 
.A(n_1707),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1757),
.B(n_533),
.Y(n_2279)
);

OAI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_1791),
.A2(n_534),
.B(n_535),
.Y(n_2280)
);

NAND2x1p5_ASAP7_75t_L g2281 ( 
.A(n_1912),
.B(n_534),
.Y(n_2281)
);

BUFx2_ASAP7_75t_SL g2282 ( 
.A(n_1707),
.Y(n_2282)
);

OAI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_1791),
.A2(n_536),
.B(n_538),
.Y(n_2283)
);

O2A1O1Ixp5_ASAP7_75t_L g2284 ( 
.A1(n_1730),
.A2(n_541),
.B(n_539),
.C(n_540),
.Y(n_2284)
);

AO31x2_ASAP7_75t_L g2285 ( 
.A1(n_1730),
.A2(n_542),
.A3(n_539),
.B(n_541),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_1946),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1696),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1696),
.Y(n_2288)
);

AOI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_1795),
.A2(n_542),
.B(n_545),
.Y(n_2289)
);

INVx2_ASAP7_75t_SL g2290 ( 
.A(n_1831),
.Y(n_2290)
);

AOI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_1795),
.A2(n_546),
.B(n_547),
.Y(n_2291)
);

AOI21xp5_ASAP7_75t_L g2292 ( 
.A1(n_1795),
.A2(n_549),
.B(n_550),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1757),
.B(n_549),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1757),
.B(n_551),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1701),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1701),
.Y(n_2296)
);

BUFx3_ASAP7_75t_L g2297 ( 
.A(n_1831),
.Y(n_2297)
);

INVx1_ASAP7_75t_SL g2298 ( 
.A(n_1946),
.Y(n_2298)
);

AOI21xp33_ASAP7_75t_L g2299 ( 
.A1(n_1902),
.A2(n_551),
.B(n_552),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_1757),
.B(n_552),
.Y(n_2300)
);

BUFx12f_ASAP7_75t_L g2301 ( 
.A(n_1739),
.Y(n_2301)
);

INVx2_ASAP7_75t_SL g2302 ( 
.A(n_1831),
.Y(n_2302)
);

OAI21xp5_ASAP7_75t_L g2303 ( 
.A1(n_1791),
.A2(n_553),
.B(n_554),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1701),
.Y(n_2304)
);

OAI21x1_ASAP7_75t_L g2305 ( 
.A1(n_1689),
.A2(n_555),
.B(n_556),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_1757),
.B(n_555),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1757),
.B(n_558),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1757),
.B(n_559),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1757),
.B(n_559),
.Y(n_2309)
);

OAI21xp5_ASAP7_75t_L g2310 ( 
.A1(n_1791),
.A2(n_560),
.B(n_561),
.Y(n_2310)
);

OAI21x1_ASAP7_75t_SL g2311 ( 
.A1(n_1917),
.A2(n_561),
.B(n_562),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1757),
.B(n_562),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_1716),
.B(n_563),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1701),
.Y(n_2314)
);

OA22x2_ASAP7_75t_L g2315 ( 
.A1(n_1716),
.A2(n_566),
.B1(n_567),
.B2(n_568),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1757),
.B(n_567),
.Y(n_2316)
);

INVx3_ASAP7_75t_L g2317 ( 
.A(n_1912),
.Y(n_2317)
);

INVx2_ASAP7_75t_SL g2318 ( 
.A(n_1831),
.Y(n_2318)
);

OAI21x1_ASAP7_75t_L g2319 ( 
.A1(n_1689),
.A2(n_569),
.B(n_570),
.Y(n_2319)
);

NAND2x1p5_ASAP7_75t_L g2320 ( 
.A(n_1912),
.B(n_570),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_1716),
.B(n_571),
.Y(n_2321)
);

OAI21x1_ASAP7_75t_L g2322 ( 
.A1(n_1689),
.A2(n_574),
.B(n_575),
.Y(n_2322)
);

INVx2_ASAP7_75t_SL g2323 ( 
.A(n_1831),
.Y(n_2323)
);

BUFx2_ASAP7_75t_L g2324 ( 
.A(n_1946),
.Y(n_2324)
);

OAI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_1757),
.A2(n_575),
.B1(n_576),
.B2(n_577),
.Y(n_2325)
);

AO31x2_ASAP7_75t_L g2326 ( 
.A1(n_1730),
.A2(n_576),
.A3(n_578),
.B(n_579),
.Y(n_2326)
);

OAI21x1_ASAP7_75t_L g2327 ( 
.A1(n_1689),
.A2(n_579),
.B(n_580),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_1696),
.Y(n_2328)
);

OAI21x1_ASAP7_75t_L g2329 ( 
.A1(n_1689),
.A2(n_581),
.B(n_582),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1696),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_1696),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1701),
.Y(n_2332)
);

AOI21xp5_ASAP7_75t_L g2333 ( 
.A1(n_1795),
.A2(n_582),
.B(n_583),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_1716),
.B(n_584),
.Y(n_2334)
);

AOI21xp5_ASAP7_75t_L g2335 ( 
.A1(n_1795),
.A2(n_585),
.B(n_586),
.Y(n_2335)
);

OAI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_1791),
.A2(n_586),
.B(n_587),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1757),
.B(n_588),
.Y(n_2337)
);

NAND2x1p5_ASAP7_75t_L g2338 ( 
.A(n_1912),
.B(n_589),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_1795),
.A2(n_589),
.B(n_590),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_1955),
.B(n_591),
.Y(n_2340)
);

AOI22x1_ASAP7_75t_L g2341 ( 
.A1(n_2128),
.A2(n_591),
.B1(n_592),
.B2(n_593),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_1949),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_1962),
.B(n_592),
.Y(n_2343)
);

OAI21x1_ASAP7_75t_L g2344 ( 
.A1(n_2025),
.A2(n_593),
.B(n_594),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_1954),
.Y(n_2345)
);

INVxp67_ASAP7_75t_L g2346 ( 
.A(n_2286),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1965),
.B(n_2197),
.Y(n_2347)
);

AO21x2_ASAP7_75t_L g2348 ( 
.A1(n_2189),
.A2(n_594),
.B(n_595),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2206),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_1970),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1966),
.Y(n_2351)
);

AOI21xp5_ASAP7_75t_L g2352 ( 
.A1(n_2040),
.A2(n_596),
.B(n_598),
.Y(n_2352)
);

NAND3xp33_ASAP7_75t_L g2353 ( 
.A(n_2123),
.B(n_2132),
.C(n_2027),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2231),
.Y(n_2354)
);

OAI22xp5_ASAP7_75t_L g2355 ( 
.A1(n_2099),
.A2(n_598),
.B1(n_599),
.B2(n_600),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_2236),
.B(n_599),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2226),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2242),
.Y(n_2358)
);

OAI22xp33_ASAP7_75t_L g2359 ( 
.A1(n_2099),
.A2(n_603),
.B1(n_604),
.B2(n_605),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2324),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2259),
.Y(n_2361)
);

INVx3_ASAP7_75t_L g2362 ( 
.A(n_2211),
.Y(n_2362)
);

OAI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2060),
.A2(n_603),
.B(n_604),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2295),
.Y(n_2364)
);

INVx4_ASAP7_75t_L g2365 ( 
.A(n_2022),
.Y(n_2365)
);

O2A1O1Ixp33_ASAP7_75t_SL g2366 ( 
.A1(n_1973),
.A2(n_605),
.B(n_606),
.C(n_608),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2296),
.B(n_606),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2304),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2314),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2332),
.Y(n_2370)
);

OAI21x1_ASAP7_75t_L g2371 ( 
.A1(n_1950),
.A2(n_609),
.B(n_610),
.Y(n_2371)
);

OAI21x1_ASAP7_75t_L g2372 ( 
.A1(n_2207),
.A2(n_611),
.B(n_612),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2017),
.Y(n_2373)
);

OAI21x1_ASAP7_75t_L g2374 ( 
.A1(n_2208),
.A2(n_613),
.B(n_615),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_1969),
.Y(n_2375)
);

AOI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2030),
.A2(n_616),
.B1(n_617),
.B2(n_618),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2000),
.A2(n_617),
.B(n_618),
.Y(n_2377)
);

OAI21x1_ASAP7_75t_L g2378 ( 
.A1(n_2229),
.A2(n_619),
.B(n_620),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1969),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2162),
.B(n_621),
.Y(n_2380)
);

INVx5_ASAP7_75t_L g2381 ( 
.A(n_1948),
.Y(n_2381)
);

OAI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2000),
.A2(n_2162),
.B(n_2052),
.Y(n_2382)
);

CKINVDCx20_ASAP7_75t_R g2383 ( 
.A(n_2278),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2038),
.Y(n_2384)
);

OR2x2_ASAP7_75t_L g2385 ( 
.A(n_2226),
.B(n_2240),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_L g2386 ( 
.A(n_2274),
.B(n_622),
.Y(n_2386)
);

BUFx6f_ASAP7_75t_L g2387 ( 
.A(n_1949),
.Y(n_2387)
);

AOI22xp33_ASAP7_75t_SL g2388 ( 
.A1(n_2046),
.A2(n_622),
.B1(n_623),
.B2(n_624),
.Y(n_2388)
);

OAI21xp5_ASAP7_75t_L g2389 ( 
.A1(n_2052),
.A2(n_2203),
.B(n_1957),
.Y(n_2389)
);

OAI21x1_ASAP7_75t_SL g2390 ( 
.A1(n_1973),
.A2(n_624),
.B(n_625),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2055),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2081),
.A2(n_625),
.B(n_626),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2287),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2135),
.B(n_626),
.Y(n_2394)
);

INVx4_ASAP7_75t_L g2395 ( 
.A(n_2022),
.Y(n_2395)
);

NAND2x1p5_ASAP7_75t_L g2396 ( 
.A(n_2022),
.B(n_627),
.Y(n_2396)
);

OAI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2245),
.A2(n_628),
.B(n_629),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2288),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2058),
.B(n_630),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2055),
.Y(n_2400)
);

OAI21xp5_ASAP7_75t_L g2401 ( 
.A1(n_2247),
.A2(n_631),
.B(n_632),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1990),
.Y(n_2402)
);

AOI22xp5_ASAP7_75t_L g2403 ( 
.A1(n_2004),
.A2(n_631),
.B1(n_632),
.B2(n_633),
.Y(n_2403)
);

OAI21x1_ASAP7_75t_L g2404 ( 
.A1(n_2250),
.A2(n_633),
.B(n_634),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_1999),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2328),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2127),
.B(n_634),
.Y(n_2407)
);

BUFx2_ASAP7_75t_L g2408 ( 
.A(n_1953),
.Y(n_2408)
);

INVx1_ASAP7_75t_SL g2409 ( 
.A(n_2240),
.Y(n_2409)
);

OAI21x1_ASAP7_75t_L g2410 ( 
.A1(n_2265),
.A2(n_636),
.B(n_637),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1986),
.Y(n_2411)
);

A2O1A1Ixp33_ASAP7_75t_L g2412 ( 
.A1(n_2252),
.A2(n_637),
.B(n_638),
.C(n_639),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_1986),
.Y(n_2413)
);

NAND2x1_ASAP7_75t_L g2414 ( 
.A(n_1948),
.B(n_640),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_2261),
.Y(n_2415)
);

AOI22xp33_ASAP7_75t_L g2416 ( 
.A1(n_1998),
.A2(n_643),
.B1(n_644),
.B2(n_645),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_1985),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2330),
.Y(n_2418)
);

OAI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2183),
.A2(n_643),
.B1(n_644),
.B2(n_645),
.C(n_646),
.Y(n_2419)
);

OAI22xp33_ASAP7_75t_L g2420 ( 
.A1(n_2137),
.A2(n_647),
.B1(n_648),
.B2(n_649),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1985),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_1972),
.Y(n_2422)
);

AO31x2_ASAP7_75t_L g2423 ( 
.A1(n_1975),
.A2(n_647),
.A3(n_649),
.B(n_650),
.Y(n_2423)
);

OAI21x1_ASAP7_75t_L g2424 ( 
.A1(n_2305),
.A2(n_651),
.B(n_652),
.Y(n_2424)
);

BUFx8_ASAP7_75t_L g2425 ( 
.A(n_2077),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2331),
.Y(n_2426)
);

AOI22xp5_ASAP7_75t_L g2427 ( 
.A1(n_2261),
.A2(n_653),
.B1(n_654),
.B2(n_655),
.Y(n_2427)
);

OAI21x1_ASAP7_75t_SL g2428 ( 
.A1(n_1979),
.A2(n_654),
.B(n_655),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2298),
.B(n_657),
.Y(n_2429)
);

AOI221x1_ASAP7_75t_L g2430 ( 
.A1(n_2193),
.A2(n_657),
.B1(n_659),
.B2(n_660),
.C(n_662),
.Y(n_2430)
);

BUFx2_ASAP7_75t_L g2431 ( 
.A(n_2298),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_1976),
.Y(n_2432)
);

INVx5_ASAP7_75t_L g2433 ( 
.A(n_1948),
.Y(n_2433)
);

OAI21x1_ASAP7_75t_L g2434 ( 
.A1(n_2319),
.A2(n_659),
.B(n_660),
.Y(n_2434)
);

CKINVDCx5p33_ASAP7_75t_R g2435 ( 
.A(n_2238),
.Y(n_2435)
);

OAI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_2254),
.A2(n_662),
.B(n_663),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_1992),
.Y(n_2437)
);

NAND3xp33_ASAP7_75t_L g2438 ( 
.A(n_2079),
.B(n_664),
.C(n_665),
.Y(n_2438)
);

NAND2x1p5_ASAP7_75t_L g2439 ( 
.A(n_2022),
.B(n_664),
.Y(n_2439)
);

OAI22xp5_ASAP7_75t_SL g2440 ( 
.A1(n_2263),
.A2(n_667),
.B1(n_668),
.B2(n_669),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2145),
.B(n_667),
.Y(n_2441)
);

OAI21x1_ASAP7_75t_L g2442 ( 
.A1(n_2322),
.A2(n_668),
.B(n_670),
.Y(n_2442)
);

OAI22xp33_ASAP7_75t_L g2443 ( 
.A1(n_2137),
.A2(n_2258),
.B1(n_2315),
.B2(n_2154),
.Y(n_2443)
);

BUFx10_ASAP7_75t_L g2444 ( 
.A(n_2039),
.Y(n_2444)
);

AOI22xp33_ASAP7_75t_L g2445 ( 
.A1(n_2258),
.A2(n_670),
.B1(n_671),
.B2(n_673),
.Y(n_2445)
);

AOI22xp33_ASAP7_75t_L g2446 ( 
.A1(n_2315),
.A2(n_671),
.B1(n_673),
.B2(n_674),
.Y(n_2446)
);

CKINVDCx20_ASAP7_75t_R g2447 ( 
.A(n_2233),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_1958),
.B(n_674),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2108),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_L g2450 ( 
.A(n_1963),
.B(n_675),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_1967),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2182),
.B(n_677),
.Y(n_2452)
);

AO31x2_ASAP7_75t_L g2453 ( 
.A1(n_2256),
.A2(n_678),
.A3(n_679),
.B(n_681),
.Y(n_2453)
);

OAI21x1_ASAP7_75t_L g2454 ( 
.A1(n_2327),
.A2(n_678),
.B(n_679),
.Y(n_2454)
);

BUFx2_ASAP7_75t_L g2455 ( 
.A(n_2057),
.Y(n_2455)
);

OAI21xp5_ASAP7_75t_L g2456 ( 
.A1(n_2270),
.A2(n_682),
.B(n_683),
.Y(n_2456)
);

NAND2x1p5_ASAP7_75t_L g2457 ( 
.A(n_2205),
.B(n_682),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2002),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1967),
.Y(n_2459)
);

OAI21x1_ASAP7_75t_L g2460 ( 
.A1(n_2329),
.A2(n_684),
.B(n_686),
.Y(n_2460)
);

NAND2x1p5_ASAP7_75t_L g2461 ( 
.A(n_2205),
.B(n_684),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2127),
.B(n_686),
.Y(n_2462)
);

A2O1A1Ixp33_ASAP7_75t_L g2463 ( 
.A1(n_2271),
.A2(n_687),
.B(n_689),
.C(n_690),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2196),
.Y(n_2464)
);

OAI22xp5_ASAP7_75t_L g2465 ( 
.A1(n_1968),
.A2(n_687),
.B1(n_690),
.B2(n_691),
.Y(n_2465)
);

AOI21x1_ASAP7_75t_L g2466 ( 
.A1(n_2041),
.A2(n_691),
.B(n_692),
.Y(n_2466)
);

AO21x2_ASAP7_75t_L g2467 ( 
.A1(n_2264),
.A2(n_2311),
.B(n_2195),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2196),
.Y(n_2468)
);

OAI22xp33_ASAP7_75t_L g2469 ( 
.A1(n_2137),
.A2(n_692),
.B1(n_693),
.B2(n_694),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2047),
.Y(n_2470)
);

AOI21x1_ASAP7_75t_L g2471 ( 
.A1(n_2170),
.A2(n_693),
.B(n_694),
.Y(n_2471)
);

BUFx2_ASAP7_75t_SL g2472 ( 
.A(n_2091),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2200),
.Y(n_2473)
);

OAI21xp33_ASAP7_75t_SL g2474 ( 
.A1(n_1979),
.A2(n_695),
.B(n_696),
.Y(n_2474)
);

AOI22xp33_ASAP7_75t_L g2475 ( 
.A1(n_2036),
.A2(n_698),
.B1(n_700),
.B2(n_701),
.Y(n_2475)
);

NOR2xp33_ASAP7_75t_L g2476 ( 
.A(n_2139),
.B(n_2186),
.Y(n_2476)
);

BUFx3_ASAP7_75t_L g2477 ( 
.A(n_2233),
.Y(n_2477)
);

INVxp67_ASAP7_75t_L g2478 ( 
.A(n_2104),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2200),
.Y(n_2479)
);

BUFx2_ASAP7_75t_L g2480 ( 
.A(n_2062),
.Y(n_2480)
);

BUFx3_ASAP7_75t_L g2481 ( 
.A(n_2014),
.Y(n_2481)
);

OA21x2_ASAP7_75t_L g2482 ( 
.A1(n_2090),
.A2(n_702),
.B(n_703),
.Y(n_2482)
);

OAI21x1_ASAP7_75t_SL g2483 ( 
.A1(n_2237),
.A2(n_702),
.B(n_704),
.Y(n_2483)
);

OAI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_1968),
.A2(n_705),
.B1(n_706),
.B2(n_707),
.Y(n_2484)
);

OAI22xp33_ASAP7_75t_L g2485 ( 
.A1(n_2154),
.A2(n_706),
.B1(n_707),
.B2(n_708),
.Y(n_2485)
);

OA21x2_ASAP7_75t_L g2486 ( 
.A1(n_2198),
.A2(n_708),
.B(n_709),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2049),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_2018),
.Y(n_2488)
);

A2O1A1Ixp33_ASAP7_75t_L g2489 ( 
.A1(n_2272),
.A2(n_709),
.B(n_710),
.C(n_711),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2061),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2205),
.B(n_711),
.Y(n_2491)
);

INVx3_ASAP7_75t_L g2492 ( 
.A(n_2211),
.Y(n_2492)
);

HB1xp67_ASAP7_75t_L g2493 ( 
.A(n_2139),
.Y(n_2493)
);

OAI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_2289),
.A2(n_714),
.B(n_715),
.Y(n_2494)
);

AOI22xp33_ASAP7_75t_L g2495 ( 
.A1(n_2044),
.A2(n_715),
.B1(n_716),
.B2(n_717),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2205),
.B(n_716),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2204),
.Y(n_2497)
);

INVx6_ASAP7_75t_L g2498 ( 
.A(n_2073),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2131),
.B(n_2059),
.Y(n_2499)
);

OR2x6_ASAP7_75t_L g2500 ( 
.A(n_2062),
.B(n_719),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2204),
.Y(n_2501)
);

NAND2xp33_ASAP7_75t_L g2502 ( 
.A(n_1948),
.B(n_721),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2282),
.Y(n_2503)
);

CKINVDCx20_ASAP7_75t_R g2504 ( 
.A(n_2133),
.Y(n_2504)
);

NAND3xp33_ASAP7_75t_L g2505 ( 
.A(n_2079),
.B(n_1993),
.C(n_2003),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2214),
.Y(n_2506)
);

OAI21xp5_ASAP7_75t_L g2507 ( 
.A1(n_2291),
.A2(n_722),
.B(n_723),
.Y(n_2507)
);

AO21x2_ASAP7_75t_L g2508 ( 
.A1(n_2237),
.A2(n_722),
.B(n_725),
.Y(n_2508)
);

OAI22xp5_ASAP7_75t_L g2509 ( 
.A1(n_2214),
.A2(n_725),
.B1(n_726),
.B2(n_727),
.Y(n_2509)
);

AOI21x1_ASAP7_75t_L g2510 ( 
.A1(n_2142),
.A2(n_726),
.B(n_728),
.Y(n_2510)
);

NOR2xp33_ASAP7_75t_L g2511 ( 
.A(n_2035),
.B(n_728),
.Y(n_2511)
);

AOI22xp33_ASAP7_75t_L g2512 ( 
.A1(n_2044),
.A2(n_2160),
.B1(n_2173),
.B2(n_1988),
.Y(n_2512)
);

OAI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2215),
.A2(n_729),
.B1(n_731),
.B2(n_733),
.Y(n_2513)
);

OAI21x1_ASAP7_75t_L g2514 ( 
.A1(n_2118),
.A2(n_731),
.B(n_733),
.Y(n_2514)
);

OAI21x1_ASAP7_75t_L g2515 ( 
.A1(n_2021),
.A2(n_734),
.B(n_735),
.Y(n_2515)
);

AND2x4_ASAP7_75t_L g2516 ( 
.A(n_2317),
.B(n_1978),
.Y(n_2516)
);

OAI21x1_ASAP7_75t_L g2517 ( 
.A1(n_2026),
.A2(n_736),
.B(n_737),
.Y(n_2517)
);

OAI22xp5_ASAP7_75t_L g2518 ( 
.A1(n_2215),
.A2(n_736),
.B1(n_737),
.B2(n_741),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2219),
.Y(n_2519)
);

O2A1O1Ixp33_ASAP7_75t_SL g2520 ( 
.A1(n_1952),
.A2(n_2201),
.B(n_2257),
.C(n_2243),
.Y(n_2520)
);

INVx3_ASAP7_75t_L g2521 ( 
.A(n_2317),
.Y(n_2521)
);

AOI21x1_ASAP7_75t_L g2522 ( 
.A1(n_2142),
.A2(n_741),
.B(n_742),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2219),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2221),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2024),
.A2(n_2183),
.B(n_1980),
.Y(n_2525)
);

OAI21xp5_ASAP7_75t_L g2526 ( 
.A1(n_2292),
.A2(n_744),
.B(n_745),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2107),
.B(n_744),
.Y(n_2527)
);

AO21x2_ASAP7_75t_L g2528 ( 
.A1(n_2255),
.A2(n_746),
.B(n_747),
.Y(n_2528)
);

INVx1_ASAP7_75t_SL g2529 ( 
.A(n_2101),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2087),
.B(n_746),
.Y(n_2530)
);

OAI21xp5_ASAP7_75t_L g2531 ( 
.A1(n_2333),
.A2(n_2339),
.B(n_2335),
.Y(n_2531)
);

OAI21xp5_ASAP7_75t_L g2532 ( 
.A1(n_2221),
.A2(n_747),
.B(n_748),
.Y(n_2532)
);

AND2x4_ASAP7_75t_L g2533 ( 
.A(n_1978),
.B(n_749),
.Y(n_2533)
);

CKINVDCx20_ASAP7_75t_R g2534 ( 
.A(n_2070),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2172),
.B(n_750),
.Y(n_2535)
);

AOI22xp33_ASAP7_75t_L g2536 ( 
.A1(n_2160),
.A2(n_751),
.B1(n_753),
.B2(n_754),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2225),
.Y(n_2537)
);

OR2x2_ASAP7_75t_L g2538 ( 
.A(n_2062),
.B(n_754),
.Y(n_2538)
);

OA21x2_ASAP7_75t_L g2539 ( 
.A1(n_2019),
.A2(n_2280),
.B(n_2255),
.Y(n_2539)
);

CKINVDCx20_ASAP7_75t_R g2540 ( 
.A(n_2209),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_2173),
.A2(n_756),
.B1(n_757),
.B2(n_758),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_SL g2542 ( 
.A(n_2222),
.B(n_762),
.Y(n_2542)
);

OAI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_1981),
.A2(n_763),
.B1(n_765),
.B2(n_766),
.Y(n_2543)
);

AO21x2_ASAP7_75t_L g2544 ( 
.A1(n_2280),
.A2(n_766),
.B(n_767),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_2301),
.Y(n_2545)
);

OAI21x1_ASAP7_75t_L g2546 ( 
.A1(n_2037),
.A2(n_768),
.B(n_2110),
.Y(n_2546)
);

OA21x2_ASAP7_75t_L g2547 ( 
.A1(n_2283),
.A2(n_2310),
.B(n_2303),
.Y(n_2547)
);

BUFx8_ASAP7_75t_L g2548 ( 
.A(n_2216),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2172),
.B(n_2225),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_1996),
.Y(n_2550)
);

OAI22xp33_ASAP7_75t_L g2551 ( 
.A1(n_1984),
.A2(n_2210),
.B1(n_2235),
.B2(n_2220),
.Y(n_2551)
);

O2A1O1Ixp5_ASAP7_75t_SL g2552 ( 
.A1(n_2193),
.A2(n_2184),
.B(n_2299),
.C(n_2234),
.Y(n_2552)
);

O2A1O1Ixp33_ASAP7_75t_L g2553 ( 
.A1(n_2156),
.A2(n_2034),
.B(n_1974),
.C(n_2067),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2232),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2239),
.Y(n_2555)
);

INVxp67_ASAP7_75t_SL g2556 ( 
.A(n_2192),
.Y(n_2556)
);

OAI22xp5_ASAP7_75t_L g2557 ( 
.A1(n_2239),
.A2(n_2268),
.B1(n_2273),
.B2(n_2248),
.Y(n_2557)
);

OA21x2_ASAP7_75t_L g2558 ( 
.A1(n_2283),
.A2(n_2310),
.B(n_2303),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2248),
.B(n_2268),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2273),
.Y(n_2560)
);

AND2x4_ASAP7_75t_L g2561 ( 
.A(n_2151),
.B(n_2035),
.Y(n_2561)
);

A2O1A1Ixp33_ASAP7_75t_L g2562 ( 
.A1(n_1983),
.A2(n_1980),
.B(n_2199),
.C(n_2336),
.Y(n_2562)
);

NAND3xp33_ASAP7_75t_SL g2563 ( 
.A(n_2338),
.B(n_2281),
.C(n_2222),
.Y(n_2563)
);

HB1xp67_ASAP7_75t_L g2564 ( 
.A(n_1991),
.Y(n_2564)
);

BUFx3_ASAP7_75t_L g2565 ( 
.A(n_2297),
.Y(n_2565)
);

BUFx6f_ASAP7_75t_L g2566 ( 
.A(n_1949),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2188),
.Y(n_2567)
);

INVx6_ASAP7_75t_L g2568 ( 
.A(n_2073),
.Y(n_2568)
);

AOI22xp33_ASAP7_75t_SL g2569 ( 
.A1(n_2210),
.A2(n_2235),
.B1(n_2241),
.B2(n_2220),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2275),
.Y(n_2570)
);

OAI21xp5_ASAP7_75t_L g2571 ( 
.A1(n_2276),
.A2(n_2293),
.B(n_2279),
.Y(n_2571)
);

AND2x4_ASAP7_75t_L g2572 ( 
.A(n_1964),
.B(n_2098),
.Y(n_2572)
);

AO21x1_ASAP7_75t_L g2573 ( 
.A1(n_2179),
.A2(n_2147),
.B(n_1961),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2213),
.B(n_2218),
.Y(n_2574)
);

INVx3_ASAP7_75t_L g2575 ( 
.A(n_1996),
.Y(n_2575)
);

AO31x2_ASAP7_75t_L g2576 ( 
.A1(n_2086),
.A2(n_2054),
.A3(n_2089),
.B(n_2260),
.Y(n_2576)
);

AOI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2029),
.A2(n_2088),
.B1(n_2244),
.B2(n_2230),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2279),
.Y(n_2578)
);

OAI21x1_ASAP7_75t_SL g2579 ( 
.A1(n_2116),
.A2(n_1960),
.B(n_2136),
.Y(n_2579)
);

AND2x4_ASAP7_75t_L g2580 ( 
.A(n_1964),
.B(n_2098),
.Y(n_2580)
);

NOR2xp67_ASAP7_75t_SL g2581 ( 
.A(n_2136),
.B(n_2066),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2293),
.Y(n_2582)
);

HB1xp67_ASAP7_75t_L g2583 ( 
.A(n_1991),
.Y(n_2583)
);

OA21x2_ASAP7_75t_L g2584 ( 
.A1(n_2033),
.A2(n_2075),
.B(n_2015),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2294),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2294),
.B(n_2300),
.Y(n_2586)
);

OAI21xp5_ASAP7_75t_L g2587 ( 
.A1(n_2300),
.A2(n_2307),
.B(n_2306),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2306),
.B(n_2307),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2308),
.Y(n_2589)
);

OAI21xp5_ASAP7_75t_L g2590 ( 
.A1(n_2308),
.A2(n_2312),
.B(n_2309),
.Y(n_2590)
);

OAI21x1_ASAP7_75t_L g2591 ( 
.A1(n_2075),
.A2(n_1982),
.B(n_2013),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2309),
.Y(n_2592)
);

OA21x2_ASAP7_75t_L g2593 ( 
.A1(n_2033),
.A2(n_2284),
.B(n_2159),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2316),
.Y(n_2594)
);

CKINVDCx8_ASAP7_75t_R g2595 ( 
.A(n_2119),
.Y(n_2595)
);

AND2x2_ASAP7_75t_SL g2596 ( 
.A(n_2249),
.B(n_2266),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_2129),
.B(n_2063),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2134),
.Y(n_2598)
);

NOR2xp33_ASAP7_75t_L g2599 ( 
.A(n_2085),
.B(n_2106),
.Y(n_2599)
);

AO31x2_ASAP7_75t_L g2600 ( 
.A1(n_2267),
.A2(n_2179),
.A3(n_2115),
.B(n_2096),
.Y(n_2600)
);

OAI21xp5_ASAP7_75t_L g2601 ( 
.A1(n_2005),
.A2(n_2007),
.B(n_2031),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2249),
.Y(n_2602)
);

O2A1O1Ixp33_ASAP7_75t_SL g2603 ( 
.A1(n_2120),
.A2(n_2105),
.B(n_2124),
.C(n_2176),
.Y(n_2603)
);

AOI221xp5_ASAP7_75t_L g2604 ( 
.A1(n_2156),
.A2(n_2100),
.B1(n_2277),
.B2(n_2325),
.C(n_2241),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2130),
.B(n_2155),
.Y(n_2605)
);

OAI21xp5_ASAP7_75t_L g2606 ( 
.A1(n_2005),
.A2(n_2007),
.B(n_2031),
.Y(n_2606)
);

NOR2xp33_ASAP7_75t_L g2607 ( 
.A(n_2178),
.B(n_2158),
.Y(n_2607)
);

AO31x2_ASAP7_75t_L g2608 ( 
.A1(n_2169),
.A2(n_2140),
.A3(n_2325),
.B(n_2277),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2082),
.Y(n_2609)
);

INVx5_ASAP7_75t_L g2610 ( 
.A(n_2093),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2266),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2246),
.Y(n_2612)
);

BUFx2_ASAP7_75t_L g2613 ( 
.A(n_2119),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2246),
.Y(n_2614)
);

OR2x2_ASAP7_75t_L g2615 ( 
.A(n_2313),
.B(n_2321),
.Y(n_2615)
);

OAI21xp5_ASAP7_75t_L g2616 ( 
.A1(n_2092),
.A2(n_2337),
.B(n_1951),
.Y(n_2616)
);

OAI21x1_ASAP7_75t_SL g2617 ( 
.A1(n_1960),
.A2(n_2097),
.B(n_2147),
.Y(n_2617)
);

INVx1_ASAP7_75t_SL g2618 ( 
.A(n_2152),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2251),
.Y(n_2619)
);

NOR2xp67_ASAP7_75t_L g2620 ( 
.A(n_2212),
.B(n_2290),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_2302),
.Y(n_2621)
);

OAI211xp5_ASAP7_75t_L g2622 ( 
.A1(n_2016),
.A2(n_2053),
.B(n_2032),
.C(n_2067),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2251),
.Y(n_2623)
);

CKINVDCx6p67_ASAP7_75t_R g2624 ( 
.A(n_2119),
.Y(n_2624)
);

OAI22xp5_ASAP7_75t_L g2625 ( 
.A1(n_2281),
.A2(n_2338),
.B1(n_2320),
.B2(n_2192),
.Y(n_2625)
);

OAI21xp5_ASAP7_75t_L g2626 ( 
.A1(n_2092),
.A2(n_2155),
.B(n_2130),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2334),
.B(n_2074),
.Y(n_2627)
);

AO31x2_ASAP7_75t_L g2628 ( 
.A1(n_2169),
.A2(n_2140),
.A3(n_2071),
.B(n_2181),
.Y(n_2628)
);

OR2x2_ASAP7_75t_L g2629 ( 
.A(n_2174),
.B(n_2065),
.Y(n_2629)
);

AND2x4_ASAP7_75t_L g2630 ( 
.A(n_2010),
.B(n_2023),
.Y(n_2630)
);

OA21x2_ASAP7_75t_L g2631 ( 
.A1(n_2164),
.A2(n_2157),
.B(n_2177),
.Y(n_2631)
);

AOI22xp5_ASAP7_75t_L g2632 ( 
.A1(n_2141),
.A2(n_2126),
.B1(n_2269),
.B2(n_2262),
.Y(n_2632)
);

INVx5_ASAP7_75t_L g2633 ( 
.A(n_2093),
.Y(n_2633)
);

AOI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2165),
.A2(n_1994),
.B1(n_2053),
.B2(n_2051),
.Y(n_2634)
);

HB1xp67_ASAP7_75t_L g2635 ( 
.A(n_2152),
.Y(n_2635)
);

OR2x2_ASAP7_75t_L g2636 ( 
.A(n_2318),
.B(n_2323),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2119),
.Y(n_2637)
);

NAND3xp33_ASAP7_75t_L g2638 ( 
.A(n_2080),
.B(n_2177),
.C(n_2012),
.Y(n_2638)
);

NAND2xp33_ASAP7_75t_SL g2639 ( 
.A(n_2051),
.B(n_2192),
.Y(n_2639)
);

AO31x2_ASAP7_75t_L g2640 ( 
.A1(n_2181),
.A2(n_2112),
.A3(n_2122),
.B(n_2125),
.Y(n_2640)
);

OR2x6_ASAP7_75t_L g2641 ( 
.A(n_2114),
.B(n_2175),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2109),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2180),
.B(n_1956),
.Y(n_2643)
);

OAI21xp5_ASAP7_75t_L g2644 ( 
.A1(n_2042),
.A2(n_2050),
.B(n_2048),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2180),
.B(n_1956),
.Y(n_2645)
);

OR2x2_ASAP7_75t_L g2646 ( 
.A(n_2102),
.B(n_2187),
.Y(n_2646)
);

NOR2xp67_ASAP7_75t_L g2647 ( 
.A(n_2191),
.B(n_1959),
.Y(n_2647)
);

AOI221xp5_ASAP7_75t_SL g2648 ( 
.A1(n_1977),
.A2(n_2113),
.B1(n_2094),
.B2(n_2121),
.C(n_2150),
.Y(n_2648)
);

A2O1A1Ixp33_ASAP7_75t_L g2649 ( 
.A1(n_2149),
.A2(n_2161),
.B(n_2185),
.C(n_2020),
.Y(n_2649)
);

INVx2_ASAP7_75t_SL g2650 ( 
.A(n_2152),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2056),
.B(n_2068),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2109),
.Y(n_2652)
);

AOI22xp33_ASAP7_75t_SL g2653 ( 
.A1(n_2166),
.A2(n_2043),
.B1(n_2144),
.B2(n_2175),
.Y(n_2653)
);

AOI21xp5_ASAP7_75t_L g2654 ( 
.A1(n_2168),
.A2(n_2171),
.B(n_2143),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2112),
.Y(n_2655)
);

OAI22xp33_ASAP7_75t_L g2656 ( 
.A1(n_1994),
.A2(n_2165),
.B1(n_2163),
.B2(n_2048),
.Y(n_2656)
);

OAI21x1_ASAP7_75t_L g2657 ( 
.A1(n_2122),
.A2(n_2125),
.B(n_2084),
.Y(n_2657)
);

BUFx2_ASAP7_75t_L g2658 ( 
.A(n_2008),
.Y(n_2658)
);

O2A1O1Ixp33_ASAP7_75t_L g2659 ( 
.A1(n_2234),
.A2(n_2299),
.B(n_2042),
.C(n_2050),
.Y(n_2659)
);

OAI21x1_ASAP7_75t_L g2660 ( 
.A1(n_1989),
.A2(n_1995),
.B(n_2228),
.Y(n_2660)
);

OAI21x1_ASAP7_75t_L g2661 ( 
.A1(n_2223),
.A2(n_2023),
.B(n_2028),
.Y(n_2661)
);

OAI21x1_ASAP7_75t_L g2662 ( 
.A1(n_2045),
.A2(n_2153),
.B(n_2072),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2082),
.Y(n_2663)
);

OAI21xp5_ASAP7_75t_L g2664 ( 
.A1(n_2045),
.A2(n_2194),
.B(n_2190),
.Y(n_2664)
);

INVx4_ASAP7_75t_L g2665 ( 
.A(n_2103),
.Y(n_2665)
);

AOI22xp33_ASAP7_75t_L g2666 ( 
.A1(n_2043),
.A2(n_2076),
.B1(n_2190),
.B2(n_2191),
.Y(n_2666)
);

INVx4_ASAP7_75t_L g2667 ( 
.A(n_2103),
.Y(n_2667)
);

AO21x2_ASAP7_75t_L g2668 ( 
.A1(n_2217),
.A2(n_2078),
.B(n_2224),
.Y(n_2668)
);

AO21x1_ASAP7_75t_L g2669 ( 
.A1(n_2011),
.A2(n_1997),
.B(n_2144),
.Y(n_2669)
);

NOR2x1_ASAP7_75t_SL g2670 ( 
.A(n_1971),
.B(n_2202),
.Y(n_2670)
);

AOI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2217),
.A2(n_2078),
.B1(n_2095),
.B2(n_2148),
.Y(n_2671)
);

AOI332xp33_ASAP7_75t_L g2672 ( 
.A1(n_1997),
.A2(n_2011),
.A3(n_2009),
.B1(n_2069),
.B2(n_2064),
.B3(n_2326),
.C1(n_2227),
.C2(n_2253),
.Y(n_2672)
);

OAI21x1_ASAP7_75t_L g2673 ( 
.A1(n_2202),
.A2(n_2111),
.B(n_1956),
.Y(n_2673)
);

BUFx3_ASAP7_75t_L g2674 ( 
.A(n_2117),
.Y(n_2674)
);

AND2x4_ASAP7_75t_L g2675 ( 
.A(n_2117),
.B(n_2148),
.Y(n_2675)
);

BUFx2_ASAP7_75t_R g2676 ( 
.A(n_1997),
.Y(n_2676)
);

HB1xp67_ASAP7_75t_L g2677 ( 
.A(n_2111),
.Y(n_2677)
);

CKINVDCx9p33_ASAP7_75t_R g2678 ( 
.A(n_2011),
.Y(n_2678)
);

OAI221xp5_ASAP7_75t_L g2679 ( 
.A1(n_2117),
.A2(n_2148),
.B1(n_2009),
.B2(n_2001),
.C(n_1987),
.Y(n_2679)
);

NOR3xp33_ASAP7_75t_L g2680 ( 
.A(n_2009),
.B(n_2069),
.C(n_2001),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2138),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2138),
.Y(n_2682)
);

O2A1O1Ixp33_ASAP7_75t_SL g2683 ( 
.A1(n_1987),
.A2(n_2001),
.B(n_2006),
.C(n_2285),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_1987),
.B(n_2006),
.Y(n_2684)
);

BUFx6f_ASAP7_75t_L g2685 ( 
.A(n_2083),
.Y(n_2685)
);

OR2x2_ASAP7_75t_L g2686 ( 
.A(n_2385),
.B(n_2138),
.Y(n_2686)
);

AOI221xp5_ASAP7_75t_L g2687 ( 
.A1(n_2551),
.A2(n_2006),
.B1(n_2146),
.B2(n_2083),
.C(n_2227),
.Y(n_2687)
);

INVx3_ASAP7_75t_L g2688 ( 
.A(n_2365),
.Y(n_2688)
);

HB1xp67_ASAP7_75t_L g2689 ( 
.A(n_2493),
.Y(n_2689)
);

OAI21x1_ASAP7_75t_L g2690 ( 
.A1(n_2673),
.A2(n_2146),
.B(n_2167),
.Y(n_2690)
);

INVx2_ASAP7_75t_SL g2691 ( 
.A(n_2425),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2347),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2347),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2478),
.B(n_2146),
.Y(n_2694)
);

INVx3_ASAP7_75t_L g2695 ( 
.A(n_2365),
.Y(n_2695)
);

INVx3_ASAP7_75t_SL g2696 ( 
.A(n_2447),
.Y(n_2696)
);

HB1xp67_ASAP7_75t_L g2697 ( 
.A(n_2493),
.Y(n_2697)
);

INVx2_ASAP7_75t_SL g2698 ( 
.A(n_2425),
.Y(n_2698)
);

INVx3_ASAP7_75t_L g2699 ( 
.A(n_2395),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2574),
.B(n_2357),
.Y(n_2700)
);

HB1xp67_ASAP7_75t_L g2701 ( 
.A(n_2357),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2499),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_L g2703 ( 
.A(n_2478),
.B(n_2167),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2499),
.Y(n_2704)
);

INVx3_ASAP7_75t_L g2705 ( 
.A(n_2395),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2345),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_L g2707 ( 
.A1(n_2604),
.A2(n_2167),
.B1(n_2569),
.B2(n_2551),
.Y(n_2707)
);

OAI21xp5_ASAP7_75t_L g2708 ( 
.A1(n_2552),
.A2(n_2562),
.B(n_2525),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2349),
.Y(n_2709)
);

OR2x6_ASAP7_75t_L g2710 ( 
.A(n_2500),
.B(n_2613),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2354),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2415),
.B(n_2596),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2361),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2343),
.B(n_2399),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2364),
.Y(n_2715)
);

INVx2_ASAP7_75t_SL g2716 ( 
.A(n_2477),
.Y(n_2716)
);

HB1xp67_ASAP7_75t_L g2717 ( 
.A(n_2415),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_L g2718 ( 
.A1(n_2604),
.A2(n_2569),
.B1(n_2443),
.B2(n_2512),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2386),
.B(n_2612),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2595),
.Y(n_2720)
);

AOI22xp33_ASAP7_75t_L g2721 ( 
.A1(n_2443),
.A2(n_2512),
.B1(n_2355),
.B2(n_2614),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2368),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2369),
.Y(n_2723)
);

INVx2_ASAP7_75t_SL g2724 ( 
.A(n_2548),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2386),
.B(n_2619),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2409),
.B(n_2431),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2677),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2370),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_2624),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2409),
.B(n_2429),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2373),
.Y(n_2731)
);

INVx1_ASAP7_75t_SL g2732 ( 
.A(n_2455),
.Y(n_2732)
);

BUFx2_ASAP7_75t_L g2733 ( 
.A(n_2480),
.Y(n_2733)
);

NAND2x1p5_ASAP7_75t_L g2734 ( 
.A(n_2381),
.B(n_2433),
.Y(n_2734)
);

BUFx3_ASAP7_75t_L g2735 ( 
.A(n_2561),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2384),
.Y(n_2736)
);

OAI22xp5_ASAP7_75t_L g2737 ( 
.A1(n_2577),
.A2(n_2615),
.B1(n_2500),
.B2(n_2340),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2402),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2405),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2356),
.Y(n_2740)
);

AO31x2_ASAP7_75t_L g2741 ( 
.A1(n_2669),
.A2(n_2684),
.A3(n_2609),
.B(n_2663),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2356),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2367),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2367),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2530),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2530),
.Y(n_2746)
);

AO21x1_ASAP7_75t_SL g2747 ( 
.A1(n_2564),
.A2(n_2583),
.B(n_2433),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2394),
.Y(n_2748)
);

CKINVDCx20_ASAP7_75t_R g2749 ( 
.A(n_2383),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2623),
.B(n_2607),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2394),
.Y(n_2751)
);

BUFx3_ASAP7_75t_L g2752 ( 
.A(n_2561),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2441),
.Y(n_2753)
);

BUFx3_ASAP7_75t_L g2754 ( 
.A(n_2548),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2441),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2642),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2452),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2452),
.Y(n_2758)
);

BUFx2_ASAP7_75t_L g2759 ( 
.A(n_2641),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2448),
.B(n_2340),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2351),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2358),
.Y(n_2762)
);

BUFx2_ASAP7_75t_L g2763 ( 
.A(n_2641),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2381),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2652),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2655),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2393),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2529),
.B(n_2500),
.Y(n_2768)
);

BUFx6f_ASAP7_75t_L g2769 ( 
.A(n_2342),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2677),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2398),
.Y(n_2771)
);

INVx2_ASAP7_75t_SL g2772 ( 
.A(n_2498),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2406),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2418),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2582),
.Y(n_2775)
);

INVx2_ASAP7_75t_L g2776 ( 
.A(n_2585),
.Y(n_2776)
);

HB1xp67_ASAP7_75t_L g2777 ( 
.A(n_2549),
.Y(n_2777)
);

INVx3_ASAP7_75t_L g2778 ( 
.A(n_2381),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2426),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2589),
.Y(n_2780)
);

HB1xp67_ASAP7_75t_SL g2781 ( 
.A(n_2625),
.Y(n_2781)
);

BUFx6f_ASAP7_75t_L g2782 ( 
.A(n_2342),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2432),
.Y(n_2783)
);

BUFx4f_ASAP7_75t_SL g2784 ( 
.A(n_2540),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2529),
.B(n_2360),
.Y(n_2785)
);

AOI22xp33_ASAP7_75t_L g2786 ( 
.A1(n_2355),
.A2(n_2359),
.B1(n_2653),
.B2(n_2627),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2437),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2449),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2594),
.Y(n_2789)
);

INVx2_ASAP7_75t_SL g2790 ( 
.A(n_2498),
.Y(n_2790)
);

NAND2x1_ASAP7_75t_L g2791 ( 
.A(n_2625),
.B(n_2665),
.Y(n_2791)
);

INVx1_ASAP7_75t_SL g2792 ( 
.A(n_2472),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2458),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2685),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2685),
.Y(n_2795)
);

BUFx3_ASAP7_75t_L g2796 ( 
.A(n_2610),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2470),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2346),
.B(n_2408),
.Y(n_2798)
);

INVx1_ASAP7_75t_SL g2799 ( 
.A(n_2481),
.Y(n_2799)
);

HB1xp67_ASAP7_75t_L g2800 ( 
.A(n_2549),
.Y(n_2800)
);

BUFx6f_ASAP7_75t_L g2801 ( 
.A(n_2342),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2487),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2490),
.Y(n_2803)
);

NOR2x1_ASAP7_75t_SL g2804 ( 
.A(n_2381),
.B(n_2433),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2346),
.B(n_2629),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2451),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2627),
.B(n_2380),
.Y(n_2807)
);

HB1xp67_ASAP7_75t_L g2808 ( 
.A(n_2564),
.Y(n_2808)
);

AOI21xp5_ASAP7_75t_SL g2809 ( 
.A1(n_2563),
.A2(n_2439),
.B(n_2396),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2380),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2597),
.Y(n_2811)
);

INVx2_ASAP7_75t_SL g2812 ( 
.A(n_2498),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2476),
.B(n_2533),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2459),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2491),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2491),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2496),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2533),
.B(n_2511),
.Y(n_2818)
);

A2O1A1Ixp33_ASAP7_75t_L g2819 ( 
.A1(n_2553),
.A2(n_2474),
.B(n_2659),
.C(n_2352),
.Y(n_2819)
);

AND2x4_ASAP7_75t_L g2820 ( 
.A(n_2433),
.B(n_2637),
.Y(n_2820)
);

AND2x4_ASAP7_75t_L g2821 ( 
.A(n_2675),
.B(n_2610),
.Y(n_2821)
);

A2O1A1Ixp33_ASAP7_75t_L g2822 ( 
.A1(n_2553),
.A2(n_2659),
.B(n_2352),
.C(n_2363),
.Y(n_2822)
);

HB1xp67_ASAP7_75t_L g2823 ( 
.A(n_2583),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2464),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2496),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2468),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2473),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2516),
.B(n_2572),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_2479),
.Y(n_2829)
);

INVx4_ASAP7_75t_L g2830 ( 
.A(n_2545),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2634),
.A2(n_2495),
.B1(n_2653),
.B2(n_2536),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2598),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2602),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_2362),
.Y(n_2834)
);

INVx2_ASAP7_75t_SL g2835 ( 
.A(n_2568),
.Y(n_2835)
);

OAI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2525),
.A2(n_2505),
.B(n_2353),
.Y(n_2836)
);

INVxp67_ASAP7_75t_L g2837 ( 
.A(n_2542),
.Y(n_2837)
);

HB1xp67_ASAP7_75t_L g2838 ( 
.A(n_2535),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2634),
.B(n_2375),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2611),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2497),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2501),
.Y(n_2842)
);

BUFx2_ASAP7_75t_L g2843 ( 
.A(n_2641),
.Y(n_2843)
);

OAI21x1_ASAP7_75t_L g2844 ( 
.A1(n_2664),
.A2(n_2657),
.B(n_2591),
.Y(n_2844)
);

INVx3_ASAP7_75t_L g2845 ( 
.A(n_2362),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2516),
.B(n_2572),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2506),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2465),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2519),
.Y(n_2849)
);

NOR2x1_ASAP7_75t_R g2850 ( 
.A(n_2350),
.B(n_2435),
.Y(n_2850)
);

AND2x4_ASAP7_75t_L g2851 ( 
.A(n_2675),
.B(n_2610),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2465),
.Y(n_2852)
);

CKINVDCx20_ASAP7_75t_R g2853 ( 
.A(n_2534),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2580),
.B(n_2388),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2484),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2484),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2396),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2439),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2457),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2523),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2457),
.Y(n_2861)
);

INVx3_ASAP7_75t_L g2862 ( 
.A(n_2492),
.Y(n_2862)
);

BUFx6f_ASAP7_75t_L g2863 ( 
.A(n_2387),
.Y(n_2863)
);

INVx3_ASAP7_75t_L g2864 ( 
.A(n_2492),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2524),
.Y(n_2865)
);

HB1xp67_ASAP7_75t_L g2866 ( 
.A(n_2535),
.Y(n_2866)
);

BUFx2_ASAP7_75t_L g2867 ( 
.A(n_2568),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2580),
.B(n_2388),
.Y(n_2868)
);

OAI21x1_ASAP7_75t_L g2869 ( 
.A1(n_2389),
.A2(n_2382),
.B(n_2510),
.Y(n_2869)
);

INVx2_ASAP7_75t_SL g2870 ( 
.A(n_2568),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2461),
.Y(n_2871)
);

AND2x2_ASAP7_75t_L g2872 ( 
.A(n_2538),
.B(n_2527),
.Y(n_2872)
);

AOI22xp5_ASAP7_75t_L g2873 ( 
.A1(n_2651),
.A2(n_2407),
.B1(n_2632),
.B2(n_2527),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2461),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2509),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2537),
.Y(n_2876)
);

INVx2_ASAP7_75t_SL g2877 ( 
.A(n_2444),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2509),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2513),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2513),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2518),
.Y(n_2881)
);

HB1xp67_ASAP7_75t_L g2882 ( 
.A(n_2556),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2407),
.B(n_2599),
.Y(n_2883)
);

INVx2_ASAP7_75t_SL g2884 ( 
.A(n_2444),
.Y(n_2884)
);

OA21x2_ASAP7_75t_L g2885 ( 
.A1(n_2684),
.A2(n_2682),
.B(n_2681),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2518),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2554),
.Y(n_2887)
);

INVxp33_ASAP7_75t_L g2888 ( 
.A(n_2635),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2348),
.Y(n_2889)
);

BUFx3_ASAP7_75t_L g2890 ( 
.A(n_2610),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2555),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2560),
.Y(n_2892)
);

BUFx2_ASAP7_75t_L g2893 ( 
.A(n_2674),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2348),
.Y(n_2894)
);

BUFx10_ASAP7_75t_L g2895 ( 
.A(n_2503),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2403),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2379),
.B(n_2391),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2570),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2515),
.Y(n_2899)
);

NAND2x1p5_ASAP7_75t_L g2900 ( 
.A(n_2633),
.B(n_2414),
.Y(n_2900)
);

INVx2_ASAP7_75t_SL g2901 ( 
.A(n_2488),
.Y(n_2901)
);

AOI21x1_ASAP7_75t_L g2902 ( 
.A1(n_2522),
.A2(n_2581),
.B(n_2654),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2578),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2592),
.Y(n_2904)
);

HB1xp67_ASAP7_75t_L g2905 ( 
.A(n_2556),
.Y(n_2905)
);

AOI22xp33_ASAP7_75t_L g2906 ( 
.A1(n_2359),
.A2(n_2573),
.B1(n_2543),
.B2(n_2495),
.Y(n_2906)
);

CKINVDCx6p67_ASAP7_75t_R g2907 ( 
.A(n_2504),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2517),
.Y(n_2908)
);

INVx3_ASAP7_75t_L g2909 ( 
.A(n_2633),
.Y(n_2909)
);

INVx5_ASAP7_75t_L g2910 ( 
.A(n_2633),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2411),
.Y(n_2911)
);

OAI22xp5_ASAP7_75t_L g2912 ( 
.A1(n_2536),
.A2(n_2541),
.B1(n_2666),
.B2(n_2469),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2413),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2532),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_2633),
.Y(n_2915)
);

AND2x2_ASAP7_75t_L g2916 ( 
.A(n_2450),
.B(n_2416),
.Y(n_2916)
);

OR2x2_ASAP7_75t_L g2917 ( 
.A(n_2646),
.B(n_2605),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2532),
.Y(n_2918)
);

HB1xp67_ASAP7_75t_L g2919 ( 
.A(n_2640),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2416),
.B(n_2462),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2521),
.B(n_2445),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2622),
.B(n_2400),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2371),
.Y(n_2923)
);

OAI21x1_ASAP7_75t_L g2924 ( 
.A1(n_2546),
.A2(n_2514),
.B(n_2661),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2417),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2521),
.B(n_2445),
.Y(n_2926)
);

INVx4_ASAP7_75t_L g2927 ( 
.A(n_2621),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2421),
.Y(n_2928)
);

INVx3_ASAP7_75t_L g2929 ( 
.A(n_2665),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2387),
.Y(n_2930)
);

OAI21x1_ASAP7_75t_L g2931 ( 
.A1(n_2531),
.A2(n_2645),
.B(n_2643),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2387),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2372),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2566),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2605),
.B(n_2422),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2566),
.Y(n_2936)
);

BUFx3_ASAP7_75t_L g2937 ( 
.A(n_2565),
.Y(n_2937)
);

INVx3_ASAP7_75t_L g2938 ( 
.A(n_2667),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2566),
.Y(n_2939)
);

BUFx4f_ASAP7_75t_SL g2940 ( 
.A(n_2667),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2374),
.Y(n_2941)
);

HB1xp67_ASAP7_75t_L g2942 ( 
.A(n_2640),
.Y(n_2942)
);

CKINVDCx5p33_ASAP7_75t_R g2943 ( 
.A(n_2567),
.Y(n_2943)
);

OR2x6_ASAP7_75t_L g2944 ( 
.A(n_2647),
.B(n_2579),
.Y(n_2944)
);

INVx2_ASAP7_75t_SL g2945 ( 
.A(n_2636),
.Y(n_2945)
);

OAI21xp33_ASAP7_75t_SL g2946 ( 
.A1(n_2363),
.A2(n_2586),
.B(n_2559),
.Y(n_2946)
);

OR2x6_ASAP7_75t_L g2947 ( 
.A(n_2658),
.B(n_2630),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2378),
.Y(n_2948)
);

OAI21x1_ASAP7_75t_L g2949 ( 
.A1(n_2531),
.A2(n_2645),
.B(n_2643),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_2630),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2543),
.A2(n_2469),
.B1(n_2420),
.B2(n_2485),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2446),
.B(n_2635),
.Y(n_2952)
);

INVx3_ASAP7_75t_L g2953 ( 
.A(n_2550),
.Y(n_2953)
);

NAND2x1p5_ASAP7_75t_L g2954 ( 
.A(n_2618),
.B(n_2620),
.Y(n_2954)
);

OR2x2_ASAP7_75t_L g2955 ( 
.A(n_2650),
.B(n_2559),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2404),
.Y(n_2956)
);

AOI22xp33_ASAP7_75t_L g2957 ( 
.A1(n_2420),
.A2(n_2485),
.B1(n_2446),
.B2(n_2541),
.Y(n_2957)
);

AND2x4_ASAP7_75t_L g2958 ( 
.A(n_2644),
.B(n_2670),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2410),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2608),
.B(n_2618),
.Y(n_2960)
);

NAND2x1_ASAP7_75t_L g2961 ( 
.A(n_2483),
.B(n_2390),
.Y(n_2961)
);

INVx3_ASAP7_75t_L g2962 ( 
.A(n_2550),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2424),
.Y(n_2963)
);

INVx2_ASAP7_75t_SL g2964 ( 
.A(n_2575),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2434),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2442),
.Y(n_2966)
);

OAI21x1_ASAP7_75t_L g2967 ( 
.A1(n_2601),
.A2(n_2606),
.B(n_2539),
.Y(n_2967)
);

BUFx2_ASAP7_75t_SL g2968 ( 
.A(n_2575),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2454),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2460),
.Y(n_2970)
);

HB1xp67_ASAP7_75t_L g2971 ( 
.A(n_2640),
.Y(n_2971)
);

HB1xp67_ASAP7_75t_L g2972 ( 
.A(n_2547),
.Y(n_2972)
);

CKINVDCx5p33_ASAP7_75t_R g2973 ( 
.A(n_2440),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2423),
.Y(n_2974)
);

INVx4_ASAP7_75t_SL g2975 ( 
.A(n_2608),
.Y(n_2975)
);

INVx1_ASAP7_75t_SL g2976 ( 
.A(n_2502),
.Y(n_2976)
);

OR2x2_ASAP7_75t_L g2977 ( 
.A(n_2586),
.B(n_2588),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2608),
.B(n_2376),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2423),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2423),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2453),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2706),
.Y(n_2982)
);

BUFx3_ASAP7_75t_L g2983 ( 
.A(n_2940),
.Y(n_2983)
);

BUFx6f_ASAP7_75t_L g2984 ( 
.A(n_2734),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2709),
.Y(n_2985)
);

AND2x2_ASAP7_75t_L g2986 ( 
.A(n_2960),
.B(n_2680),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2975),
.B(n_2680),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2975),
.B(n_2453),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2711),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2713),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2700),
.B(n_2427),
.Y(n_2991)
);

AND2x4_ASAP7_75t_L g2992 ( 
.A(n_2958),
.B(n_2601),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2805),
.B(n_2475),
.Y(n_2993)
);

INVx1_ASAP7_75t_SL g2994 ( 
.A(n_2792),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2760),
.B(n_2475),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2730),
.B(n_2666),
.Y(n_2996)
);

AND2x4_ASAP7_75t_L g2997 ( 
.A(n_2958),
.B(n_2606),
.Y(n_2997)
);

AND2x2_ASAP7_75t_L g2998 ( 
.A(n_2726),
.B(n_2542),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2715),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2737),
.B(n_2622),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2722),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2723),
.Y(n_3002)
);

INVx3_ASAP7_75t_SL g3003 ( 
.A(n_2696),
.Y(n_3003)
);

INVx3_ASAP7_75t_L g3004 ( 
.A(n_2734),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2813),
.B(n_2453),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2728),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2818),
.B(n_2397),
.Y(n_3007)
);

HB1xp67_ASAP7_75t_L g3008 ( 
.A(n_2882),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2798),
.B(n_2397),
.Y(n_3009)
);

INVxp67_ASAP7_75t_L g3010 ( 
.A(n_2727),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2702),
.B(n_2588),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_2883),
.B(n_2401),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2872),
.B(n_2401),
.Y(n_3013)
);

BUFx2_ASAP7_75t_L g3014 ( 
.A(n_2940),
.Y(n_3014)
);

AND2x2_ASAP7_75t_L g3015 ( 
.A(n_2811),
.B(n_2436),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2945),
.B(n_2436),
.Y(n_3016)
);

BUFx3_ASAP7_75t_L g3017 ( 
.A(n_2910),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2731),
.Y(n_3018)
);

INVxp67_ASAP7_75t_L g3019 ( 
.A(n_2727),
.Y(n_3019)
);

HB1xp67_ASAP7_75t_L g3020 ( 
.A(n_2882),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2718),
.B(n_2456),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2736),
.Y(n_3022)
);

OAI221xp5_ASAP7_75t_L g3023 ( 
.A1(n_2718),
.A2(n_2626),
.B1(n_2419),
.B2(n_2671),
.C(n_2654),
.Y(n_3023)
);

AND2x2_ASAP7_75t_L g3024 ( 
.A(n_2828),
.B(n_2456),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2738),
.Y(n_3025)
);

AND2x2_ASAP7_75t_L g3026 ( 
.A(n_2846),
.B(n_2494),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2785),
.B(n_2557),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2712),
.B(n_2494),
.Y(n_3028)
);

AND2x4_ASAP7_75t_L g3029 ( 
.A(n_2958),
.B(n_2644),
.Y(n_3029)
);

HB1xp67_ASAP7_75t_L g3030 ( 
.A(n_2905),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2739),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2704),
.Y(n_3032)
);

INVxp67_ASAP7_75t_L g3033 ( 
.A(n_2770),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2917),
.B(n_2557),
.Y(n_3034)
);

AND2x2_ASAP7_75t_L g3035 ( 
.A(n_2768),
.B(n_2507),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2761),
.Y(n_3036)
);

OR2x2_ASAP7_75t_L g3037 ( 
.A(n_2732),
.B(n_2419),
.Y(n_3037)
);

INVx4_ASAP7_75t_L g3038 ( 
.A(n_2910),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2762),
.Y(n_3039)
);

OR2x2_ASAP7_75t_L g3040 ( 
.A(n_2701),
.B(n_2679),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2767),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2701),
.B(n_2507),
.Y(n_3042)
);

AND2x4_ASAP7_75t_L g3043 ( 
.A(n_2975),
.B(n_2467),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2692),
.B(n_2626),
.Y(n_3044)
);

NOR2xp67_ASAP7_75t_L g3045 ( 
.A(n_2910),
.B(n_2563),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2717),
.B(n_2526),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_2717),
.B(n_2526),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2854),
.B(n_2868),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2735),
.B(n_2377),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2735),
.B(n_2377),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2771),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2752),
.B(n_2628),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2773),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2752),
.B(n_2693),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2774),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2733),
.B(n_2628),
.Y(n_3056)
);

OR2x2_ASAP7_75t_L g3057 ( 
.A(n_2977),
.B(n_2679),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2750),
.B(n_2628),
.Y(n_3058)
);

NOR2x1_ASAP7_75t_L g3059 ( 
.A(n_2809),
.B(n_2528),
.Y(n_3059)
);

INVx2_ASAP7_75t_SL g3060 ( 
.A(n_2910),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2893),
.B(n_2508),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2779),
.B(n_2508),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2783),
.Y(n_3063)
);

OAI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2786),
.A2(n_2676),
.B1(n_2438),
.B2(n_2671),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_2787),
.B(n_2544),
.Y(n_3065)
);

AOI21xp33_ASAP7_75t_L g3066 ( 
.A1(n_2831),
.A2(n_2648),
.B(n_2638),
.Y(n_3066)
);

OA21x2_ASAP7_75t_L g3067 ( 
.A1(n_2708),
.A2(n_2836),
.B(n_2844),
.Y(n_3067)
);

BUFx3_ASAP7_75t_L g3068 ( 
.A(n_2937),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2788),
.Y(n_3069)
);

INVx4_ASAP7_75t_L g3070 ( 
.A(n_2710),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2793),
.Y(n_3071)
);

INVxp67_ASAP7_75t_L g3072 ( 
.A(n_2770),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2978),
.B(n_2547),
.Y(n_3073)
);

OAI22xp5_ASAP7_75t_L g3074 ( 
.A1(n_2786),
.A2(n_2676),
.B1(n_2558),
.B2(n_2341),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2797),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_2777),
.B(n_2558),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2802),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2803),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2806),
.Y(n_3079)
);

OR2x2_ASAP7_75t_L g3080 ( 
.A(n_2777),
.B(n_2571),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_2800),
.B(n_2528),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2806),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_2800),
.B(n_2544),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2867),
.B(n_2463),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2807),
.B(n_2719),
.Y(n_3085)
);

AND2x2_ASAP7_75t_L g3086 ( 
.A(n_2937),
.B(n_2412),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2814),
.Y(n_3087)
);

INVx4_ASAP7_75t_L g3088 ( 
.A(n_2710),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2814),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2725),
.B(n_2571),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2824),
.Y(n_3091)
);

HB1xp67_ASAP7_75t_L g3092 ( 
.A(n_2905),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2824),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_2955),
.B(n_2489),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2756),
.Y(n_3095)
);

INVx3_ASAP7_75t_L g3096 ( 
.A(n_2769),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2756),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2826),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2826),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2765),
.Y(n_3100)
);

INVx4_ASAP7_75t_L g3101 ( 
.A(n_2710),
.Y(n_3101)
);

BUFx3_ASAP7_75t_L g3102 ( 
.A(n_2796),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2766),
.Y(n_3103)
);

BUFx3_ASAP7_75t_L g3104 ( 
.A(n_2796),
.Y(n_3104)
);

BUFx5_ASAP7_75t_L g3105 ( 
.A(n_2890),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2827),
.Y(n_3106)
);

AND2x4_ASAP7_75t_L g3107 ( 
.A(n_2820),
.B(n_2467),
.Y(n_3107)
);

INVxp67_ASAP7_75t_L g3108 ( 
.A(n_2689),
.Y(n_3108)
);

INVx6_ASAP7_75t_L g3109 ( 
.A(n_2915),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2832),
.B(n_2616),
.Y(n_3110)
);

HB1xp67_ASAP7_75t_L g3111 ( 
.A(n_2689),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2827),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_2808),
.B(n_2616),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2829),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2808),
.B(n_2600),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2829),
.Y(n_3116)
);

AND2x2_ASAP7_75t_L g3117 ( 
.A(n_2823),
.B(n_2775),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2823),
.B(n_2600),
.Y(n_3118)
);

INVx4_ASAP7_75t_L g3119 ( 
.A(n_2915),
.Y(n_3119)
);

AND2x2_ASAP7_75t_L g3120 ( 
.A(n_2775),
.B(n_2600),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2841),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_2776),
.B(n_2590),
.Y(n_3122)
);

HB1xp67_ASAP7_75t_L g3123 ( 
.A(n_2697),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2885),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_2776),
.B(n_2780),
.Y(n_3125)
);

BUFx2_ASAP7_75t_L g3126 ( 
.A(n_2759),
.Y(n_3126)
);

AND2x4_ASAP7_75t_L g3127 ( 
.A(n_2820),
.B(n_2344),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2841),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2842),
.Y(n_3129)
);

INVx3_ASAP7_75t_L g3130 ( 
.A(n_2782),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2780),
.B(n_2587),
.Y(n_3131)
);

BUFx2_ASAP7_75t_L g3132 ( 
.A(n_2763),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2842),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2707),
.B(n_2587),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2847),
.Y(n_3135)
);

HB1xp67_ASAP7_75t_L g3136 ( 
.A(n_2697),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2972),
.Y(n_3137)
);

INVx3_ASAP7_75t_L g3138 ( 
.A(n_2782),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2847),
.Y(n_3139)
);

BUFx2_ASAP7_75t_L g3140 ( 
.A(n_2843),
.Y(n_3140)
);

INVx3_ASAP7_75t_L g3141 ( 
.A(n_2782),
.Y(n_3141)
);

HB1xp67_ASAP7_75t_L g3142 ( 
.A(n_2919),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2849),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_2789),
.B(n_2590),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2849),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2707),
.B(n_2656),
.Y(n_3146)
);

OR2x2_ASAP7_75t_L g3147 ( 
.A(n_2789),
.B(n_2576),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2935),
.B(n_2656),
.Y(n_3148)
);

OR2x2_ASAP7_75t_L g3149 ( 
.A(n_2839),
.B(n_2860),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2860),
.B(n_2430),
.Y(n_3150)
);

BUFx2_ASAP7_75t_SL g3151 ( 
.A(n_2853),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2972),
.Y(n_3152)
);

OAI22xp5_ASAP7_75t_L g3153 ( 
.A1(n_2951),
.A2(n_2649),
.B1(n_2392),
.B2(n_2584),
.Y(n_3153)
);

AND2x2_ASAP7_75t_L g3154 ( 
.A(n_2703),
.B(n_2694),
.Y(n_3154)
);

AND2x2_ASAP7_75t_L g3155 ( 
.A(n_2703),
.B(n_2584),
.Y(n_3155)
);

INVx4_ASAP7_75t_L g3156 ( 
.A(n_2764),
.Y(n_3156)
);

OR2x2_ASAP7_75t_L g3157 ( 
.A(n_2865),
.B(n_2576),
.Y(n_3157)
);

BUFx2_ASAP7_75t_L g3158 ( 
.A(n_2821),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2865),
.B(n_2392),
.Y(n_3159)
);

OR2x2_ASAP7_75t_L g3160 ( 
.A(n_2876),
.B(n_2576),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2887),
.B(n_2683),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2891),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2891),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2892),
.Y(n_3164)
);

HB1xp67_ASAP7_75t_L g3165 ( 
.A(n_2942),
.Y(n_3165)
);

BUFx4f_ASAP7_75t_SL g3166 ( 
.A(n_2853),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_2898),
.B(n_2466),
.Y(n_3167)
);

INVx3_ASAP7_75t_L g3168 ( 
.A(n_2801),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2903),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2904),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2890),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2741),
.Y(n_3172)
);

HB1xp67_ASAP7_75t_L g3173 ( 
.A(n_2942),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_2911),
.B(n_2913),
.Y(n_3174)
);

INVx2_ASAP7_75t_SL g3175 ( 
.A(n_2821),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2741),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_2913),
.B(n_2925),
.Y(n_3177)
);

INVx6_ASAP7_75t_L g3178 ( 
.A(n_2927),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2928),
.Y(n_3179)
);

BUFx3_ASAP7_75t_L g3180 ( 
.A(n_2821),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_2772),
.B(n_2648),
.Y(n_3181)
);

AND2x2_ASAP7_75t_L g3182 ( 
.A(n_2790),
.B(n_2471),
.Y(n_3182)
);

HB1xp67_ASAP7_75t_L g3183 ( 
.A(n_2971),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2897),
.Y(n_3184)
);

INVxp67_ASAP7_75t_SL g3185 ( 
.A(n_2971),
.Y(n_3185)
);

NOR2x1_ASAP7_75t_L g3186 ( 
.A(n_2754),
.B(n_2668),
.Y(n_3186)
);

INVx3_ASAP7_75t_L g3187 ( 
.A(n_2801),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2833),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2840),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_2812),
.B(n_2662),
.Y(n_3190)
);

BUFx2_ASAP7_75t_L g3191 ( 
.A(n_2851),
.Y(n_3191)
);

HB1xp67_ASAP7_75t_L g3192 ( 
.A(n_2838),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2835),
.B(n_2593),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2686),
.Y(n_3194)
);

AND2x2_ASAP7_75t_L g3195 ( 
.A(n_2694),
.B(n_2482),
.Y(n_3195)
);

OR2x2_ASAP7_75t_L g3196 ( 
.A(n_2838),
.B(n_2639),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_2866),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2896),
.B(n_2366),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_2866),
.B(n_2482),
.Y(n_3199)
);

OAI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_2951),
.A2(n_2957),
.B1(n_2906),
.B2(n_2721),
.Y(n_3200)
);

BUFx3_ASAP7_75t_L g3201 ( 
.A(n_2851),
.Y(n_3201)
);

AOI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_2912),
.A2(n_2428),
.B1(n_2617),
.B2(n_2486),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2954),
.Y(n_3203)
);

AND2x4_ASAP7_75t_L g3204 ( 
.A(n_2820),
.B(n_2660),
.Y(n_3204)
);

AND2x2_ASAP7_75t_L g3205 ( 
.A(n_3048),
.B(n_2888),
.Y(n_3205)
);

OR2x2_ASAP7_75t_L g3206 ( 
.A(n_3027),
.B(n_2696),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3058),
.B(n_2848),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2982),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_3154),
.B(n_2852),
.Y(n_3209)
);

OR2x2_ASAP7_75t_L g3210 ( 
.A(n_3192),
.B(n_2888),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_3174),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_3177),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2985),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2989),
.Y(n_3214)
);

INVx3_ASAP7_75t_L g3215 ( 
.A(n_3156),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2990),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_2996),
.B(n_2952),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_3054),
.B(n_2921),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3007),
.B(n_2926),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2999),
.Y(n_3220)
);

AND2x2_ASAP7_75t_L g3221 ( 
.A(n_3068),
.B(n_2950),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3001),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3002),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_3125),
.Y(n_3224)
);

AND2x2_ASAP7_75t_L g3225 ( 
.A(n_3068),
.B(n_2922),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_2998),
.B(n_2922),
.Y(n_3226)
);

AND2x6_ASAP7_75t_SL g3227 ( 
.A(n_3003),
.B(n_3000),
.Y(n_3227)
);

AND2x4_ASAP7_75t_SL g3228 ( 
.A(n_3119),
.B(n_2927),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_3200),
.A2(n_2916),
.B1(n_2973),
.B2(n_2957),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3006),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3117),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3018),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3154),
.B(n_2855),
.Y(n_3233)
);

AND2x2_ASAP7_75t_L g3234 ( 
.A(n_3005),
.B(n_2815),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_3194),
.B(n_2856),
.Y(n_3235)
);

INVx3_ASAP7_75t_L g3236 ( 
.A(n_3156),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_3158),
.B(n_2816),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3148),
.B(n_2687),
.Y(n_3238)
);

AND2x4_ASAP7_75t_L g3239 ( 
.A(n_3070),
.B(n_3088),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3022),
.Y(n_3240)
);

AND2x2_ASAP7_75t_L g3241 ( 
.A(n_3191),
.B(n_2817),
.Y(n_3241)
);

INVx3_ASAP7_75t_L g3242 ( 
.A(n_3156),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_3113),
.B(n_2875),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3015),
.B(n_2878),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3025),
.Y(n_3245)
);

AND2x4_ASAP7_75t_SL g3246 ( 
.A(n_3119),
.B(n_2691),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3031),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_3188),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_3175),
.B(n_2825),
.Y(n_3249)
);

AND2x4_ASAP7_75t_L g3250 ( 
.A(n_3070),
.B(n_2944),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_3166),
.B(n_2799),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3095),
.Y(n_3252)
);

NAND4xp25_ASAP7_75t_L g3253 ( 
.A(n_3000),
.B(n_2721),
.C(n_2906),
.D(n_2873),
.Y(n_3253)
);

AND2x4_ASAP7_75t_L g3254 ( 
.A(n_3070),
.B(n_2944),
.Y(n_3254)
);

BUFx4f_ASAP7_75t_SL g3255 ( 
.A(n_2983),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_3095),
.Y(n_3256)
);

AND2x4_ASAP7_75t_L g3257 ( 
.A(n_3088),
.B(n_2944),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3090),
.B(n_2879),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3056),
.B(n_2880),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3175),
.B(n_3024),
.Y(n_3260)
);

BUFx2_ASAP7_75t_L g3261 ( 
.A(n_3119),
.Y(n_3261)
);

OR2x2_ASAP7_75t_L g3262 ( 
.A(n_3192),
.B(n_2810),
.Y(n_3262)
);

OR2x2_ASAP7_75t_L g3263 ( 
.A(n_3008),
.B(n_2947),
.Y(n_3263)
);

OAI21xp33_ASAP7_75t_L g3264 ( 
.A1(n_3066),
.A2(n_2973),
.B(n_2946),
.Y(n_3264)
);

AND2x2_ASAP7_75t_L g3265 ( 
.A(n_3026),
.B(n_2851),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3189),
.Y(n_3266)
);

AND2x2_ASAP7_75t_L g3267 ( 
.A(n_3180),
.B(n_2947),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_3180),
.B(n_2947),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_3201),
.B(n_2837),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_3097),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_3122),
.B(n_2881),
.Y(n_3271)
);

AND2x2_ASAP7_75t_L g3272 ( 
.A(n_3201),
.B(n_2837),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3009),
.B(n_3035),
.Y(n_3273)
);

INVx2_ASAP7_75t_L g3274 ( 
.A(n_3097),
.Y(n_3274)
);

AOI22xp33_ASAP7_75t_L g3275 ( 
.A1(n_3021),
.A2(n_2920),
.B1(n_2714),
.B2(n_2886),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3036),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_3100),
.Y(n_3277)
);

AND2x2_ASAP7_75t_L g3278 ( 
.A(n_3012),
.B(n_3184),
.Y(n_3278)
);

AND2x2_ASAP7_75t_L g3279 ( 
.A(n_3013),
.B(n_2688),
.Y(n_3279)
);

INVx3_ASAP7_75t_L g3280 ( 
.A(n_3038),
.Y(n_3280)
);

HB1xp67_ASAP7_75t_L g3281 ( 
.A(n_3008),
.Y(n_3281)
);

INVxp67_ASAP7_75t_SL g3282 ( 
.A(n_3020),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3039),
.Y(n_3283)
);

AND2x4_ASAP7_75t_SL g3284 ( 
.A(n_3038),
.B(n_2698),
.Y(n_3284)
);

INVx1_ASAP7_75t_SL g3285 ( 
.A(n_3102),
.Y(n_3285)
);

AND2x2_ASAP7_75t_L g3286 ( 
.A(n_2995),
.B(n_2688),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3131),
.B(n_2914),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3041),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3100),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3144),
.B(n_2918),
.Y(n_3290)
);

BUFx2_ASAP7_75t_SL g3291 ( 
.A(n_2983),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3051),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_2993),
.B(n_2695),
.Y(n_3293)
);

AND2x4_ASAP7_75t_L g3294 ( 
.A(n_3088),
.B(n_3101),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3053),
.Y(n_3295)
);

AOI22xp33_ASAP7_75t_L g3296 ( 
.A1(n_3146),
.A2(n_2755),
.B1(n_2748),
.B2(n_2753),
.Y(n_3296)
);

OR2x2_ASAP7_75t_L g3297 ( 
.A(n_3020),
.B(n_3030),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3055),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3149),
.B(n_2974),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_2991),
.B(n_2695),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3030),
.B(n_2699),
.Y(n_3301)
);

AND2x2_ASAP7_75t_L g3302 ( 
.A(n_3092),
.B(n_2699),
.Y(n_3302)
);

AND2x4_ASAP7_75t_L g3303 ( 
.A(n_3101),
.B(n_2804),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3103),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3092),
.B(n_2705),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3063),
.Y(n_3306)
);

NAND2x1_ASAP7_75t_L g3307 ( 
.A(n_3101),
.B(n_2764),
.Y(n_3307)
);

BUFx2_ASAP7_75t_L g3308 ( 
.A(n_3102),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3069),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3197),
.B(n_3042),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3016),
.B(n_2705),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3046),
.B(n_2979),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3071),
.Y(n_3313)
);

AND2x4_ASAP7_75t_L g3314 ( 
.A(n_3186),
.B(n_2794),
.Y(n_3314)
);

NOR2x1_ASAP7_75t_L g3315 ( 
.A(n_3038),
.B(n_2754),
.Y(n_3315)
);

OR2x2_ASAP7_75t_L g3316 ( 
.A(n_3080),
.B(n_2740),
.Y(n_3316)
);

INVxp67_ASAP7_75t_L g3317 ( 
.A(n_3111),
.Y(n_3317)
);

AND2x2_ASAP7_75t_L g3318 ( 
.A(n_2986),
.B(n_3032),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3075),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3047),
.B(n_2980),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3077),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3044),
.B(n_2981),
.Y(n_3322)
);

OR2x2_ASAP7_75t_L g3323 ( 
.A(n_3057),
.B(n_2742),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_2986),
.B(n_2747),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3078),
.Y(n_3325)
);

OR2x2_ASAP7_75t_L g3326 ( 
.A(n_3010),
.B(n_2743),
.Y(n_3326)
);

NOR2xp67_ASAP7_75t_L g3327 ( 
.A(n_3060),
.B(n_2724),
.Y(n_3327)
);

INVxp67_ASAP7_75t_SL g3328 ( 
.A(n_3124),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3110),
.B(n_2834),
.Y(n_3329)
);

BUFx3_ASAP7_75t_L g3330 ( 
.A(n_3014),
.Y(n_3330)
);

OR2x2_ASAP7_75t_L g3331 ( 
.A(n_3010),
.B(n_2744),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3111),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3034),
.B(n_2822),
.Y(n_3333)
);

AND2x2_ASAP7_75t_L g3334 ( 
.A(n_3104),
.B(n_2834),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_3104),
.B(n_2845),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_3171),
.B(n_2845),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3123),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_3123),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3134),
.B(n_2822),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3136),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3073),
.B(n_2931),
.Y(n_3341)
);

OR2x2_ASAP7_75t_L g3342 ( 
.A(n_3019),
.B(n_2751),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_3045),
.B(n_2976),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3136),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3171),
.B(n_2862),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3079),
.Y(n_3346)
);

INVx3_ASAP7_75t_SL g3347 ( 
.A(n_3003),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3082),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_3087),
.Y(n_3349)
);

OR2x2_ASAP7_75t_L g3350 ( 
.A(n_3019),
.B(n_3033),
.Y(n_3350)
);

AND2x2_ASAP7_75t_L g3351 ( 
.A(n_3028),
.B(n_2862),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3089),
.Y(n_3352)
);

INVx1_ASAP7_75t_SL g3353 ( 
.A(n_3109),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3091),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3093),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3098),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_3073),
.B(n_2931),
.Y(n_3357)
);

AND2x4_ASAP7_75t_L g3358 ( 
.A(n_2992),
.B(n_2795),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3099),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3052),
.B(n_2864),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3181),
.B(n_2949),
.Y(n_3361)
);

BUFx3_ASAP7_75t_L g3362 ( 
.A(n_3166),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3106),
.Y(n_3363)
);

NOR2xp33_ASAP7_75t_L g3364 ( 
.A(n_2994),
.B(n_2716),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3115),
.B(n_2949),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3112),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3114),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3126),
.B(n_2864),
.Y(n_3368)
);

BUFx2_ASAP7_75t_L g3369 ( 
.A(n_3017),
.Y(n_3369)
);

OR2x2_ASAP7_75t_L g3370 ( 
.A(n_3033),
.B(n_2757),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3116),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3121),
.Y(n_3372)
);

NOR2xp33_ASAP7_75t_L g3373 ( 
.A(n_3037),
.B(n_2758),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3132),
.B(n_2954),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3118),
.B(n_2889),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3128),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3140),
.B(n_2929),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3129),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_2992),
.B(n_2929),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_3133),
.B(n_2894),
.Y(n_3380)
);

INVx2_ASAP7_75t_L g3381 ( 
.A(n_3135),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3208),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_3218),
.B(n_2997),
.Y(n_3383)
);

NAND2x1_ASAP7_75t_SL g3384 ( 
.A(n_3347),
.B(n_3059),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3213),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_3252),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3273),
.B(n_3108),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_3278),
.B(n_3108),
.Y(n_3388)
);

INVxp67_ASAP7_75t_SL g3389 ( 
.A(n_3328),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3318),
.B(n_3072),
.Y(n_3390)
);

AND2x4_ASAP7_75t_L g3391 ( 
.A(n_3250),
.B(n_3107),
.Y(n_3391)
);

AND2x2_ASAP7_75t_L g3392 ( 
.A(n_3209),
.B(n_3155),
.Y(n_3392)
);

AND2x2_ASAP7_75t_L g3393 ( 
.A(n_3209),
.B(n_3155),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3214),
.Y(n_3394)
);

BUFx2_ASAP7_75t_L g3395 ( 
.A(n_3261),
.Y(n_3395)
);

OR2x2_ASAP7_75t_L g3396 ( 
.A(n_3231),
.B(n_3072),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3260),
.B(n_2997),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3205),
.B(n_2997),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3233),
.B(n_3195),
.Y(n_3399)
);

OR2x2_ASAP7_75t_L g3400 ( 
.A(n_3310),
.B(n_3040),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3216),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3220),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3222),
.Y(n_3403)
);

HB1xp67_ASAP7_75t_L g3404 ( 
.A(n_3281),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3233),
.B(n_3195),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3256),
.Y(n_3406)
);

CKINVDCx5p33_ASAP7_75t_R g3407 ( 
.A(n_3291),
.Y(n_3407)
);

AND2x2_ASAP7_75t_L g3408 ( 
.A(n_3219),
.B(n_3076),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3265),
.B(n_3029),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3223),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_3234),
.B(n_3076),
.Y(n_3411)
);

AND2x2_ASAP7_75t_L g3412 ( 
.A(n_3351),
.B(n_3029),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3275),
.B(n_3373),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_3253),
.B(n_3085),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3275),
.B(n_3139),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3373),
.B(n_3143),
.Y(n_3416)
);

AND2x4_ASAP7_75t_L g3417 ( 
.A(n_3250),
.B(n_3107),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3230),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3279),
.B(n_3226),
.Y(n_3419)
);

AND2x4_ASAP7_75t_L g3420 ( 
.A(n_3254),
.B(n_3107),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3270),
.Y(n_3421)
);

OR2x2_ASAP7_75t_L g3422 ( 
.A(n_3310),
.B(n_3137),
.Y(n_3422)
);

OR2x2_ASAP7_75t_L g3423 ( 
.A(n_3211),
.B(n_3137),
.Y(n_3423)
);

BUFx2_ASAP7_75t_L g3424 ( 
.A(n_3308),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3232),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3217),
.B(n_3145),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3240),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3324),
.B(n_3029),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3243),
.B(n_3162),
.Y(n_3429)
);

INVx3_ASAP7_75t_L g3430 ( 
.A(n_3215),
.Y(n_3430)
);

AND2x2_ASAP7_75t_L g3431 ( 
.A(n_3341),
.B(n_3067),
.Y(n_3431)
);

OR2x2_ASAP7_75t_L g3432 ( 
.A(n_3212),
.B(n_3152),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_3274),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_SL g3434 ( 
.A(n_3255),
.B(n_2784),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3245),
.Y(n_3435)
);

OR2x2_ASAP7_75t_L g3436 ( 
.A(n_3297),
.B(n_3152),
.Y(n_3436)
);

BUFx2_ASAP7_75t_L g3437 ( 
.A(n_3215),
.Y(n_3437)
);

AND2x2_ASAP7_75t_L g3438 ( 
.A(n_3293),
.B(n_3061),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3247),
.Y(n_3439)
);

INVxp67_ASAP7_75t_L g3440 ( 
.A(n_3281),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3248),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3300),
.B(n_2987),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3286),
.B(n_2987),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3266),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3243),
.B(n_3163),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3277),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3289),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3244),
.B(n_3164),
.Y(n_3448)
);

INVx1_ASAP7_75t_SL g3449 ( 
.A(n_3246),
.Y(n_3449)
);

AND2x2_ASAP7_75t_L g3450 ( 
.A(n_3311),
.B(n_3193),
.Y(n_3450)
);

OR2x2_ASAP7_75t_L g3451 ( 
.A(n_3224),
.B(n_3142),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_3360),
.B(n_3190),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_3304),
.Y(n_3453)
);

NOR2x1_ASAP7_75t_L g3454 ( 
.A(n_3315),
.B(n_3017),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3276),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3283),
.Y(n_3456)
);

AND2x4_ASAP7_75t_L g3457 ( 
.A(n_3254),
.B(n_3043),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3244),
.B(n_3169),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3323),
.B(n_3170),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_3341),
.B(n_3067),
.Y(n_3460)
);

AND2x2_ASAP7_75t_L g3461 ( 
.A(n_3357),
.B(n_3067),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3288),
.Y(n_3462)
);

AND2x4_ASAP7_75t_L g3463 ( 
.A(n_3257),
.B(n_3043),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3292),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3271),
.B(n_3179),
.Y(n_3465)
);

AND2x2_ASAP7_75t_L g3466 ( 
.A(n_3357),
.B(n_2988),
.Y(n_3466)
);

HB1xp67_ASAP7_75t_L g3467 ( 
.A(n_3282),
.Y(n_3467)
);

INVx2_ASAP7_75t_SL g3468 ( 
.A(n_3236),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3225),
.B(n_3120),
.Y(n_3469)
);

OR2x2_ASAP7_75t_L g3470 ( 
.A(n_3350),
.B(n_3142),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3295),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_3419),
.B(n_3408),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_3467),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3408),
.B(n_3379),
.Y(n_3474)
);

AOI32xp33_ASAP7_75t_L g3475 ( 
.A1(n_3449),
.A2(n_3228),
.A3(n_3284),
.B1(n_3264),
.B2(n_3330),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3382),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3385),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3394),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3467),
.Y(n_3479)
);

NAND2x1p5_ASAP7_75t_L g3480 ( 
.A(n_3454),
.B(n_3236),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3401),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3402),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3403),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3431),
.B(n_3339),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3410),
.Y(n_3485)
);

AND2x2_ASAP7_75t_L g3486 ( 
.A(n_3438),
.B(n_3269),
.Y(n_3486)
);

AND2x2_ASAP7_75t_L g3487 ( 
.A(n_3443),
.B(n_3272),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3418),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3395),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3425),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3431),
.B(n_3339),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3427),
.Y(n_3492)
);

OR2x2_ASAP7_75t_L g3493 ( 
.A(n_3400),
.B(n_3375),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3435),
.Y(n_3494)
);

NAND2x2_ASAP7_75t_L g3495 ( 
.A(n_3413),
.B(n_3362),
.Y(n_3495)
);

AND2x4_ASAP7_75t_L g3496 ( 
.A(n_3457),
.B(n_3285),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3411),
.B(n_3206),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3439),
.Y(n_3498)
);

OR2x2_ASAP7_75t_L g3499 ( 
.A(n_3387),
.B(n_3426),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3441),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3411),
.B(n_3392),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3444),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3460),
.B(n_3333),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3455),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3460),
.B(n_3333),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3456),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3392),
.B(n_3329),
.Y(n_3507)
);

NAND2xp33_ASAP7_75t_SL g3508 ( 
.A(n_3384),
.B(n_3242),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3462),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3464),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3471),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3422),
.Y(n_3512)
);

OR2x2_ASAP7_75t_L g3513 ( 
.A(n_3388),
.B(n_3375),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_L g3514 ( 
.A(n_3414),
.B(n_3253),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3461),
.B(n_3332),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3396),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3389),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3404),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_3407),
.B(n_3178),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3461),
.B(n_3337),
.Y(n_3520)
);

NOR2xp67_ASAP7_75t_SL g3521 ( 
.A(n_3407),
.B(n_3178),
.Y(n_3521)
);

INVx2_ASAP7_75t_SL g3522 ( 
.A(n_3424),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3404),
.Y(n_3523)
);

AOI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3414),
.A2(n_3229),
.B1(n_3264),
.B2(n_3074),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3470),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3465),
.Y(n_3526)
);

INVx2_ASAP7_75t_SL g3527 ( 
.A(n_3437),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3393),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3389),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3451),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3393),
.Y(n_3531)
);

NOR2xp67_ASAP7_75t_L g3532 ( 
.A(n_3430),
.B(n_3242),
.Y(n_3532)
);

AND2x2_ASAP7_75t_L g3533 ( 
.A(n_3450),
.B(n_3301),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3448),
.Y(n_3534)
);

OR2x2_ASAP7_75t_L g3535 ( 
.A(n_3390),
.B(n_3365),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3399),
.B(n_3338),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3458),
.Y(n_3537)
);

OR2x2_ASAP7_75t_L g3538 ( 
.A(n_3399),
.B(n_3365),
.Y(n_3538)
);

NOR2x1_ASAP7_75t_L g3539 ( 
.A(n_3430),
.B(n_3327),
.Y(n_3539)
);

OR2x2_ASAP7_75t_L g3540 ( 
.A(n_3405),
.B(n_3259),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3484),
.B(n_3405),
.Y(n_3541)
);

NOR2xp33_ASAP7_75t_L g3542 ( 
.A(n_3514),
.B(n_3434),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3484),
.B(n_3440),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3515),
.Y(n_3544)
);

INVx1_ASAP7_75t_SL g3545 ( 
.A(n_3496),
.Y(n_3545)
);

OR2x2_ASAP7_75t_L g3546 ( 
.A(n_3538),
.B(n_3491),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3515),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3517),
.Y(n_3548)
);

INVx1_ASAP7_75t_SL g3549 ( 
.A(n_3522),
.Y(n_3549)
);

AND2x2_ASAP7_75t_SL g3550 ( 
.A(n_3496),
.B(n_3519),
.Y(n_3550)
);

OAI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3514),
.A2(n_3229),
.B(n_3364),
.Y(n_3551)
);

OAI21xp33_ASAP7_75t_L g3552 ( 
.A1(n_3524),
.A2(n_3415),
.B(n_3251),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3486),
.B(n_3469),
.Y(n_3553)
);

OAI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_3524),
.A2(n_3468),
.B(n_3285),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_3501),
.B(n_3442),
.Y(n_3555)
);

INVx2_ASAP7_75t_SL g3556 ( 
.A(n_3527),
.Y(n_3556)
);

OAI22xp5_ASAP7_75t_L g3557 ( 
.A1(n_3495),
.A2(n_3255),
.B1(n_3468),
.B2(n_3430),
.Y(n_3557)
);

AO21x1_ASAP7_75t_L g3558 ( 
.A1(n_3508),
.A2(n_3343),
.B(n_3282),
.Y(n_3558)
);

AND2x4_ASAP7_75t_L g3559 ( 
.A(n_3532),
.B(n_3539),
.Y(n_3559)
);

INVxp67_ASAP7_75t_L g3560 ( 
.A(n_3489),
.Y(n_3560)
);

OAI21xp33_ASAP7_75t_L g3561 ( 
.A1(n_3475),
.A2(n_3416),
.B(n_3296),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3520),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3520),
.Y(n_3563)
);

OAI22xp33_ASAP7_75t_L g3564 ( 
.A1(n_3532),
.A2(n_3369),
.B1(n_3280),
.B2(n_3353),
.Y(n_3564)
);

O2A1O1Ixp33_ASAP7_75t_L g3565 ( 
.A1(n_3518),
.A2(n_2877),
.B(n_2884),
.C(n_2819),
.Y(n_3565)
);

AOI21x1_ASAP7_75t_L g3566 ( 
.A1(n_3521),
.A2(n_3529),
.B(n_3307),
.Y(n_3566)
);

OR2x2_ASAP7_75t_L g3567 ( 
.A(n_3491),
.B(n_3436),
.Y(n_3567)
);

OAI21xp33_ASAP7_75t_L g3568 ( 
.A1(n_3503),
.A2(n_3296),
.B(n_3429),
.Y(n_3568)
);

NAND2x1_ASAP7_75t_L g3569 ( 
.A(n_3472),
.B(n_3280),
.Y(n_3569)
);

OAI32xp33_ASAP7_75t_L g3570 ( 
.A1(n_3480),
.A2(n_3353),
.A3(n_3263),
.B1(n_3440),
.B2(n_3428),
.Y(n_3570)
);

OAI21xp5_ASAP7_75t_SL g3571 ( 
.A1(n_3480),
.A2(n_3303),
.B(n_2729),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3476),
.Y(n_3572)
);

AOI21xp33_ASAP7_75t_L g3573 ( 
.A1(n_3523),
.A2(n_3331),
.B(n_3326),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3497),
.B(n_3383),
.Y(n_3574)
);

OR2x2_ASAP7_75t_L g3575 ( 
.A(n_3503),
.B(n_3423),
.Y(n_3575)
);

HB1xp67_ASAP7_75t_L g3576 ( 
.A(n_3473),
.Y(n_3576)
);

OR2x2_ASAP7_75t_L g3577 ( 
.A(n_3505),
.B(n_3432),
.Y(n_3577)
);

INVx1_ASAP7_75t_SL g3578 ( 
.A(n_3533),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3505),
.B(n_3466),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3477),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_3474),
.B(n_3466),
.Y(n_3581)
);

OR2x2_ASAP7_75t_L g3582 ( 
.A(n_3535),
.B(n_3493),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3479),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3478),
.Y(n_3584)
);

INVx2_ASAP7_75t_SL g3585 ( 
.A(n_3487),
.Y(n_3585)
);

AND2x2_ASAP7_75t_L g3586 ( 
.A(n_3507),
.B(n_3452),
.Y(n_3586)
);

OAI322xp33_ASAP7_75t_L g3587 ( 
.A1(n_3526),
.A2(n_3316),
.A3(n_3459),
.B1(n_3445),
.B2(n_3238),
.C1(n_3370),
.C2(n_3342),
.Y(n_3587)
);

AOI21xp5_ASAP7_75t_SL g3588 ( 
.A1(n_3481),
.A2(n_3303),
.B(n_3257),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3482),
.Y(n_3589)
);

NAND3xp33_ASAP7_75t_SL g3590 ( 
.A(n_3540),
.B(n_2749),
.C(n_2672),
.Y(n_3590)
);

HB1xp67_ASAP7_75t_L g3591 ( 
.A(n_3530),
.Y(n_3591)
);

OAI221xp5_ASAP7_75t_L g3592 ( 
.A1(n_3534),
.A2(n_3537),
.B1(n_3151),
.B2(n_3525),
.C(n_3488),
.Y(n_3592)
);

OR2x2_ASAP7_75t_L g3593 ( 
.A(n_3513),
.B(n_3259),
.Y(n_3593)
);

A2O1A1Ixp33_ASAP7_75t_L g3594 ( 
.A1(n_3499),
.A2(n_3060),
.B(n_2729),
.C(n_3374),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3483),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3528),
.B(n_3398),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3485),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3490),
.Y(n_3598)
);

INVx1_ASAP7_75t_SL g3599 ( 
.A(n_3516),
.Y(n_3599)
);

OAI22xp33_ASAP7_75t_L g3600 ( 
.A1(n_3531),
.A2(n_3536),
.B1(n_3178),
.B2(n_3317),
.Y(n_3600)
);

INVx2_ASAP7_75t_SL g3601 ( 
.A(n_3512),
.Y(n_3601)
);

AOI321xp33_ASAP7_75t_L g3602 ( 
.A1(n_3552),
.A2(n_3542),
.A3(n_3561),
.B1(n_3570),
.B2(n_3592),
.C(n_3565),
.Y(n_3602)
);

OR2x2_ASAP7_75t_L g3603 ( 
.A(n_3546),
.B(n_3536),
.Y(n_3603)
);

O2A1O1Ixp33_ASAP7_75t_L g3604 ( 
.A1(n_3551),
.A2(n_2819),
.B(n_3023),
.C(n_3064),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3567),
.Y(n_3605)
);

OAI21xp5_ASAP7_75t_SL g3606 ( 
.A1(n_3571),
.A2(n_2720),
.B(n_3227),
.Y(n_3606)
);

OR2x2_ASAP7_75t_L g3607 ( 
.A(n_3582),
.B(n_3492),
.Y(n_3607)
);

OAI22xp5_ASAP7_75t_L g3608 ( 
.A1(n_3550),
.A2(n_2781),
.B1(n_3397),
.B2(n_3391),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3568),
.B(n_3552),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3575),
.Y(n_3610)
);

OAI322xp33_ASAP7_75t_SL g3611 ( 
.A1(n_3541),
.A2(n_3511),
.A3(n_3510),
.B1(n_3494),
.B2(n_3498),
.C1(n_3500),
.C2(n_3502),
.Y(n_3611)
);

AOI222xp33_ASAP7_75t_L g3612 ( 
.A1(n_3590),
.A2(n_3509),
.B1(n_3506),
.B2(n_3504),
.C1(n_3309),
.C2(n_3298),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3577),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3588),
.A2(n_3317),
.B(n_3457),
.Y(n_3614)
);

AOI22xp33_ASAP7_75t_SL g3615 ( 
.A1(n_3554),
.A2(n_3391),
.B1(n_3420),
.B2(n_3417),
.Y(n_3615)
);

AOI22xp5_ASAP7_75t_L g3616 ( 
.A1(n_3561),
.A2(n_3412),
.B1(n_3409),
.B2(n_3391),
.Y(n_3616)
);

AND2x2_ASAP7_75t_L g3617 ( 
.A(n_3545),
.B(n_3457),
.Y(n_3617)
);

HB1xp67_ASAP7_75t_L g3618 ( 
.A(n_3591),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3545),
.B(n_3463),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3569),
.B(n_3463),
.Y(n_3620)
);

AOI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_3568),
.A2(n_3420),
.B1(n_3417),
.B2(n_3377),
.Y(n_3621)
);

AOI21xp33_ASAP7_75t_L g3622 ( 
.A1(n_3549),
.A2(n_2870),
.B(n_3262),
.Y(n_3622)
);

OAI22xp33_ASAP7_75t_L g3623 ( 
.A1(n_3571),
.A2(n_3196),
.B1(n_3109),
.B2(n_3238),
.Y(n_3623)
);

NAND3xp33_ASAP7_75t_SL g3624 ( 
.A(n_3558),
.B(n_2749),
.C(n_2943),
.Y(n_3624)
);

OAI22xp5_ASAP7_75t_L g3625 ( 
.A1(n_3594),
.A2(n_2781),
.B1(n_3420),
.B2(n_3417),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3544),
.B(n_3340),
.Y(n_3626)
);

INVx1_ASAP7_75t_SL g3627 ( 
.A(n_3556),
.Y(n_3627)
);

OAI332xp33_ASAP7_75t_L g3628 ( 
.A1(n_3599),
.A2(n_3153),
.A3(n_2901),
.B1(n_3313),
.B2(n_3306),
.B3(n_3325),
.C1(n_3319),
.C2(n_3321),
.Y(n_3628)
);

AND2x4_ASAP7_75t_L g3629 ( 
.A(n_3559),
.B(n_3463),
.Y(n_3629)
);

AOI22xp33_ASAP7_75t_L g3630 ( 
.A1(n_3587),
.A2(n_3086),
.B1(n_3268),
.B2(n_3267),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3589),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3543),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3547),
.B(n_3344),
.Y(n_3633)
);

AOI211x1_ASAP7_75t_L g3634 ( 
.A1(n_3600),
.A2(n_3227),
.B(n_3221),
.C(n_3368),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_3581),
.B(n_3302),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3562),
.B(n_3312),
.Y(n_3636)
);

OAI22xp5_ASAP7_75t_L g3637 ( 
.A1(n_3578),
.A2(n_3294),
.B1(n_3239),
.B2(n_3109),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3586),
.B(n_3305),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3563),
.Y(n_3639)
);

OAI21xp33_ASAP7_75t_L g3640 ( 
.A1(n_3601),
.A2(n_3361),
.B(n_3320),
.Y(n_3640)
);

NOR2xp67_ASAP7_75t_L g3641 ( 
.A(n_3559),
.B(n_2830),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3579),
.B(n_3312),
.Y(n_3642)
);

OAI221xp5_ASAP7_75t_L g3643 ( 
.A1(n_3602),
.A2(n_3557),
.B1(n_3560),
.B2(n_3573),
.C(n_3566),
.Y(n_3643)
);

AOI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_3609),
.A2(n_3624),
.B1(n_3625),
.B2(n_3616),
.Y(n_3644)
);

O2A1O1Ixp33_ASAP7_75t_L g3645 ( 
.A1(n_3627),
.A2(n_3587),
.B(n_3564),
.C(n_3580),
.Y(n_3645)
);

NAND4xp25_ASAP7_75t_L g3646 ( 
.A(n_3634),
.B(n_3604),
.C(n_3606),
.D(n_3615),
.Y(n_3646)
);

NAND3xp33_ASAP7_75t_L g3647 ( 
.A(n_3612),
.B(n_3584),
.C(n_3572),
.Y(n_3647)
);

AOI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_3606),
.A2(n_3585),
.B(n_3576),
.Y(n_3648)
);

NOR2xp33_ASAP7_75t_L g3649 ( 
.A(n_3632),
.B(n_2907),
.Y(n_3649)
);

NOR2xp33_ASAP7_75t_SL g3650 ( 
.A(n_3641),
.B(n_2784),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3618),
.Y(n_3651)
);

OAI221xp5_ASAP7_75t_L g3652 ( 
.A1(n_3621),
.A2(n_3598),
.B1(n_3597),
.B2(n_3595),
.C(n_3593),
.Y(n_3652)
);

AOI221xp5_ASAP7_75t_L g3653 ( 
.A1(n_3611),
.A2(n_3596),
.B1(n_3548),
.B2(n_3583),
.C(n_3553),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3639),
.B(n_3555),
.Y(n_3654)
);

OAI222xp33_ASAP7_75t_L g3655 ( 
.A1(n_3608),
.A2(n_3574),
.B1(n_3271),
.B2(n_3258),
.C1(n_3207),
.C2(n_3320),
.Y(n_3655)
);

AOI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3623),
.A2(n_3237),
.B1(n_3241),
.B2(n_3084),
.Y(n_3656)
);

NOR4xp25_ASAP7_75t_L g3657 ( 
.A(n_3628),
.B(n_2746),
.C(n_2745),
.D(n_3011),
.Y(n_3657)
);

OAI21xp33_ASAP7_75t_SL g3658 ( 
.A1(n_3620),
.A2(n_3335),
.B(n_3334),
.Y(n_3658)
);

AOI222xp33_ASAP7_75t_L g3659 ( 
.A1(n_3640),
.A2(n_3258),
.B1(n_3207),
.B2(n_3235),
.C1(n_3094),
.C2(n_3361),
.Y(n_3659)
);

AOI222xp33_ASAP7_75t_L g3660 ( 
.A1(n_3630),
.A2(n_3235),
.B1(n_3290),
.B2(n_3287),
.C1(n_3249),
.C2(n_3299),
.Y(n_3660)
);

NAND3xp33_ASAP7_75t_L g3661 ( 
.A(n_3637),
.B(n_3182),
.C(n_3202),
.Y(n_3661)
);

NOR3xp33_ASAP7_75t_SL g3662 ( 
.A(n_3614),
.B(n_2943),
.C(n_3198),
.Y(n_3662)
);

NOR3xp33_ASAP7_75t_L g3663 ( 
.A(n_3628),
.B(n_2830),
.C(n_2850),
.Y(n_3663)
);

AOI221x1_ASAP7_75t_L g3664 ( 
.A1(n_3622),
.A2(n_3629),
.B1(n_3605),
.B2(n_3610),
.C(n_3613),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3607),
.Y(n_3665)
);

INVxp67_ASAP7_75t_L g3666 ( 
.A(n_3626),
.Y(n_3666)
);

NOR3xp33_ASAP7_75t_L g3667 ( 
.A(n_3633),
.B(n_2858),
.C(n_2857),
.Y(n_3667)
);

NOR2xp33_ASAP7_75t_L g3668 ( 
.A(n_3603),
.B(n_3642),
.Y(n_3668)
);

NOR2x1_ASAP7_75t_L g3669 ( 
.A(n_3629),
.B(n_3611),
.Y(n_3669)
);

INVx2_ASAP7_75t_SL g3670 ( 
.A(n_3617),
.Y(n_3670)
);

AOI22xp33_ASAP7_75t_L g3671 ( 
.A1(n_3619),
.A2(n_3294),
.B1(n_3239),
.B2(n_3336),
.Y(n_3671)
);

AOI211xp5_ASAP7_75t_L g3672 ( 
.A1(n_3636),
.A2(n_3345),
.B(n_2720),
.C(n_3050),
.Y(n_3672)
);

OAI311xp33_ASAP7_75t_L g3673 ( 
.A1(n_3631),
.A2(n_3202),
.A3(n_3210),
.B1(n_3287),
.C1(n_3290),
.Y(n_3673)
);

AOI321xp33_ASAP7_75t_L g3674 ( 
.A1(n_3638),
.A2(n_3049),
.A3(n_2988),
.B1(n_3299),
.B2(n_3043),
.C(n_3322),
.Y(n_3674)
);

NAND4xp25_ASAP7_75t_SL g3675 ( 
.A(n_3635),
.B(n_2861),
.C(n_2871),
.D(n_2859),
.Y(n_3675)
);

NOR3xp33_ASAP7_75t_L g3676 ( 
.A(n_3624),
.B(n_2874),
.C(n_3203),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3624),
.A2(n_2961),
.B(n_2791),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3618),
.Y(n_3678)
);

NOR2xp33_ASAP7_75t_L g3679 ( 
.A(n_3627),
.B(n_2895),
.Y(n_3679)
);

OAI21xp33_ASAP7_75t_SL g3680 ( 
.A1(n_3641),
.A2(n_3328),
.B(n_3185),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_3624),
.A2(n_3322),
.B(n_3004),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_SL g3682 ( 
.A(n_3641),
.B(n_3314),
.Y(n_3682)
);

AND5x1_ASAP7_75t_L g3683 ( 
.A(n_3602),
.B(n_2603),
.C(n_2520),
.D(n_2895),
.E(n_2678),
.Y(n_3683)
);

NAND4xp25_ASAP7_75t_L g3684 ( 
.A(n_3602),
.B(n_3004),
.C(n_3127),
.D(n_3204),
.Y(n_3684)
);

BUFx2_ASAP7_75t_L g3685 ( 
.A(n_3680),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3657),
.B(n_3346),
.Y(n_3686)
);

AND2x2_ASAP7_75t_L g3687 ( 
.A(n_3670),
.B(n_3386),
.Y(n_3687)
);

NOR3xp33_ASAP7_75t_L g3688 ( 
.A(n_3646),
.B(n_2938),
.C(n_2909),
.Y(n_3688)
);

AOI222xp33_ASAP7_75t_L g3689 ( 
.A1(n_3643),
.A2(n_3199),
.B1(n_3356),
.B2(n_3355),
.C1(n_3376),
.C2(n_3354),
.Y(n_3689)
);

AOI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_3650),
.A2(n_3004),
.B(n_3380),
.Y(n_3690)
);

AOI221x1_ASAP7_75t_SL g3691 ( 
.A1(n_3684),
.A2(n_3127),
.B1(n_3349),
.B2(n_3372),
.C(n_3348),
.Y(n_3691)
);

NOR4xp25_ASAP7_75t_L g3692 ( 
.A(n_3645),
.B(n_3673),
.C(n_3678),
.D(n_3651),
.Y(n_3692)
);

AOI222xp33_ASAP7_75t_L g3693 ( 
.A1(n_3647),
.A2(n_3199),
.B1(n_3366),
.B2(n_3359),
.C1(n_3352),
.C2(n_3367),
.Y(n_3693)
);

AOI221xp5_ASAP7_75t_L g3694 ( 
.A1(n_3663),
.A2(n_3644),
.B1(n_3666),
.B2(n_3649),
.C(n_3655),
.Y(n_3694)
);

OAI221xp5_ASAP7_75t_SL g3695 ( 
.A1(n_3683),
.A2(n_3081),
.B1(n_3083),
.B2(n_3160),
.C(n_3157),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3665),
.Y(n_3696)
);

NOR3x1_ASAP7_75t_L g3697 ( 
.A(n_3652),
.B(n_3150),
.C(n_2964),
.Y(n_3697)
);

AOI211xp5_ASAP7_75t_SL g3698 ( 
.A1(n_3677),
.A2(n_2778),
.B(n_2909),
.C(n_2938),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3654),
.Y(n_3699)
);

AND2x2_ASAP7_75t_L g3700 ( 
.A(n_3669),
.B(n_3386),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3668),
.B(n_3363),
.Y(n_3701)
);

NAND3xp33_ASAP7_75t_SL g3702 ( 
.A(n_3662),
.B(n_3676),
.C(n_3648),
.Y(n_3702)
);

NAND4xp25_ASAP7_75t_L g3703 ( 
.A(n_3664),
.B(n_3679),
.C(n_3660),
.D(n_3674),
.Y(n_3703)
);

NAND3xp33_ASAP7_75t_L g3704 ( 
.A(n_3659),
.B(n_2908),
.C(n_2899),
.Y(n_3704)
);

NOR3xp33_ASAP7_75t_L g3705 ( 
.A(n_3658),
.B(n_2778),
.C(n_2953),
.Y(n_3705)
);

AOI221xp5_ASAP7_75t_L g3706 ( 
.A1(n_3653),
.A2(n_3083),
.B1(n_3081),
.B2(n_3378),
.C(n_3371),
.Y(n_3706)
);

NOR4xp25_ASAP7_75t_L g3707 ( 
.A(n_3654),
.B(n_2953),
.C(n_2962),
.D(n_3380),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3667),
.Y(n_3708)
);

NOR2xp33_ASAP7_75t_L g3709 ( 
.A(n_3675),
.B(n_2968),
.Y(n_3709)
);

OAI211xp5_ASAP7_75t_L g3710 ( 
.A1(n_3656),
.A2(n_2902),
.B(n_2984),
.C(n_3159),
.Y(n_3710)
);

NAND4xp25_ASAP7_75t_L g3711 ( 
.A(n_3681),
.B(n_3127),
.C(n_3204),
.D(n_3314),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3672),
.B(n_3406),
.Y(n_3712)
);

NOR3xp33_ASAP7_75t_L g3713 ( 
.A(n_3661),
.B(n_2962),
.C(n_2690),
.Y(n_3713)
);

NOR3xp33_ASAP7_75t_L g3714 ( 
.A(n_3702),
.B(n_3682),
.C(n_3130),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3700),
.B(n_3671),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3696),
.Y(n_3716)
);

OAI211xp5_ASAP7_75t_SL g3717 ( 
.A1(n_3694),
.A2(n_3689),
.B(n_3698),
.C(n_3706),
.Y(n_3717)
);

NAND5xp2_ASAP7_75t_L g3718 ( 
.A(n_3694),
.B(n_2900),
.C(n_3167),
.D(n_3065),
.E(n_3062),
.Y(n_3718)
);

NOR2x1_ASAP7_75t_L g3719 ( 
.A(n_3703),
.B(n_2984),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3708),
.B(n_3692),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3687),
.Y(n_3721)
);

NOR2x1_ASAP7_75t_L g3722 ( 
.A(n_3685),
.B(n_2984),
.Y(n_3722)
);

INVxp33_ASAP7_75t_L g3723 ( 
.A(n_3688),
.Y(n_3723)
);

NOR2x1_ASAP7_75t_L g3724 ( 
.A(n_3711),
.B(n_2984),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3699),
.B(n_3406),
.Y(n_3725)
);

NOR2xp33_ASAP7_75t_L g3726 ( 
.A(n_3701),
.B(n_3421),
.Y(n_3726)
);

OAI22xp33_ASAP7_75t_L g3727 ( 
.A1(n_3686),
.A2(n_2900),
.B1(n_3447),
.B2(n_3446),
.Y(n_3727)
);

OR2x2_ASAP7_75t_L g3728 ( 
.A(n_3712),
.B(n_3704),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3693),
.B(n_3421),
.Y(n_3729)
);

NAND3xp33_ASAP7_75t_L g3730 ( 
.A(n_3713),
.B(n_2932),
.C(n_2930),
.Y(n_3730)
);

AND5x1_ASAP7_75t_L g3731 ( 
.A(n_3706),
.B(n_2678),
.C(n_3105),
.D(n_3204),
.E(n_2967),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3697),
.B(n_3433),
.Y(n_3732)
);

AND3x1_ASAP7_75t_L g3733 ( 
.A(n_3707),
.B(n_3130),
.C(n_3096),
.Y(n_3733)
);

NOR3xp33_ASAP7_75t_L g3734 ( 
.A(n_3710),
.B(n_3130),
.C(n_3096),
.Y(n_3734)
);

NOR2x1_ASAP7_75t_L g3735 ( 
.A(n_3709),
.B(n_2631),
.Y(n_3735)
);

NAND3xp33_ASAP7_75t_L g3736 ( 
.A(n_3695),
.B(n_2932),
.C(n_2930),
.Y(n_3736)
);

NOR2x1_ASAP7_75t_L g3737 ( 
.A(n_3690),
.B(n_2801),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3719),
.B(n_3691),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3721),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3725),
.Y(n_3740)
);

INVx2_ASAP7_75t_SL g3741 ( 
.A(n_3728),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3716),
.Y(n_3742)
);

AND2x2_ASAP7_75t_L g3743 ( 
.A(n_3715),
.B(n_3705),
.Y(n_3743)
);

NOR2xp33_ASAP7_75t_L g3744 ( 
.A(n_3723),
.B(n_3433),
.Y(n_3744)
);

NOR3xp33_ASAP7_75t_L g3745 ( 
.A(n_3720),
.B(n_3138),
.C(n_3096),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3726),
.B(n_3453),
.Y(n_3746)
);

NOR3xp33_ASAP7_75t_L g3747 ( 
.A(n_3717),
.B(n_3141),
.C(n_3138),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3729),
.Y(n_3748)
);

NOR2x1_ASAP7_75t_L g3749 ( 
.A(n_3722),
.B(n_3727),
.Y(n_3749)
);

NOR2xp33_ASAP7_75t_L g3750 ( 
.A(n_3718),
.B(n_3446),
.Y(n_3750)
);

INVxp67_ASAP7_75t_L g3751 ( 
.A(n_3714),
.Y(n_3751)
);

NAND4xp25_ASAP7_75t_L g3752 ( 
.A(n_3724),
.B(n_2959),
.C(n_2941),
.D(n_2948),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_SL g3753 ( 
.A1(n_3735),
.A2(n_3381),
.B(n_3161),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_SL g3754 ( 
.A(n_3733),
.B(n_3105),
.Y(n_3754)
);

NOR2x1_ASAP7_75t_L g3755 ( 
.A(n_3737),
.B(n_3730),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3732),
.Y(n_3756)
);

NOR3xp33_ASAP7_75t_L g3757 ( 
.A(n_3741),
.B(n_3736),
.C(n_3734),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3739),
.Y(n_3758)
);

NOR2x1_ASAP7_75t_L g3759 ( 
.A(n_3742),
.B(n_3733),
.Y(n_3759)
);

AND3x2_ASAP7_75t_L g3760 ( 
.A(n_3751),
.B(n_3731),
.C(n_3173),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3747),
.B(n_3453),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3740),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3748),
.B(n_3447),
.Y(n_3763)
);

OR2x6_ASAP7_75t_L g3764 ( 
.A(n_3738),
.B(n_2863),
.Y(n_3764)
);

NOR2x1_ASAP7_75t_L g3765 ( 
.A(n_3749),
.B(n_2923),
.Y(n_3765)
);

INVx4_ASAP7_75t_L g3766 ( 
.A(n_3743),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3744),
.Y(n_3767)
);

NAND2x1p5_ASAP7_75t_L g3768 ( 
.A(n_3755),
.B(n_2863),
.Y(n_3768)
);

OR2x2_ASAP7_75t_L g3769 ( 
.A(n_3756),
.B(n_3165),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3758),
.Y(n_3770)
);

NOR3xp33_ASAP7_75t_L g3771 ( 
.A(n_3766),
.B(n_3745),
.C(n_3754),
.Y(n_3771)
);

HB1xp67_ASAP7_75t_L g3772 ( 
.A(n_3762),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3763),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3767),
.Y(n_3774)
);

INVx3_ASAP7_75t_SL g3775 ( 
.A(n_3764),
.Y(n_3775)
);

OR2x6_ASAP7_75t_L g3776 ( 
.A(n_3764),
.B(n_3746),
.Y(n_3776)
);

AOI221xp5_ASAP7_75t_L g3777 ( 
.A1(n_3757),
.A2(n_3753),
.B1(n_3750),
.B2(n_3752),
.C(n_3165),
.Y(n_3777)
);

AOI22xp5_ASAP7_75t_L g3778 ( 
.A1(n_3759),
.A2(n_3752),
.B1(n_3105),
.B2(n_3358),
.Y(n_3778)
);

O2A1O1Ixp33_ASAP7_75t_L g3779 ( 
.A1(n_3768),
.A2(n_2934),
.B(n_2936),
.C(n_2939),
.Y(n_3779)
);

AOI221xp5_ASAP7_75t_L g3780 ( 
.A1(n_3761),
.A2(n_3183),
.B1(n_3173),
.B2(n_2965),
.C(n_2963),
.Y(n_3780)
);

NOR2x1p5_ASAP7_75t_L g3781 ( 
.A(n_3770),
.B(n_3769),
.Y(n_3781)
);

NOR3xp33_ASAP7_75t_L g3782 ( 
.A(n_3774),
.B(n_3765),
.C(n_3760),
.Y(n_3782)
);

OAI22x1_ASAP7_75t_L g3783 ( 
.A1(n_3775),
.A2(n_3138),
.B1(n_3168),
.B2(n_3141),
.Y(n_3783)
);

AOI221x1_ASAP7_75t_L g3784 ( 
.A1(n_3771),
.A2(n_2956),
.B1(n_2970),
.B2(n_2969),
.C(n_2966),
.Y(n_3784)
);

BUFx2_ASAP7_75t_L g3785 ( 
.A(n_3772),
.Y(n_3785)
);

XOR2xp5_ASAP7_75t_L g3786 ( 
.A(n_3773),
.B(n_2863),
.Y(n_3786)
);

OAI22xp5_ASAP7_75t_L g3787 ( 
.A1(n_3776),
.A2(n_3147),
.B1(n_3176),
.B2(n_3172),
.Y(n_3787)
);

NOR2x1_ASAP7_75t_L g3788 ( 
.A(n_3785),
.B(n_3776),
.Y(n_3788)
);

OAI22x1_ASAP7_75t_L g3789 ( 
.A1(n_3781),
.A2(n_3778),
.B1(n_3777),
.B2(n_3779),
.Y(n_3789)
);

AOI22xp5_ASAP7_75t_L g3790 ( 
.A1(n_3782),
.A2(n_3780),
.B1(n_3105),
.B2(n_3358),
.Y(n_3790)
);

OAI21x1_ASAP7_75t_L g3791 ( 
.A1(n_3788),
.A2(n_3786),
.B(n_3787),
.Y(n_3791)
);

AOI22xp5_ASAP7_75t_L g3792 ( 
.A1(n_3789),
.A2(n_3783),
.B1(n_3784),
.B2(n_3105),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3791),
.A2(n_3790),
.B(n_2933),
.Y(n_3793)
);

OA21x2_ASAP7_75t_L g3794 ( 
.A1(n_3793),
.A2(n_3792),
.B(n_2924),
.Y(n_3794)
);

OAI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3794),
.A2(n_2967),
.B(n_2869),
.Y(n_3795)
);

O2A1O1Ixp33_ASAP7_75t_L g3796 ( 
.A1(n_3795),
.A2(n_3187),
.B(n_3168),
.C(n_3141),
.Y(n_3796)
);


endmodule