module fake_jpeg_30951_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_0),
.Y(n_6)
);

INVx6_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx12_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_1),
.B(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_18),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_6),
.B(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_10),
.B(n_5),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_20),
.B(n_11),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_7),
.A2(n_0),
.B(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_9),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_26),
.B(n_4),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_11),
.C(n_12),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_29),
.B(n_31),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_23),
.B(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_12),
.B1(n_5),
.B2(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_38),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_9),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_9),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_9),
.C(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI311xp33_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_43),
.A3(n_44),
.B(n_40),
.C(n_8),
.Y(n_46)
);


endmodule