module fake_aes_3957_n_434 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_434, n_538);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_434;
output n_538;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_62), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_8), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_67), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_28), .Y(n_79) );
OR2x2_ASAP7_75t_L g80 ( .A(n_44), .B(n_23), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_74), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_53), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_20), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_4), .Y(n_84) );
CKINVDCx16_ASAP7_75t_R g85 ( .A(n_35), .Y(n_85) );
INVx1_ASAP7_75t_SL g86 ( .A(n_71), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_60), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_33), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_75), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_18), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_25), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_66), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_54), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_11), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_45), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_34), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_50), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_69), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_7), .Y(n_99) );
INVx3_ASAP7_75t_L g100 ( .A(n_7), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_9), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_0), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_47), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_29), .Y(n_104) );
INVxp33_ASAP7_75t_SL g105 ( .A(n_55), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_36), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_26), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_4), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_100), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_100), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_78), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_85), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_85), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_100), .Y(n_115) );
AND2x6_ASAP7_75t_L g116 ( .A(n_78), .B(n_37), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_101), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_78), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_100), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_104), .Y(n_120) );
OA21x2_ASAP7_75t_L g121 ( .A1(n_76), .A2(n_32), .B(n_72), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_76), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_101), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_106), .B(n_0), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_84), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_104), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_104), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_79), .B(n_1), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_87), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
NOR2xp33_ASAP7_75t_R g132 ( .A(n_93), .B(n_38), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_108), .Y(n_133) );
OR2x6_ASAP7_75t_L g134 ( .A(n_124), .B(n_77), .Y(n_134) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_122), .A2(n_109), .B1(n_77), .B2(n_94), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_110), .B(n_81), .Y(n_136) );
NAND2xp33_ASAP7_75t_L g137 ( .A(n_116), .B(n_80), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_120), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_110), .B(n_103), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_120), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_120), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_110), .B(n_109), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_117), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_110), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_115), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_115), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
INVxp67_ASAP7_75t_L g149 ( .A(n_123), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_116), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_120), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_120), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_115), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_127), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
AO22x2_ASAP7_75t_L g158 ( .A1(n_122), .A2(n_82), .B1(n_91), .B2(n_92), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_111), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_119), .Y(n_160) );
OR2x6_ASAP7_75t_L g161 ( .A(n_134), .B(n_94), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_134), .A2(n_130), .B1(n_113), .B2(n_114), .Y(n_162) );
INVx1_ASAP7_75t_SL g163 ( .A(n_139), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
OR2x2_ASAP7_75t_L g167 ( .A(n_134), .B(n_131), .Y(n_167) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
NOR2xp67_ASAP7_75t_L g169 ( .A(n_149), .B(n_119), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_143), .Y(n_170) );
BUFx12f_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_159), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_159), .Y(n_173) );
BUFx12f_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_142), .B(n_131), .Y(n_175) );
NOR3xp33_ASAP7_75t_SL g176 ( .A(n_136), .B(n_128), .C(n_102), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_159), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_158), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_142), .B(n_129), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_146), .B(n_99), .Y(n_181) );
BUFx8_ASAP7_75t_SL g182 ( .A(n_136), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_158), .B(n_129), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_146), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_147), .B(n_89), .Y(n_188) );
NOR2xp33_ASAP7_75t_R g189 ( .A(n_137), .B(n_125), .Y(n_189) );
INVx5_ASAP7_75t_L g190 ( .A(n_150), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_147), .Y(n_191) );
NOR3xp33_ASAP7_75t_SL g192 ( .A(n_154), .B(n_102), .C(n_99), .Y(n_192) );
INVx6_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_147), .B(n_129), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_147), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_182), .Y(n_196) );
BUFx8_ASAP7_75t_SL g197 ( .A(n_170), .Y(n_197) );
OR2x6_ASAP7_75t_L g198 ( .A(n_161), .B(n_158), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_170), .Y(n_200) );
INVx3_ASAP7_75t_SL g201 ( .A(n_161), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_165), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
INVxp67_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_168), .B(n_154), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_165), .Y(n_206) );
NOR2x1_ASAP7_75t_SL g207 ( .A(n_161), .B(n_80), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_162), .B(n_133), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_175), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_171), .Y(n_210) );
AOI22xp33_ASAP7_75t_SL g211 ( .A1(n_168), .A2(n_158), .B1(n_105), .B2(n_116), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_186), .A2(n_192), .B(n_176), .C(n_183), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_168), .A2(n_144), .B1(n_148), .B2(n_153), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_175), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_175), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_167), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_177), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_163), .B(n_144), .Y(n_220) );
INVx5_ASAP7_75t_L g221 ( .A(n_174), .Y(n_221) );
INVx5_ASAP7_75t_L g222 ( .A(n_174), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_167), .Y(n_223) );
O2A1O1Ixp5_ASAP7_75t_L g224 ( .A1(n_188), .A2(n_148), .B(n_153), .C(n_160), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_166), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_180), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_177), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_179), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_164), .B(n_135), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_220), .Y(n_230) );
NAND2xp33_ASAP7_75t_L g231 ( .A(n_201), .B(n_166), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_199), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_220), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_221), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_198), .A2(n_178), .B1(n_183), .B2(n_186), .Y(n_235) );
OAI221xp5_ASAP7_75t_L g236 ( .A1(n_214), .A2(n_169), .B1(n_178), .B2(n_194), .C(n_191), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_218), .B(n_181), .Y(n_237) );
BUFx10_ASAP7_75t_L g238 ( .A(n_198), .Y(n_238) );
NAND3xp33_ASAP7_75t_SL g239 ( .A(n_200), .B(n_189), .C(n_132), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_223), .B(n_181), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_209), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_221), .B(n_181), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_198), .B(n_185), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_199), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_198), .B(n_185), .Y(n_247) );
NOR3xp33_ASAP7_75t_SL g248 ( .A(n_196), .B(n_95), .C(n_83), .Y(n_248) );
BUFx4f_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_197), .Y(n_250) );
CKINVDCx8_ASAP7_75t_R g251 ( .A(n_196), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_204), .A2(n_173), .B1(n_172), .B2(n_179), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_221), .B(n_185), .Y(n_253) );
NAND2x1_ASAP7_75t_L g254 ( .A(n_219), .B(n_172), .Y(n_254) );
AOI21xp33_ASAP7_75t_SL g255 ( .A1(n_208), .A2(n_1), .B(n_2), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_230), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_233), .A2(n_214), .B1(n_216), .B2(n_217), .C(n_229), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_236), .A2(n_224), .B(n_205), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_235), .A2(n_211), .B1(n_226), .B2(n_205), .Y(n_259) );
OAI221xp5_ASAP7_75t_L g260 ( .A1(n_248), .A2(n_210), .B1(n_213), .B2(n_215), .C(n_221), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_238), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_241), .Y(n_262) );
OAI221xp5_ASAP7_75t_L g263 ( .A1(n_255), .A2(n_213), .B1(n_222), .B2(n_184), .C(n_187), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_244), .A2(n_197), .B1(n_222), .B2(n_187), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_244), .B(n_207), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_238), .Y(n_266) );
AOI222xp33_ASAP7_75t_L g267 ( .A1(n_249), .A2(n_222), .B1(n_160), .B2(n_108), .C1(n_92), .C2(n_91), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_232), .A2(n_121), .B(n_227), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_242), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_237), .A2(n_222), .B1(n_227), .B2(n_228), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_232), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_247), .B(n_222), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_246), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_238), .B(n_219), .Y(n_274) );
AOI222xp33_ASAP7_75t_L g275 ( .A1(n_249), .A2(n_108), .B1(n_82), .B2(n_96), .C1(n_97), .C2(n_116), .Y(n_275) );
BUFx6f_ASAP7_75t_SL g276 ( .A(n_243), .Y(n_276) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_246), .A2(n_126), .B(n_112), .Y(n_277) );
OAI221xp5_ASAP7_75t_L g278 ( .A1(n_259), .A2(n_249), .B1(n_240), .B2(n_251), .C(n_239), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_277), .Y(n_279) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_267), .B(n_231), .C(n_127), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_269), .Y(n_281) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_258), .A2(n_252), .B(n_126), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_269), .Y(n_284) );
AOI21x1_ASAP7_75t_L g285 ( .A1(n_268), .A2(n_254), .B(n_112), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_257), .A2(n_250), .B1(n_108), .B2(n_243), .C(n_245), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_256), .Y(n_287) );
OAI321xp33_ASAP7_75t_L g288 ( .A1(n_260), .A2(n_108), .A3(n_97), .B1(n_96), .B2(n_107), .C(n_234), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_277), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_277), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_256), .B(n_243), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_277), .Y(n_292) );
NAND4xp25_ASAP7_75t_L g293 ( .A(n_267), .B(n_112), .C(n_118), .D(n_126), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_265), .B(n_234), .Y(n_294) );
OAI211xp5_ASAP7_75t_L g295 ( .A1(n_275), .A2(n_251), .B(n_250), .C(n_88), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_259), .A2(n_247), .B1(n_253), .B2(n_231), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_272), .B(n_253), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_271), .Y(n_298) );
NAND4xp25_ASAP7_75t_L g299 ( .A(n_264), .B(n_118), .C(n_98), .D(n_86), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_271), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_281), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_281), .B(n_273), .Y(n_302) );
AOI211xp5_ASAP7_75t_L g303 ( .A1(n_299), .A2(n_265), .B(n_262), .C(n_272), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_284), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_284), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_279), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_279), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_287), .B(n_274), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_298), .B(n_270), .Y(n_310) );
OAI31xp33_ASAP7_75t_SL g311 ( .A1(n_280), .A2(n_274), .A3(n_263), .B(n_253), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_298), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_280), .B(n_270), .C(n_127), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_283), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_296), .A2(n_276), .B1(n_266), .B2(n_261), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_289), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_289), .Y(n_317) );
NOR4xp25_ASAP7_75t_L g318 ( .A(n_278), .B(n_118), .C(n_98), .D(n_90), .Y(n_318) );
OAI33xp33_ASAP7_75t_L g319 ( .A1(n_299), .A2(n_2), .A3(n_3), .B1(n_5), .B2(n_6), .B3(n_8), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_300), .B(n_273), .Y(n_320) );
BUFx12f_ASAP7_75t_L g321 ( .A(n_297), .Y(n_321) );
OAI33xp33_ASAP7_75t_L g322 ( .A1(n_293), .A2(n_3), .A3(n_5), .B1(n_6), .B2(n_9), .B3(n_10), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_300), .B(n_261), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_291), .B(n_266), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_294), .B(n_266), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_283), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_290), .Y(n_327) );
AND2x2_ASAP7_75t_SL g328 ( .A(n_290), .B(n_261), .Y(n_328) );
XNOR2xp5_ASAP7_75t_L g329 ( .A(n_295), .B(n_10), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_292), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_297), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_292), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_317), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_307), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_301), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_331), .B(n_286), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_301), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_317), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_326), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_323), .B(n_108), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_304), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_303), .A2(n_276), .B1(n_261), .B2(n_288), .Y(n_342) );
OAI33xp33_ASAP7_75t_L g343 ( .A1(n_304), .A2(n_293), .A3(n_12), .B1(n_13), .B2(n_14), .B3(n_15), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_305), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_306), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_312), .B(n_282), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_303), .A2(n_276), .B1(n_282), .B2(n_116), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_326), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_309), .B(n_282), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_302), .B(n_11), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_307), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_13), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_319), .B(n_14), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_302), .B(n_15), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_313), .B(n_285), .Y(n_358) );
INVxp67_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_308), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
NAND2xp33_ASAP7_75t_R g363 ( .A(n_310), .B(n_121), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_323), .B(n_16), .Y(n_364) );
OAI33xp33_ASAP7_75t_L g365 ( .A1(n_324), .A2(n_16), .A3(n_157), .B1(n_156), .B2(n_152), .B3(n_155), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_320), .B(n_332), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_332), .B(n_285), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_316), .B(n_127), .Y(n_368) );
NOR2x1_ASAP7_75t_L g369 ( .A(n_313), .B(n_121), .Y(n_369) );
NAND2xp33_ASAP7_75t_R g370 ( .A(n_310), .B(n_121), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_321), .B(n_17), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_316), .B(n_228), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_320), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_330), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_330), .B(n_268), .Y(n_375) );
NAND2xp33_ASAP7_75t_L g376 ( .A(n_315), .B(n_116), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_328), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_321), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_373), .B(n_328), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_343), .B(n_322), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_342), .A2(n_325), .B1(n_329), .B2(n_314), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_356), .A2(n_318), .B1(n_329), .B2(n_138), .C(n_140), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_335), .Y(n_384) );
OR4x1_ASAP7_75t_L g385 ( .A(n_377), .B(n_311), .C(n_21), .D(n_22), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_356), .A2(n_140), .B1(n_138), .B2(n_145), .C(n_151), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_340), .B(n_116), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_337), .B(n_116), .Y(n_388) );
AOI21xp33_ASAP7_75t_SL g389 ( .A1(n_379), .A2(n_19), .B(n_24), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_359), .B(n_27), .Y(n_390) );
BUFx2_ASAP7_75t_L g391 ( .A(n_339), .Y(n_391) );
AND3x2_ASAP7_75t_L g392 ( .A(n_371), .B(n_157), .C(n_156), .Y(n_392) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_338), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_341), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_333), .Y(n_395) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_355), .A2(n_157), .B(n_156), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_348), .A2(n_225), .B1(n_212), .B2(n_206), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_349), .B(n_366), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_333), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_344), .Y(n_400) );
AOI211xp5_ASAP7_75t_L g401 ( .A1(n_376), .A2(n_141), .B(n_152), .C(n_155), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_345), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_334), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_334), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_346), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_350), .B(n_155), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_364), .B(n_30), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_352), .B(n_138), .C(n_140), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_379), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_372), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_358), .Y(n_411) );
BUFx2_ASAP7_75t_L g412 ( .A(n_374), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_378), .B(n_362), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_351), .B(n_152), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_353), .Y(n_416) );
AOI322xp5_ASAP7_75t_L g417 ( .A1(n_336), .A2(n_141), .A3(n_191), .B1(n_184), .B2(n_138), .C1(n_145), .C2(n_151), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_353), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_358), .Y(n_419) );
AOI31xp33_ASAP7_75t_L g420 ( .A1(n_365), .A2(n_141), .A3(n_39), .B(n_40), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_357), .A2(n_225), .B(n_212), .Y(n_421) );
A2O1A1Ixp33_ASAP7_75t_L g422 ( .A1(n_376), .A2(n_195), .B(n_212), .C(n_206), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_347), .A2(n_138), .B1(n_140), .B2(n_145), .C(n_151), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_354), .Y(n_424) );
OAI33xp33_ASAP7_75t_L g425 ( .A1(n_375), .A2(n_173), .A3(n_195), .B1(n_42), .B2(n_43), .B3(n_46), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_354), .B(n_31), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_367), .A2(n_138), .B1(n_140), .B2(n_145), .C(n_151), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_360), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_367), .A2(n_140), .B(n_145), .Y(n_429) );
NAND2xp33_ASAP7_75t_L g430 ( .A(n_360), .B(n_225), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_363), .A2(n_145), .B1(n_151), .B2(n_206), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_368), .B(n_151), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_393), .B(n_368), .Y(n_433) );
UNKNOWN g434 ( );
O2A1O1Ixp33_ASAP7_75t_L g435 ( .A1(n_420), .A2(n_369), .B(n_370), .C(n_363), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_384), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_394), .Y(n_437) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_391), .B(n_370), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_398), .B(n_41), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_382), .A2(n_381), .B1(n_390), .B2(n_407), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_402), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_405), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_412), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_410), .B(n_48), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_393), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_395), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_399), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_380), .B(n_49), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_411), .B(n_225), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_403), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_404), .Y(n_454) );
XOR2x2_ASAP7_75t_L g455 ( .A(n_409), .B(n_51), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_416), .B(n_52), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_428), .B(n_56), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_424), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_411), .B(n_57), .Y(n_460) );
XOR2x2_ASAP7_75t_L g461 ( .A(n_390), .B(n_58), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_419), .B(n_59), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_381), .B(n_61), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_419), .B(n_63), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_386), .B(n_212), .C(n_206), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_415), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_421), .A2(n_203), .B1(n_202), .B2(n_199), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_406), .B(n_64), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
XNOR2xp5_ASAP7_75t_L g470 ( .A(n_392), .B(n_65), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_423), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_392), .B(n_68), .Y(n_472) );
AOI21xp33_ASAP7_75t_SL g473 ( .A1(n_385), .A2(n_70), .B(n_73), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_408), .B(n_199), .Y(n_474) );
XNOR2xp5_ASAP7_75t_L g475 ( .A(n_455), .B(n_401), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_447), .B(n_429), .Y(n_476) );
OAI211xp5_ASAP7_75t_L g477 ( .A1(n_441), .A2(n_389), .B(n_422), .C(n_431), .Y(n_477) );
XNOR2xp5_ASAP7_75t_L g478 ( .A(n_455), .B(n_397), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_463), .A2(n_425), .B(n_397), .C(n_396), .Y(n_479) );
XOR2xp5_ASAP7_75t_L g480 ( .A(n_461), .B(n_387), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_436), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_437), .Y(n_482) );
AOI21xp33_ASAP7_75t_L g483 ( .A1(n_471), .A2(n_426), .B(n_432), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_433), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_444), .Y(n_485) );
NAND3xp33_ASAP7_75t_L g486 ( .A(n_471), .B(n_417), .C(n_427), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_442), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_457), .B(n_388), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_443), .B(n_425), .Y(n_490) );
AOI321xp33_ASAP7_75t_L g491 ( .A1(n_438), .A2(n_202), .A3(n_203), .B1(n_190), .B2(n_193), .C(n_166), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_448), .B(n_202), .Y(n_492) );
NAND3x1_ASAP7_75t_SL g493 ( .A(n_461), .B(n_202), .C(n_203), .Y(n_493) );
AOI211x1_ASAP7_75t_SL g494 ( .A1(n_434), .A2(n_203), .B(n_166), .C(n_190), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_466), .B(n_166), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_433), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_473), .B(n_190), .C(n_193), .Y(n_498) );
OAI31xp33_ASAP7_75t_SL g499 ( .A1(n_460), .A2(n_190), .A3(n_193), .B(n_465), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_435), .A2(n_190), .B1(n_193), .B2(n_469), .C(n_470), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_433), .B(n_450), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_485), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_486), .A2(n_435), .B1(n_449), .B2(n_440), .C(n_453), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_475), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_481), .Y(n_505) );
AOI221xp5_ASAP7_75t_L g506 ( .A1(n_483), .A2(n_459), .B1(n_453), .B2(n_454), .C(n_464), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_490), .B(n_459), .Y(n_507) );
NOR2x1p5_ASAP7_75t_L g508 ( .A(n_498), .B(n_472), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_501), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_499), .A2(n_460), .B(n_467), .C(n_445), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_490), .B(n_454), .Y(n_511) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_495), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_484), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_482), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_487), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_488), .Y(n_516) );
NAND4xp25_ASAP7_75t_L g517 ( .A(n_500), .B(n_451), .C(n_462), .D(n_460), .Y(n_517) );
OAI221xp5_ASAP7_75t_L g518 ( .A1(n_478), .A2(n_452), .B1(n_468), .B2(n_458), .C(n_456), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_483), .A2(n_452), .B1(n_474), .B2(n_496), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_497), .B(n_492), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_477), .A2(n_480), .B1(n_476), .B2(n_479), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_491), .B(n_476), .Y(n_522) );
OR3x2_ASAP7_75t_L g523 ( .A(n_493), .B(n_494), .C(n_489), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_489), .B(n_409), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_485), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_504), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_513), .B(n_509), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_502), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_521), .A2(n_503), .B1(n_522), .B2(n_517), .Y(n_529) );
OAI211xp5_ASAP7_75t_SL g530 ( .A1(n_506), .A2(n_519), .B(n_518), .C(n_510), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_529), .B(n_512), .C(n_507), .Y(n_531) );
OA22x2_ASAP7_75t_L g532 ( .A1(n_526), .A2(n_525), .B1(n_511), .B2(n_509), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_528), .Y(n_533) );
OAI221xp5_ASAP7_75t_L g534 ( .A1(n_531), .A2(n_530), .B1(n_527), .B2(n_524), .C(n_512), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_533), .Y(n_535) );
OAI222xp33_ASAP7_75t_L g536 ( .A1(n_534), .A2(n_532), .B1(n_505), .B2(n_516), .C1(n_515), .C2(n_514), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_536), .A2(n_535), .B1(n_512), .B2(n_508), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_537), .A2(n_520), .B(n_523), .Y(n_538) );
endmodule