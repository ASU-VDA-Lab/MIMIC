module real_aes_8380_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_841;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_316;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_725;
wire n_310;
wire n_455;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_397;
wire n_749;
wire n_358;
wire n_293;
wire n_385;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_753;
wire n_314;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_SL g337 ( .A1(n_0), .A2(n_237), .B1(n_338), .B2(n_342), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_1), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_2), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_3), .A2(n_246), .B1(n_625), .B2(n_626), .Y(n_624) );
AOI222xp33_ASAP7_75t_L g410 ( .A1(n_4), .A2(n_86), .B1(n_260), .B2(n_366), .C1(n_411), .C2(n_413), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_5), .A2(n_113), .B1(n_357), .B2(n_409), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_6), .A2(n_24), .B1(n_369), .B2(n_577), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_7), .A2(n_59), .B1(n_370), .B2(n_479), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_8), .B(n_405), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_9), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_10), .A2(n_271), .B1(n_710), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_11), .A2(n_71), .B1(n_601), .B2(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g457 ( .A(n_12), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_13), .A2(n_257), .B1(n_536), .B2(n_753), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_14), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_15), .A2(n_123), .B1(n_536), .B2(n_564), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_16), .A2(n_266), .B1(n_405), .B2(n_620), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_17), .A2(n_144), .B1(n_489), .B2(n_560), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_18), .A2(n_120), .B1(n_487), .B2(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_19), .A2(n_111), .B1(n_407), .B2(n_473), .Y(n_621) );
AOI22xp33_ASAP7_75t_SL g853 ( .A1(n_20), .A2(n_163), .B1(n_472), .B2(n_473), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_21), .A2(n_178), .B1(n_306), .B2(n_499), .Y(n_801) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_22), .A2(n_55), .B1(n_710), .B2(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g788 ( .A(n_23), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_25), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_26), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_27), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_28), .A2(n_167), .B1(n_396), .B2(n_529), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_29), .A2(n_274), .B1(n_565), .B2(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_30), .A2(n_240), .B1(n_357), .B2(n_773), .Y(n_793) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_31), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_32), .B(n_555), .Y(n_554) );
AO22x2_ASAP7_75t_L g312 ( .A1(n_33), .A2(n_88), .B1(n_313), .B2(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g839 ( .A(n_33), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_34), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_35), .A2(n_142), .B1(n_528), .B2(n_753), .Y(n_752) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_36), .A2(n_209), .B1(n_366), .B2(n_369), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_37), .A2(n_162), .B1(n_487), .B2(n_530), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_38), .A2(n_157), .B1(n_334), .B2(n_345), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_39), .A2(n_259), .B1(n_323), .B2(n_645), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_40), .A2(n_121), .B1(n_388), .B2(n_631), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_41), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_42), .A2(n_247), .B1(n_388), .B2(n_389), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_43), .A2(n_189), .B1(n_472), .B2(n_557), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_44), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_45), .Y(n_480) );
INVx1_ASAP7_75t_L g771 ( .A(n_46), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_47), .A2(n_175), .B1(n_370), .B2(n_557), .Y(n_556) );
AO22x2_ASAP7_75t_L g316 ( .A1(n_48), .A2(n_91), .B1(n_313), .B2(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g840 ( .A(n_48), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_49), .A2(n_128), .B1(n_358), .B2(n_362), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_50), .Y(n_497) );
INVx1_ASAP7_75t_L g736 ( .A(n_51), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_52), .A2(n_270), .B1(n_374), .B2(n_553), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_53), .A2(n_159), .B1(n_345), .B2(n_347), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_54), .Y(n_549) );
AOI22xp33_ASAP7_75t_SL g714 ( .A1(n_56), .A2(n_60), .B1(n_715), .B2(n_716), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_57), .A2(n_255), .B1(n_413), .B2(n_851), .Y(n_850) );
AOI222xp33_ASAP7_75t_L g653 ( .A1(n_58), .A2(n_188), .B1(n_262), .B2(n_366), .C1(n_411), .C2(n_482), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_61), .Y(n_599) );
AOI22xp5_ASAP7_75t_SL g329 ( .A1(n_62), .A2(n_156), .B1(n_330), .B2(n_334), .Y(n_329) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_63), .A2(n_256), .B1(n_323), .B2(n_631), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_64), .A2(n_268), .B1(n_616), .B2(n_617), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_65), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_66), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_67), .A2(n_222), .B1(n_384), .B2(n_386), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_68), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_69), .A2(n_278), .B1(n_532), .B2(n_533), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_70), .A2(n_195), .B1(n_396), .B2(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_72), .A2(n_182), .B1(n_347), .B2(n_560), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_73), .A2(n_198), .B1(n_533), .B2(n_560), .Y(n_559) );
AOI22xp5_ASAP7_75t_SL g305 ( .A1(n_74), .A2(n_137), .B1(n_306), .B2(n_323), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_75), .A2(n_221), .B1(n_374), .B2(n_377), .Y(n_373) );
XNOR2x2_ASAP7_75t_L g380 ( .A(n_76), .B(n_381), .Y(n_380) );
AO22x2_ASAP7_75t_L g503 ( .A1(n_77), .A2(n_504), .B1(n_537), .B2(n_538), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_77), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_78), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_79), .A2(n_235), .B1(n_528), .B2(n_529), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_80), .Y(n_467) );
AOI211xp5_ASAP7_75t_L g464 ( .A1(n_81), .A2(n_465), .B(n_466), .C(n_476), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_82), .A2(n_104), .B1(n_536), .B2(n_718), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_83), .Y(n_875) );
AO22x1_ASAP7_75t_L g877 ( .A1(n_83), .A2(n_875), .B1(n_878), .B2(n_879), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_84), .A2(n_145), .B1(n_564), .B2(n_565), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_85), .A2(n_99), .B1(n_777), .B2(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g781 ( .A(n_87), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_89), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_90), .A2(n_135), .B1(n_577), .B2(n_578), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_92), .A2(n_203), .B1(n_348), .B2(n_530), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_93), .A2(n_661), .B1(n_694), .B2(n_695), .Y(n_660) );
INVx1_ASAP7_75t_L g694 ( .A(n_93), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_94), .Y(n_654) );
INVx1_ASAP7_75t_L g293 ( .A(n_95), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_96), .A2(n_611), .B1(n_635), .B2(n_636), .Y(n_610) );
INVx1_ASAP7_75t_L g636 ( .A(n_96), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_97), .A2(n_124), .B1(n_392), .B2(n_393), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_98), .A2(n_202), .B1(n_560), .B2(n_749), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_100), .A2(n_205), .B1(n_487), .B2(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g290 ( .A(n_101), .Y(n_290) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_102), .A2(n_143), .B1(n_358), .B2(n_366), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_103), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_105), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g821 ( .A1(n_106), .A2(n_168), .B1(n_634), .B2(n_822), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_107), .A2(n_185), .B1(n_396), .B2(n_397), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_108), .A2(n_241), .B1(n_645), .B2(n_728), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_109), .B(n_553), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_110), .A2(n_226), .B1(n_683), .B2(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g428 ( .A(n_112), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_114), .A2(n_158), .B1(n_557), .B2(n_649), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_115), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_116), .Y(n_573) );
AOI211xp5_ASAP7_75t_L g719 ( .A1(n_117), .A2(n_601), .B(n_720), .C(n_725), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_118), .A2(n_150), .B1(n_491), .B2(n_633), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g895 ( .A1(n_119), .A2(n_138), .B1(n_273), .B2(n_577), .C1(n_617), .C2(n_669), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_122), .A2(n_225), .B1(n_338), .B2(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g458 ( .A(n_125), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_126), .A2(n_204), .B1(n_689), .B2(n_690), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_127), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_129), .A2(n_279), .B1(n_393), .B2(n_749), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_130), .A2(n_181), .B1(n_357), .B2(n_362), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_131), .A2(n_212), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_132), .A2(n_276), .B1(n_589), .B2(n_592), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_133), .A2(n_166), .B1(n_323), .B2(n_891), .Y(n_890) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_134), .Y(n_670) );
AOI22xp5_ASAP7_75t_SL g568 ( .A1(n_136), .A2(n_569), .B1(n_603), .B2(n_604), .Y(n_568) );
INVx1_ASAP7_75t_L g604 ( .A(n_136), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_139), .A2(n_843), .B1(n_844), .B2(n_864), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_139), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_140), .B(n_405), .Y(n_470) );
INVx2_ASAP7_75t_L g294 ( .A(n_141), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_146), .Y(n_702) );
INVx1_ASAP7_75t_L g744 ( .A(n_147), .Y(n_744) );
AOI22xp33_ASAP7_75t_SL g860 ( .A1(n_148), .A2(n_180), .B1(n_491), .B2(n_589), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_149), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_151), .A2(n_208), .B1(n_407), .B2(n_409), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_152), .Y(n_572) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_153), .Y(n_462) );
AND2x6_ASAP7_75t_L g289 ( .A(n_154), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_154), .Y(n_833) );
AO22x2_ASAP7_75t_L g320 ( .A1(n_155), .A2(n_232), .B1(n_313), .B2(n_317), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_160), .Y(n_704) );
INVx1_ASAP7_75t_L g745 ( .A(n_161), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_164), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_165), .A2(n_201), .B1(n_306), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_169), .A2(n_230), .B1(n_374), .B2(n_620), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_170), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_171), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_172), .Y(n_664) );
AOI22xp33_ASAP7_75t_SL g779 ( .A1(n_173), .A2(n_263), .B1(n_345), .B2(n_749), .Y(n_779) );
OA22x2_ASAP7_75t_L g730 ( .A1(n_174), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_174), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_176), .Y(n_675) );
AOI22xp33_ASAP7_75t_SL g755 ( .A1(n_177), .A2(n_283), .B1(n_397), .B2(n_533), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_179), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_183), .A2(n_261), .B1(n_535), .B2(n_536), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_184), .A2(n_252), .B1(n_564), .B2(n_565), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_186), .A2(n_215), .B1(n_882), .B2(n_883), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_187), .Y(n_567) );
AO22x2_ASAP7_75t_L g322 ( .A1(n_190), .A2(n_250), .B1(n_313), .B2(n_314), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_191), .A2(n_218), .B1(n_413), .B2(n_475), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_192), .A2(n_219), .B1(n_587), .B2(n_601), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_193), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_194), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_196), .A2(n_253), .B1(n_482), .B2(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g500 ( .A(n_197), .Y(n_500) );
INVx1_ASAP7_75t_L g423 ( .A(n_199), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_200), .Y(n_849) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_206), .A2(n_280), .B1(n_672), .B2(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g454 ( .A(n_207), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_210), .B(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_211), .A2(n_254), .B1(n_306), .B2(n_334), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_213), .B(n_342), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_214), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_216), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_217), .A2(n_251), .B1(n_528), .B2(n_530), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_220), .A2(n_272), .B1(n_389), .B2(n_393), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_223), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_224), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_227), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_228), .A2(n_239), .B1(n_777), .B2(n_778), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_229), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_231), .A2(n_248), .B1(n_362), .B2(n_472), .Y(n_894) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_232), .B(n_838), .Y(n_837) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_233), .A2(n_287), .B(n_295), .C(n_841), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_234), .B(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g594 ( .A(n_236), .Y(n_594) );
INVx1_ASAP7_75t_L g741 ( .A(n_238), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_242), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_243), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_244), .A2(n_258), .B1(n_405), .B2(n_553), .Y(n_647) );
INVx1_ASAP7_75t_L g738 ( .A(n_245), .Y(n_738) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_249), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g836 ( .A(n_250), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_264), .Y(n_792) );
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_265), .A2(n_285), .B1(n_393), .B2(n_499), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_267), .Y(n_673) );
INVx1_ASAP7_75t_L g313 ( .A(n_269), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_269), .Y(n_315) );
INVx1_ASAP7_75t_L g790 ( .A(n_275), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_277), .A2(n_284), .B1(n_633), .B2(n_686), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_281), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_282), .Y(n_706) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_290), .Y(n_832) );
OA21x2_ASAP7_75t_L g873 ( .A1(n_291), .A2(n_831), .B(n_874), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_657), .B1(n_826), .B2(n_827), .C(n_828), .Y(n_295) );
INVxp67_ASAP7_75t_L g826 ( .A(n_296), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B1(n_541), .B2(n_656), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
XOR2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_414), .Y(n_298) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_379), .B2(n_380), .Y(n_301) );
OAI22xp5_ASAP7_75t_SL g416 ( .A1(n_302), .A2(n_303), .B1(n_417), .B2(n_418), .Y(n_416) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
XOR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_378), .Y(n_303) );
NAND4xp75_ASAP7_75t_SL g304 ( .A(n_305), .B(n_329), .C(n_336), .D(n_350), .Y(n_304) );
INVx1_ASAP7_75t_L g494 ( .A(n_306), .Y(n_494) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_SL g689 ( .A(n_307), .Y(n_689) );
INVx4_ASAP7_75t_L g728 ( .A(n_307), .Y(n_728) );
INVx11_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx11_ASAP7_75t_L g385 ( .A(n_308), .Y(n_385) );
AND2x6_ASAP7_75t_L g308 ( .A(n_309), .B(n_318), .Y(n_308) );
AND2x4_ASAP7_75t_L g376 ( .A(n_309), .B(n_349), .Y(n_376) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g424 ( .A(n_310), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_316), .Y(n_310) );
AND2x2_ASAP7_75t_L g328 ( .A(n_311), .B(n_316), .Y(n_328) );
AND2x2_ASAP7_75t_L g332 ( .A(n_311), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_316), .Y(n_355) );
AND2x2_ASAP7_75t_L g361 ( .A(n_312), .B(n_320), .Y(n_361) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g317 ( .A(n_315), .Y(n_317) );
INVx2_ASAP7_75t_L g333 ( .A(n_316), .Y(n_333) );
INVx1_ASAP7_75t_L g372 ( .A(n_316), .Y(n_372) );
AND2x2_ASAP7_75t_L g331 ( .A(n_318), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g335 ( .A(n_318), .B(n_328), .Y(n_335) );
AND2x6_ASAP7_75t_L g354 ( .A(n_318), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
AND2x2_ASAP7_75t_L g349 ( .A(n_319), .B(n_322), .Y(n_349) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g326 ( .A(n_320), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_320), .B(n_322), .Y(n_341) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g327 ( .A(n_322), .Y(n_327) );
INVx1_ASAP7_75t_L g360 ( .A(n_322), .Y(n_360) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g396 ( .A(n_324), .Y(n_396) );
INVx2_ASAP7_75t_L g528 ( .A(n_324), .Y(n_528) );
INVx4_ASAP7_75t_L g591 ( .A(n_324), .Y(n_591) );
INVx5_ASAP7_75t_L g634 ( .A(n_324), .Y(n_634) );
INVx8_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g346 ( .A(n_326), .B(n_332), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_326), .B(n_328), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_326), .B(n_332), .Y(n_455) );
INVx1_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
AND2x6_ASAP7_75t_L g377 ( .A(n_328), .B(n_349), .Y(n_377) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_328), .B(n_349), .Y(n_403) );
BUFx2_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_331), .Y(n_392) );
INVx2_ASAP7_75t_L g443 ( .A(n_331), .Y(n_443) );
BUFx2_ASAP7_75t_SL g601 ( .A(n_331), .Y(n_601) );
AND2x4_ASAP7_75t_L g339 ( .A(n_332), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g348 ( .A(n_332), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g343 ( .A(n_333), .Y(n_343) );
AND2x2_ASAP7_75t_L g368 ( .A(n_333), .B(n_360), .Y(n_368) );
BUFx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx3_ASAP7_75t_L g386 ( .A(n_335), .Y(n_386) );
INVx6_ASAP7_75t_L g445 ( .A(n_335), .Y(n_445) );
BUFx3_ASAP7_75t_L g715 ( .A(n_335), .Y(n_715) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_344), .Y(n_336) );
BUFx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_SL g389 ( .A(n_339), .Y(n_389) );
INVx1_ASAP7_75t_L g450 ( .A(n_339), .Y(n_450) );
BUFx2_ASAP7_75t_L g489 ( .A(n_339), .Y(n_489) );
BUFx3_ASAP7_75t_L g536 ( .A(n_339), .Y(n_536) );
BUFx3_ASAP7_75t_L g565 ( .A(n_339), .Y(n_565) );
BUFx3_ASAP7_75t_L g587 ( .A(n_339), .Y(n_587) );
BUFx2_ASAP7_75t_SL g626 ( .A(n_339), .Y(n_626) );
AND2x2_ASAP7_75t_L g342 ( .A(n_340), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x6_ASAP7_75t_L g398 ( .A(n_341), .B(n_372), .Y(n_398) );
NAND2x1p5_ASAP7_75t_L g431 ( .A(n_343), .B(n_361), .Y(n_431) );
BUFx2_ASAP7_75t_L g716 ( .A(n_345), .Y(n_716) );
INVx1_ASAP7_75t_L g884 ( .A(n_345), .Y(n_884) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g394 ( .A(n_346), .Y(n_394) );
BUFx3_ASAP7_75t_L g564 ( .A(n_346), .Y(n_564) );
BUFx3_ASAP7_75t_L g628 ( .A(n_346), .Y(n_628) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_347), .Y(n_718) );
BUFx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_348), .Y(n_388) );
INVx2_ASAP7_75t_L g439 ( .A(n_348), .Y(n_439) );
BUFx3_ASAP7_75t_L g533 ( .A(n_348), .Y(n_533) );
BUFx3_ASAP7_75t_L g777 ( .A(n_348), .Y(n_777) );
INVx1_ASAP7_75t_L g425 ( .A(n_349), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_364), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B(n_356), .Y(n_351) );
OAI222xp33_ASAP7_75t_L g701 ( .A1(n_353), .A2(n_702), .B1(n_703), .B2(n_704), .C1(n_705), .C2(n_706), .Y(n_701) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx4_ASAP7_75t_L g412 ( .A(n_354), .Y(n_412) );
INVx2_ASAP7_75t_SL g434 ( .A(n_354), .Y(n_434) );
BUFx3_ASAP7_75t_L g465 ( .A(n_354), .Y(n_465) );
INVx2_ASAP7_75t_L g548 ( .A(n_354), .Y(n_548) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_354), .Y(n_669) );
AND2x4_ASAP7_75t_L g362 ( .A(n_355), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g523 ( .A(n_355), .Y(n_523) );
INVx2_ASAP7_75t_L g483 ( .A(n_357), .Y(n_483) );
BUFx4f_ASAP7_75t_SL g617 ( .A(n_357), .Y(n_617) );
BUFx12f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_358), .Y(n_413) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_358), .Y(n_672) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g367 ( .A(n_361), .B(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g370 ( .A(n_361), .B(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_SL g409 ( .A(n_362), .Y(n_409) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_362), .Y(n_475) );
BUFx3_ASAP7_75t_L g557 ( .A(n_362), .Y(n_557) );
BUFx2_ASAP7_75t_SL g773 ( .A(n_362), .Y(n_773) );
INVx1_ASAP7_75t_L g524 ( .A(n_363), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_373), .Y(n_364) );
INVx4_ASAP7_75t_L g436 ( .A(n_366), .Y(n_436) );
BUFx2_ASAP7_75t_L g851 ( .A(n_366), .Y(n_851) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_367), .Y(n_479) );
BUFx2_ASAP7_75t_L g516 ( .A(n_367), .Y(n_516) );
BUFx4f_ASAP7_75t_SL g577 ( .A(n_367), .Y(n_577) );
BUFx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g408 ( .A(n_370), .Y(n_408) );
BUFx2_ASAP7_75t_L g472 ( .A(n_370), .Y(n_472) );
BUFx2_ASAP7_75t_L g649 ( .A(n_370), .Y(n_649) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_374), .Y(n_710) );
INVx5_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g405 ( .A(n_375), .Y(n_405) );
INVx2_ASAP7_75t_L g555 ( .A(n_375), .Y(n_555) );
INVx2_ASAP7_75t_L g767 ( .A(n_375), .Y(n_767) );
INVx4_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx4f_ASAP7_75t_L g553 ( .A(n_377), .Y(n_553) );
BUFx2_ASAP7_75t_L g620 ( .A(n_377), .Y(n_620) );
INVx1_ASAP7_75t_SL g856 ( .A(n_377), .Y(n_856) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND4xp75_ASAP7_75t_L g381 ( .A(n_382), .B(n_390), .C(n_399), .D(n_410), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_387), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_385), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_SL g535 ( .A(n_385), .Y(n_535) );
INVx4_ASAP7_75t_L g596 ( .A(n_385), .Y(n_596) );
INVx2_ASAP7_75t_L g625 ( .A(n_385), .Y(n_625) );
INVx5_ASAP7_75t_SL g749 ( .A(n_385), .Y(n_749) );
HB1xp67_ASAP7_75t_L g889 ( .A(n_385), .Y(n_889) );
INVx3_ASAP7_75t_L g754 ( .A(n_386), .Y(n_754) );
INVx4_ASAP7_75t_L g488 ( .A(n_388), .Y(n_488) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_392), .Y(n_499) );
BUFx3_ASAP7_75t_L g683 ( .A(n_392), .Y(n_683) );
BUFx3_ASAP7_75t_L g882 ( .A(n_392), .Y(n_882) );
BUFx4f_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g491 ( .A(n_398), .Y(n_491) );
INVx6_ASAP7_75t_SL g530 ( .A(n_398), .Y(n_530) );
INVx1_ASAP7_75t_SL g778 ( .A(n_398), .Y(n_778) );
OA211x2_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B(n_404), .C(n_406), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g511 ( .A(n_402), .Y(n_511) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx3_ASAP7_75t_L g429 ( .A(n_403), .Y(n_429) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx4_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI21xp5_ASAP7_75t_SL g574 ( .A1(n_412), .A2(n_575), .B(n_576), .Y(n_574) );
BUFx4f_ASAP7_75t_L g578 ( .A(n_413), .Y(n_578) );
INVx1_ASAP7_75t_L g705 ( .A(n_413), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_459), .B2(n_460), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
XNOR2x1_ASAP7_75t_L g419 ( .A(n_420), .B(n_458), .Y(n_419) );
AND3x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_437), .C(n_447), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_427), .C(n_432), .Y(n_421) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B(n_426), .Y(n_422) );
INVx2_ASAP7_75t_L g509 ( .A(n_424), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g571 ( .A1(n_424), .A2(n_429), .B1(n_572), .B2(n_573), .Y(n_571) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_424), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_427) );
INVx2_ASAP7_75t_L g469 ( .A(n_429), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_429), .A2(n_508), .B1(n_664), .B2(n_665), .Y(n_663) );
BUFx3_ASAP7_75t_L g739 ( .A(n_429), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_429), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_787) );
INVx4_ASAP7_75t_L g520 ( .A(n_431), .Y(n_520) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_431), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_431), .A2(n_478), .B1(n_744), .B2(n_745), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_435), .B2(n_436), .Y(n_432) );
OAI222xp33_ASAP7_75t_L g666 ( .A1(n_436), .A2(n_667), .B1(n_668), .B2(n_670), .C1(n_671), .C2(n_673), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_442), .Y(n_437) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_440), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g684 ( .A(n_439), .Y(n_684) );
INVx2_ASAP7_75t_L g859 ( .A(n_439), .Y(n_859) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_444), .B1(n_445), .B2(n_446), .Y(n_442) );
INVx3_ASAP7_75t_L g532 ( .A(n_443), .Y(n_532) );
INVx3_ASAP7_75t_L g560 ( .A(n_443), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_445), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_445), .A2(n_594), .B1(n_595), .B2(n_597), .Y(n_593) );
INVx2_ASAP7_75t_L g631 ( .A(n_445), .Y(n_631) );
INVx2_ASAP7_75t_L g645 ( .A(n_445), .Y(n_645) );
INVx2_ASAP7_75t_L g690 ( .A(n_445), .Y(n_690) );
INVx3_ASAP7_75t_L g822 ( .A(n_445), .Y(n_822) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_453), .C(n_456), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_451), .B2(n_452), .Y(n_448) );
BUFx2_ASAP7_75t_R g721 ( .A(n_452), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g502 ( .A(n_455), .Y(n_502) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_503), .B1(n_539), .B2(n_540), .Y(n_460) );
INVx2_ASAP7_75t_L g539 ( .A(n_461), .Y(n_539) );
XNOR2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_484), .Y(n_463) );
INVx3_ASAP7_75t_L g514 ( .A(n_465), .Y(n_514) );
OAI211xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_470), .C(n_471), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_480), .B2(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_479), .Y(n_616) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_492), .C(n_496), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_490), .Y(n_485) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_500), .B2(n_501), .Y(n_496) );
INVx1_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_501), .A2(n_599), .B1(n_600), .B2(n_602), .Y(n_598) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g540 ( .A(n_503), .Y(n_540) );
INVx1_ASAP7_75t_SL g537 ( .A(n_504), .Y(n_537) );
AND2x2_ASAP7_75t_SL g504 ( .A(n_505), .B(n_525), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_512), .C(n_517), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_510), .B2(n_511), .Y(n_506) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_SL g789 ( .A(n_509), .Y(n_789) );
OAI21xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_515), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_521), .B2(n_522), .Y(n_517) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx3_ASAP7_75t_SL g580 ( .A(n_520), .Y(n_580) );
BUFx2_ASAP7_75t_L g582 ( .A(n_522), .Y(n_582) );
CKINVDCx16_ASAP7_75t_R g679 ( .A(n_522), .Y(n_679) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
AND4x1_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .C(n_531), .D(n_534), .Y(n_525) );
BUFx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g592 ( .A(n_530), .Y(n_592) );
BUFx4f_ASAP7_75t_SL g686 ( .A(n_530), .Y(n_686) );
BUFx2_ASAP7_75t_L g891 ( .A(n_530), .Y(n_891) );
INVx1_ASAP7_75t_L g656 ( .A(n_541), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B1(n_607), .B2(n_655), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AO22x2_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_568), .B1(n_605), .B2(n_606), .Y(n_543) );
INVx4_ASAP7_75t_SL g605 ( .A(n_544), .Y(n_605) );
AO22x2_ASAP7_75t_L g638 ( .A1(n_544), .A2(n_605), .B1(n_639), .B2(n_640), .Y(n_638) );
XOR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_567), .Y(n_544) );
NAND3x1_ASAP7_75t_L g545 ( .A(n_546), .B(n_558), .C(n_562), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_551), .Y(n_546) );
OAI21xp5_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_549), .B(n_550), .Y(n_547) );
OAI21xp5_ASAP7_75t_SL g613 ( .A1(n_548), .A2(n_614), .B(n_615), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g770 ( .A1(n_548), .A2(n_771), .B(n_772), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g810 ( .A1(n_548), .A2(n_811), .B(n_812), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .C(n_556), .Y(n_551) );
INVx1_ASAP7_75t_L g712 ( .A(n_553), .Y(n_712) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_566), .Y(n_562) );
INVx1_ASAP7_75t_L g606 ( .A(n_568), .Y(n_606) );
INVx1_ASAP7_75t_L g603 ( .A(n_569), .Y(n_603) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_584), .Y(n_569) );
NOR3xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .C(n_579), .Y(n_570) );
INVx1_ASAP7_75t_L g796 ( .A(n_577), .Y(n_796) );
OAI22xp5_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_579) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_593), .C(n_598), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g723 ( .A(n_592), .Y(n_723) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g655 ( .A(n_607), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_637), .B2(n_638), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_SL g635 ( .A(n_611), .Y(n_635) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_622), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_618), .Y(n_612) );
INVx2_ASAP7_75t_SL g703 ( .A(n_616), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_619), .B(n_621), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_629), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
INVx1_ASAP7_75t_L g693 ( .A(n_628), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
XOR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_654), .Y(n_640) );
NAND4xp75_ASAP7_75t_L g641 ( .A(n_642), .B(n_646), .C(n_650), .D(n_653), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x2_ASAP7_75t_SL g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g827 ( .A(n_657), .Y(n_827) );
XOR2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_758), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_696), .B2(n_757), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g695 ( .A(n_661), .Y(n_695) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_680), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .C(n_674), .Y(n_662) );
OAI21xp33_ASAP7_75t_L g740 ( .A1(n_668), .A2(n_741), .B(n_742), .Y(n_740) );
OAI21xp33_ASAP7_75t_L g791 ( .A1(n_668), .A2(n_792), .B(n_793), .Y(n_791) );
INVx2_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g848 ( .A(n_669), .Y(n_848) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_677), .B2(n_678), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_676), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_687), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_685), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_688), .B(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g757 ( .A(n_696), .Y(n_757) );
OAI22xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_729), .B1(n_730), .B2(n_756), .Y(n_696) );
INVx1_ASAP7_75t_L g756 ( .A(n_697), .Y(n_756) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND3x1_ASAP7_75t_L g699 ( .A(n_700), .B(n_713), .C(n_719), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_707), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_717), .Y(n_713) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_721), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_746), .Y(n_733) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_740), .C(n_743), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_751), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_755), .Y(n_751) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OA22x2_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_782), .B2(n_825), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
XOR2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_781), .Y(n_762) );
NAND4xp75_ASAP7_75t_SL g763 ( .A(n_764), .B(n_774), .C(n_779), .D(n_780), .Y(n_763) );
NOR2xp67_ASAP7_75t_SL g764 ( .A(n_765), .B(n_770), .Y(n_764) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .C(n_769), .Y(n_765) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g825 ( .A(n_782), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B1(n_806), .B2(n_807), .Y(n_782) );
INVx1_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
XNOR2x1_ASAP7_75t_L g784 ( .A(n_785), .B(n_805), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_798), .Y(n_785) );
NOR3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_791), .C(n_794), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_802), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
INVx3_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
XOR2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_824), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g808 ( .A(n_809), .B(n_816), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_813), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_820), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_823), .Y(n_820) );
INVx1_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
NOR2x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_834), .Y(n_829) );
OR2x2_ASAP7_75t_SL g898 ( .A(n_830), .B(n_835), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_833), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_831), .Y(n_866) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_832), .B(n_870), .Y(n_874) );
CKINVDCx16_ASAP7_75t_R g870 ( .A(n_833), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
OAI322xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_865), .A3(n_867), .B1(n_871), .B2(n_875), .C1(n_876), .C2(n_896), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g843 ( .A(n_844), .Y(n_843) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND3xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_857), .C(n_861), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_852), .Y(n_846) );
OAI21xp5_ASAP7_75t_SL g847 ( .A1(n_848), .A2(n_849), .B(n_850), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .Y(n_852) );
INVx1_ASAP7_75t_SL g855 ( .A(n_856), .Y(n_855) );
AND2x2_ASAP7_75t_L g857 ( .A(n_858), .B(n_860), .Y(n_857) );
AND2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_SL g878 ( .A(n_879), .Y(n_878) );
NAND4xp75_ASAP7_75t_SL g879 ( .A(n_880), .B(n_886), .C(n_892), .D(n_895), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_885), .Y(n_880) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
AND2x2_ASAP7_75t_L g886 ( .A(n_887), .B(n_890), .Y(n_886) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
AND2x2_ASAP7_75t_SL g892 ( .A(n_893), .B(n_894), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_897), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_898), .Y(n_897) );
endmodule