module fake_jpeg_13702_n_379 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_379);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_379;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_50),
.B(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_53),
.Y(n_147)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_25),
.B(n_14),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_55),
.B(n_61),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_56),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_26),
.A2(n_14),
.B1(n_11),
.B2(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_57),
.A2(n_88),
.B1(n_20),
.B2(n_37),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_87),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_69),
.B(n_79),
.Y(n_128)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_30),
.B(n_1),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_73),
.A2(n_94),
.B(n_21),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx2_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_31),
.B(n_1),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_81),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

NAND2x1_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_91),
.Y(n_146)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_85),
.B(n_96),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_20),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_26),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_93),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_32),
.B(n_3),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_47),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_23),
.B(n_3),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_27),
.B1(n_48),
.B2(n_22),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_97),
.A2(n_45),
.B1(n_38),
.B2(n_18),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_134),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_5),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_111),
.B(n_131),
.CI(n_133),
.CON(n_181),
.SN(n_181)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_54),
.A2(n_27),
.B1(n_24),
.B2(n_43),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_112),
.A2(n_126),
.B1(n_109),
.B2(n_107),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_38),
.B1(n_43),
.B2(n_80),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_28),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_132),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_68),
.A2(n_24),
.B1(n_43),
.B2(n_19),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_59),
.B(n_48),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_127),
.B(n_137),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_77),
.C(n_63),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_87),
.B(n_22),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_71),
.B(n_33),
.C(n_42),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_33),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_70),
.A2(n_21),
.B(n_39),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_59),
.B(n_37),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_87),
.B(n_39),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_145),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_67),
.B(n_19),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_58),
.B(n_78),
.C(n_82),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_113),
.B(n_123),
.C(n_102),
.Y(n_191)
);

AOI32xp33_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_58),
.A3(n_95),
.B1(n_42),
.B2(n_45),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_150),
.B(n_135),
.CI(n_102),
.CON(n_195),
.SN(n_195)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_155),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_131),
.A2(n_93),
.B1(n_90),
.B2(n_81),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_158),
.B1(n_174),
.B2(n_178),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_166),
.B1(n_180),
.B2(n_118),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_136),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_101),
.C(n_135),
.Y(n_211)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_171),
.Y(n_194)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_116),
.A2(n_8),
.B(n_9),
.C(n_111),
.Y(n_167)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_130),
.A3(n_103),
.B1(n_116),
.B2(n_120),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_98),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_169),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_99),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_106),
.A2(n_9),
.B1(n_136),
.B2(n_105),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_118),
.B(n_107),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_121),
.A2(n_117),
.B1(n_104),
.B2(n_146),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_179),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_104),
.A2(n_117),
.B1(n_146),
.B2(n_148),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_183),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_98),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_184),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_213),
.B1(n_214),
.B2(n_174),
.Y(n_221)
);

AND2x4_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_113),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_209),
.C(n_211),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_191),
.A2(n_206),
.B1(n_149),
.B2(n_156),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_116),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_212),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_201),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_122),
.B1(n_129),
.B2(n_143),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_150),
.B1(n_172),
.B2(n_164),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_162),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_161),
.Y(n_230)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_181),
.C(n_170),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_162),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_122),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_159),
.A2(n_129),
.B1(n_141),
.B2(n_138),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_141),
.B1(n_138),
.B2(n_120),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_170),
.B(n_101),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_218),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_158),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_109),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_219),
.A2(n_206),
.B(n_191),
.Y(n_259)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_221),
.A2(n_231),
.B1(n_242),
.B2(n_243),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_172),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_225),
.C(n_215),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_193),
.A2(n_167),
.B1(n_149),
.B2(n_166),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_233),
.Y(n_264)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_229),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_230),
.B(n_240),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_175),
.B1(n_173),
.B2(n_169),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_193),
.A2(n_160),
.B1(n_163),
.B2(n_184),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_176),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_234),
.B(n_202),
.Y(n_245)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_171),
.B1(n_152),
.B2(n_155),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_237),
.A2(n_244),
.B1(n_200),
.B2(n_186),
.Y(n_263)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_209),
.B(n_151),
.CI(n_153),
.CON(n_240),
.SN(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_164),
.B1(n_155),
.B2(n_124),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_195),
.A2(n_100),
.B1(n_124),
.B2(n_204),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_248),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_188),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_247),
.B(n_250),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_238),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_188),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_216),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_196),
.B(n_218),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_227),
.B(n_210),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_225),
.B(n_202),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_258),
.Y(n_277)
);

AND2x6_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_209),
.Y(n_257)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_268),
.A3(n_189),
.B1(n_195),
.B2(n_201),
.C1(n_204),
.C2(n_226),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_196),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_259),
.A2(n_243),
.B(n_191),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_232),
.B(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_231),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_189),
.C(n_211),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_236),
.C(n_189),
.Y(n_283)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_203),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_228),
.B1(n_233),
.B2(n_220),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_269),
.A2(n_264),
.B1(n_256),
.B2(n_258),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_236),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_282),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_284),
.B(n_253),
.Y(n_299)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_281),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_246),
.A2(n_221),
.B1(n_219),
.B2(n_234),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_256),
.B1(n_264),
.B2(n_245),
.Y(n_301)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_247),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_232),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_286),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_218),
.B(n_216),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_262),
.Y(n_303)
);

XNOR2x2_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_262),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_289),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_205),
.C(n_194),
.Y(n_289)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_304),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_274),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_300),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_284),
.B(n_289),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_265),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_269),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_279),
.B1(n_270),
.B2(n_272),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_305),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_250),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_273),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_260),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_306),
.B(n_277),
.Y(n_309)
);

XOR2x2_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_313),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_310),
.A2(n_311),
.B1(n_314),
.B2(n_301),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_285),
.B1(n_276),
.B2(n_270),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_315),
.C(n_317),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_277),
.B1(n_275),
.B2(n_237),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_271),
.C(n_283),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_299),
.B(n_295),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_271),
.C(n_288),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_288),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_320),
.C(n_323),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_287),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_257),
.C(n_260),
.Y(n_323)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_327),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_319),
.B(n_291),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_328),
.B(n_334),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_304),
.Y(n_330)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_330),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_331),
.A2(n_317),
.B1(n_298),
.B2(n_296),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_290),
.C(n_300),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_307),
.Y(n_335)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_335),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_307),
.Y(n_336)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_336),
.Y(n_343)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_320),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_323),
.A2(n_296),
.B(n_298),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_339),
.A2(n_254),
.B(n_251),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_336),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_309),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_344),
.B(n_347),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_337),
.B(n_312),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_340),
.B(n_326),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_345),
.B(n_327),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_352),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_329),
.C(n_339),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_318),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_353),
.A2(n_343),
.B(n_332),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_358),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_329),
.C(n_332),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_359),
.C(n_333),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_346),
.B(n_330),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_356),
.A2(n_340),
.B1(n_343),
.B2(n_335),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_363),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_362),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_L g362 ( 
.A1(n_355),
.A2(n_349),
.A3(n_333),
.B1(n_251),
.B2(n_244),
.C1(n_229),
.C2(n_241),
.Y(n_362)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_365),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_353),
.A2(n_261),
.B(n_239),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_366),
.A2(n_244),
.B(n_267),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_368),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_364),
.A2(n_261),
.B(n_267),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_370),
.A2(n_207),
.B(n_242),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_L g372 ( 
.A1(n_371),
.A2(n_363),
.B(n_207),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_373),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_374),
.B(n_369),
.C(n_367),
.Y(n_375)
);

OAI321xp33_ASAP7_75t_L g377 ( 
.A1(n_375),
.A2(n_229),
.A3(n_235),
.B1(n_223),
.B2(n_200),
.C(n_190),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_376),
.C(n_194),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_378),
.A2(n_194),
.B(n_235),
.Y(n_379)
);


endmodule