module fake_jpeg_27490_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_16),
.B1(n_24),
.B2(n_30),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_17),
.B(n_22),
.C(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_59),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_18),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_53),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_18),
.B1(n_16),
.B2(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_16),
.B1(n_18),
.B2(n_31),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_16),
.B1(n_32),
.B2(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_27),
.B1(n_19),
.B2(n_23),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_27),
.B1(n_33),
.B2(n_29),
.Y(n_66)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_17),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_76),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_67),
.B1(n_73),
.B2(n_79),
.Y(n_109)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_31),
.B1(n_24),
.B2(n_30),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_72),
.B1(n_83),
.B2(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

OR2x6_ASAP7_75t_SL g110 ( 
.A(n_70),
.B(n_85),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_53),
.B1(n_51),
.B2(n_44),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_80),
.Y(n_105)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_31),
.B1(n_24),
.B2(n_30),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_28),
.B1(n_23),
.B2(n_17),
.Y(n_85)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_90),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_33),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_43),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_29),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_89),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_43),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_93),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_43),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_43),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_48),
.B(n_61),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_112),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_32),
.B1(n_58),
.B2(n_20),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_123),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_32),
.B1(n_22),
.B2(n_20),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_122),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_36),
.B(n_35),
.C(n_37),
.Y(n_118)
);

AOI211xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_74),
.B(n_91),
.C(n_69),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_42),
.B1(n_37),
.B2(n_38),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_63),
.B1(n_73),
.B2(n_67),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_69),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_126),
.B(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_65),
.B1(n_121),
.B2(n_106),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_103),
.B1(n_100),
.B2(n_124),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_131),
.A2(n_150),
.B(n_107),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_147),
.B1(n_148),
.B2(n_152),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_74),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_135),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_75),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_136),
.B(n_138),
.Y(n_184)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_65),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_98),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_146),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_81),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_82),
.B1(n_79),
.B2(n_86),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_87),
.B1(n_97),
.B2(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_155),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_110),
.A2(n_90),
.B1(n_42),
.B2(n_37),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_10),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_36),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_160),
.A2(n_178),
.B1(n_102),
.B2(n_101),
.Y(n_205)
);

AOI21x1_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_118),
.B(n_98),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_170),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_168),
.B(n_125),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_113),
.B1(n_109),
.B2(n_100),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_143),
.B1(n_187),
.B2(n_154),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_135),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_180),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_103),
.B(n_120),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_175),
.B(n_185),
.Y(n_211)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_133),
.B(n_136),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_109),
.B(n_108),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_117),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_186),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_111),
.B1(n_112),
.B2(n_101),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_36),
.C(n_38),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_181),
.C(n_183),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_113),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_131),
.B(n_104),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_104),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_104),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_125),
.B(n_1),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_132),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_145),
.B1(n_150),
.B2(n_128),
.Y(n_189)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_127),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_194),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_128),
.B1(n_146),
.B2(n_142),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_205),
.B1(n_206),
.B2(n_209),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_196),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_197),
.B(n_203),
.Y(n_234)
);

OAI21x1_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_129),
.B(n_156),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_185),
.B(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_157),
.A2(n_102),
.B1(n_125),
.B2(n_84),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_102),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_84),
.B1(n_42),
.B2(n_38),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_167),
.B(n_84),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_212),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_182),
.B(n_7),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_171),
.C(n_170),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_215),
.C(n_192),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_181),
.C(n_183),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_173),
.Y(n_218)
);

OAI322xp33_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_162),
.A3(n_189),
.B1(n_165),
.B2(n_161),
.C1(n_12),
.C2(n_5),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_180),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_220),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_166),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_160),
.B1(n_175),
.B2(n_186),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_201),
.B1(n_200),
.B2(n_189),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_177),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_229),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_233),
.Y(n_243)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_238),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_246),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_192),
.C(n_188),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_211),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_247),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_179),
.C(n_188),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_248),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_233),
.B1(n_216),
.B2(n_217),
.Y(n_252)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_5),
.B(n_14),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_161),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_165),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_190),
.C(n_176),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_223),
.C(n_232),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_6),
.C(n_14),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_251),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_227),
.B(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_SL g256 ( 
.A(n_242),
.B(n_227),
.Y(n_256)
);

OA21x2_ASAP7_75t_SL g273 ( 
.A1(n_256),
.A2(n_264),
.B(n_15),
.Y(n_273)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_8),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_216),
.B1(n_224),
.B2(n_226),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_15),
.B1(n_13),
.B2(n_11),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_221),
.B(n_225),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_237),
.B(n_5),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_230),
.B1(n_8),
.B2(n_11),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_250),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_254),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_235),
.C(n_246),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_270),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_238),
.B(n_235),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_276),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_273),
.B(n_275),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_265),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_263),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_11),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_253),
.B1(n_265),
.B2(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_278),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_283),
.B(n_285),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_254),
.B1(n_257),
.B2(n_260),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_284),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_282),
.A2(n_271),
.B(n_272),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_0),
.B(n_2),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_281),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_276),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_281),
.C(n_268),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_274),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_293),
.B(n_295),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_286),
.C1(n_290),
.C2(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_297),
.B(n_3),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_4),
.Y(n_300)
);


endmodule