module fake_jpeg_23545_n_163 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_163);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_43),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_40),
.Y(n_47)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_26),
.B1(n_17),
.B2(n_28),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_30),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_1),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_46),
.B(n_64),
.Y(n_89)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_25),
.CI(n_15),
.CON(n_48),
.SN(n_48)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_56),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_21),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_2),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_59),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_21),
.B1(n_23),
.B2(n_27),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_23),
.B1(n_15),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_41),
.B1(n_37),
.B2(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_68),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_22),
.B1(n_26),
.B2(n_17),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_69),
.B1(n_7),
.B2(n_8),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_32),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_65),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_1),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_28),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_70),
.Y(n_100)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_87),
.B(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_52),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_6),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_3),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_8),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_49),
.C(n_48),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_10),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_102),
.B(n_79),
.Y(n_113)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_59),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_109),
.B(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_54),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_89),
.B(n_78),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_121),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_115),
.C(n_123),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_50),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_91),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_93),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_47),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_125),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_72),
.B1(n_77),
.B2(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_99),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_120),
.B(n_108),
.Y(n_144)
);

AO221x1_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_103),
.B1(n_95),
.B2(n_106),
.C(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

AO221x1_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_107),
.B1(n_86),
.B2(n_104),
.C(n_81),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_139),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_125),
.B1(n_96),
.B2(n_117),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_136),
.A2(n_96),
.B1(n_118),
.B2(n_115),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_123),
.C(n_129),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_104),
.C(n_55),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_144),
.A2(n_129),
.B(n_126),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_142),
.B(n_143),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_53),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_145),
.C(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_149),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_156),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_140),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_150),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_159),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_153),
.A3(n_152),
.B1(n_81),
.B2(n_82),
.C1(n_13),
.C2(n_10),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_82),
.B(n_157),
.C(n_90),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_160),
.Y(n_163)
);


endmodule