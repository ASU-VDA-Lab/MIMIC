module fake_jpeg_20275_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

AO22x1_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_44),
.Y(n_53)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_45),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_47),
.B(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_31),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_61),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_17),
.B1(n_26),
.B2(n_18),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_62),
.B1(n_39),
.B2(n_42),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_42),
.B1(n_41),
.B2(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_35),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_66),
.C(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_26),
.B(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_17),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_74),
.Y(n_120)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_78),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_76),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_33),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_75),
.B(n_95),
.C(n_21),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_80),
.Y(n_125)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_83),
.B1(n_91),
.B2(n_93),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_33),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_87),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_42),
.B1(n_41),
.B2(n_39),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_53),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_41),
.B1(n_39),
.B2(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_22),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_18),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_28),
.B1(n_24),
.B2(n_34),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_28),
.B1(n_34),
.B2(n_27),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_112),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_110),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_102),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_26),
.B1(n_29),
.B2(n_21),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_132),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_32),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_30),
.Y(n_128)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_128),
.B(n_30),
.CI(n_22),
.CON(n_145),
.SN(n_145)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_95),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_81),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_111),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_83),
.B(n_86),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_140),
.B(n_142),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_89),
.B1(n_105),
.B2(n_83),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_137),
.A2(n_165),
.B1(n_157),
.B2(n_158),
.Y(n_198)
);

BUFx12_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_70),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_141),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_69),
.B(n_74),
.C(n_53),
.D(n_93),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_107),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_84),
.B1(n_90),
.B2(n_94),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_130),
.B(n_29),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_143),
.B(n_160),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_35),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_149),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_67),
.B1(n_1),
.B2(n_2),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_152),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_30),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_23),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_77),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_84),
.B(n_1),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_164),
.B(n_110),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_108),
.A2(n_88),
.B(n_85),
.C(n_99),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_119),
.B(n_127),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_32),
.B1(n_19),
.B2(n_98),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_113),
.B(n_77),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_121),
.Y(n_184)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_22),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_108),
.A2(n_79),
.B1(n_40),
.B2(n_38),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_135),
.C(n_127),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_170),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_128),
.C(n_129),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_178),
.C(n_193),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_124),
.B(n_117),
.C(n_134),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_160),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_179),
.Y(n_212)
);

AOI21x1_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_88),
.B(n_119),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_173),
.A2(n_175),
.B(n_182),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_151),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_188),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_121),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_189),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_134),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_142),
.B(n_146),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_144),
.B(n_14),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_40),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_190),
.A2(n_148),
.B1(n_157),
.B2(n_155),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_196),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_40),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_40),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_38),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_187),
.B1(n_191),
.B2(n_189),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_198),
.B1(n_197),
.B2(n_190),
.Y(n_227)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_157),
.B1(n_142),
.B2(n_153),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_187),
.B(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_206),
.B(n_208),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_217),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_210),
.B(n_218),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_216),
.C(n_174),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_185),
.C(n_182),
.Y(n_216)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_154),
.B(n_138),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

XNOR2x2_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_170),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_219),
.B(n_194),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_222),
.Y(n_229)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_224),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_168),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_226),
.A2(n_230),
.B(n_236),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_217),
.B1(n_221),
.B2(n_203),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_180),
.B(n_194),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_163),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_171),
.C(n_138),
.Y(n_243)
);

A2O1A1O1Ixp25_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_207),
.B(n_223),
.C(n_225),
.D(n_216),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_230),
.A2(n_207),
.B1(n_202),
.B2(n_220),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_255),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_244),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_214),
.C(n_211),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_258),
.C(n_261),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_212),
.B1(n_217),
.B2(n_215),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_259),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_234),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_222),
.C(n_166),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_242),
.A2(n_96),
.B1(n_25),
.B2(n_35),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_227),
.A2(n_25),
.B1(n_35),
.B2(n_23),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_260),
.B(n_265),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_96),
.C(n_25),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_228),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_231),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_25),
.C(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_274),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_239),
.C(n_241),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_275),
.C(n_278),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_236),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_247),
.C(n_246),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_233),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_263),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_247),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_243),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_240),
.C(n_226),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_259),
.B1(n_262),
.B2(n_248),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_281),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_270),
.A2(n_251),
.B(n_254),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_6),
.B(n_7),
.Y(n_300)
);

NOR3xp33_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_254),
.C(n_240),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_289),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_252),
.B(n_229),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_229),
.B(n_265),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_292),
.B(n_298),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_286),
.A2(n_281),
.B1(n_288),
.B2(n_274),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_300),
.B1(n_287),
.B2(n_7),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_269),
.C(n_5),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_297),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_4),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_5),
.C(n_6),
.Y(n_298)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_287),
.B(n_7),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_304),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_12),
.C2(n_13),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_293),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_301),
.B(n_305),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_299),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_310),
.A2(n_311),
.B(n_309),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_294),
.B(n_12),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_9),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_13),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_13),
.Y(n_315)
);


endmodule