module fake_netlist_1_84_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVx3_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
BUFx16f_ASAP7_75t_R g5 ( .A(n_1), .Y(n_5) );
OAI21xp5_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_6) );
OAI21x1_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_0), .B(n_2), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_4), .A2(n_0), .B(n_2), .Y(n_8) );
INVxp67_ASAP7_75t_SL g9 ( .A(n_6), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_7), .B(n_3), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_9), .B(n_7), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
NAND4xp75_ASAP7_75t_L g13 ( .A(n_11), .B(n_5), .C(n_8), .D(n_10), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_12), .B(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
OA21x2_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_11), .B(n_12), .Y(n_17) );
AOI22xp33_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_3), .B1(n_16), .B2(n_15), .Y(n_18) );
endmodule