module fake_jpeg_7826_n_226 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_2),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_47),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_25),
.B1(n_30),
.B2(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_35),
.B1(n_20),
.B2(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_57),
.A2(n_60),
.B1(n_69),
.B2(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_66),
.B1(n_26),
.B2(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_60)
);

CKINVDCx12_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_48),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_1),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_35),
.B1(n_20),
.B2(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_41),
.B1(n_22),
.B2(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_22),
.B1(n_28),
.B2(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_72),
.B(n_73),
.Y(n_121)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_76),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_75),
.B(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_79),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_46),
.B1(n_43),
.B2(n_31),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_29),
.B1(n_26),
.B2(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_84),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_76),
.B1(n_74),
.B2(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_10),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_92),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_49),
.B(n_37),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_2),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_68),
.B1(n_62),
.B2(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_24),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_97),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_24),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_95),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_89),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_84),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_109),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_24),
.B1(n_14),
.B2(n_12),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_110),
.B1(n_81),
.B2(n_71),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_1),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_120),
.B(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_3),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_124),
.B(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_71),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_129),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_120),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_134),
.C(n_136),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_128),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_95),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_132),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_141),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_73),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_91),
.C(n_98),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_75),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_83),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_142),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_78),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_77),
.C(n_5),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_5),
.Y(n_166)
);

OAI22x1_ASAP7_75t_SL g146 ( 
.A1(n_108),
.A2(n_79),
.B1(n_77),
.B2(n_99),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_77),
.B1(n_90),
.B2(n_116),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_100),
.B1(n_118),
.B2(n_110),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_152),
.B1(n_116),
.B2(n_7),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_106),
.B(n_114),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_148),
.A2(n_150),
.B(n_151),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_114),
.B(n_100),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_117),
.B(n_118),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_117),
.B1(n_105),
.B2(n_90),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_155),
.B(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_166),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_133),
.B1(n_137),
.B2(n_125),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_3),
.B(n_5),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_127),
.B(n_7),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_181),
.B1(n_149),
.B2(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_174),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_178),
.B(n_179),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_177),
.B1(n_162),
.B2(n_157),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_163),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_9),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_6),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_180),
.C(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_6),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_160),
.B(n_6),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_184),
.C(n_186),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_158),
.C(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_153),
.C(n_175),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_172),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_148),
.C(n_150),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_191),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_147),
.B1(n_152),
.B2(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_193),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_176),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_183),
.C(n_190),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_171),
.C(n_179),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_187),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_174),
.B(n_173),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_8),
.B1(n_9),
.B2(n_201),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_200),
.B(n_184),
.CI(n_191),
.CON(n_205),
.SN(n_205)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_209),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_198),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_8),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_205),
.Y(n_219)
);

NAND3xp33_ASAP7_75t_SL g216 ( 
.A(n_212),
.B(n_209),
.C(n_205),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_197),
.B(n_215),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_208),
.B(n_197),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_202),
.C(n_218),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_202),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_220),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_222),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_223),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_224),
.Y(n_226)
);


endmodule