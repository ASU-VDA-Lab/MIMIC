module fake_jpeg_1041_n_186 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_34),
.B(n_44),
.Y(n_78)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_45),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_16),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_53),
.Y(n_64)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_71),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_15),
.B1(n_22),
.B2(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_15),
.B1(n_22),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_31),
.B1(n_29),
.B2(n_24),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_23),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_51),
.B1(n_49),
.B2(n_35),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_19),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_82),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_46),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_59),
.C(n_79),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_52),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_31),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_92),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_43),
.B(n_20),
.C(n_19),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_94),
.B(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_17),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_96),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_8),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_88),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_103),
.B1(n_84),
.B2(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_2),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_65),
.B1(n_73),
.B2(n_85),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_5),
.B(n_14),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_75),
.B(n_81),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_57),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_56),
.B1(n_72),
.B2(n_59),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_100),
.Y(n_109)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_68),
.A2(n_79),
.B1(n_67),
.B2(n_55),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_95),
.Y(n_123)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_91),
.B(n_104),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_72),
.B(n_57),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_121),
.B(n_86),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_103),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_95),
.C(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_125),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_65),
.B(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_105),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_127),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_119),
.Y(n_127)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_99),
.B(n_86),
.C(n_84),
.D(n_90),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_136),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_115),
.B1(n_107),
.B2(n_110),
.Y(n_153)
);

AOI21x1_ASAP7_75t_SL g149 ( 
.A1(n_139),
.A2(n_109),
.B(n_106),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_106),
.C(n_114),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_82),
.B1(n_109),
.B2(n_107),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_141),
.A2(n_113),
.B(n_121),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_117),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_146),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_149),
.B(n_151),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_116),
.C(n_124),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_116),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_111),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_153),
.B(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_159),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_139),
.B(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

OA21x2_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_142),
.B(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_170),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_138),
.B1(n_149),
.B2(n_146),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_168),
.A2(n_140),
.B1(n_129),
.B2(n_125),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_111),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_169),
.A2(n_158),
.B(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_175),
.B(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_153),
.B1(n_157),
.B2(n_138),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_179),
.B(n_129),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_174),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_166),
.B(n_165),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_181),
.B(n_128),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_176),
.C(n_128),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_183),
.B(n_137),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_107),
.Y(n_186)
);


endmodule