module fake_jpeg_16699_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_9),
.B(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_51),
.Y(n_76)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_0),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_58),
.Y(n_72)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_72),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_57),
.B1(n_47),
.B2(n_53),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_54),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_44),
.B1(n_43),
.B2(n_48),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_55),
.B1(n_60),
.B2(n_2),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_60),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_50),
.B1(n_55),
.B2(n_46),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_96),
.B1(n_84),
.B2(n_89),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_98),
.C(n_83),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_72),
.B1(n_18),
.B2(n_19),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_100),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_5),
.Y(n_113)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_113),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_95),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_92),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_91),
.B(n_7),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_91),
.B1(n_7),
.B2(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_120),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_126),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_106),
.C(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_99),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_104),
.B1(n_109),
.B2(n_106),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_125),
.A2(n_110),
.B1(n_14),
.B2(n_15),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_13),
.B1(n_17),
.B2(n_20),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_134),
.B1(n_133),
.B2(n_124),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_134),
.A2(n_22),
.B(n_24),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_26),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_27),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_32),
.B(n_34),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_35),
.C(n_36),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_37),
.B(n_39),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_40),
.Y(n_146)
);


endmodule